module channel_reduce_4(input [0:0] clk, input [0:0] rst, output [0:0] valid, output [31:0] in_in_data, input [31:0] in_out_data, input [0:0] in_read_ready, output [0:0] in_read_valid, input [0:0] in_write_ready, output [0:0] in_write_valid, output [31:0] out_in_data, input [31:0] out_out_data, input [0:0] out_read_ready, output [0:0] out_read_valid, input [0:0] out_write_ready, output [0:0] out_write_valid);

	reg [0:0] valid_reg;
	reg [31:0] in_in_data_reg;
	reg [0:0] in_read_valid_reg;
	reg [0:0] in_write_valid_reg;
	reg [31:0] out_in_data_reg;
	reg [0:0] out_read_valid_reg;
	reg [0:0] out_write_valid_reg;

	assign valid = valid_reg;
	assign in_in_data = in_in_data_reg;
	assign in_read_valid = in_read_valid_reg;
	assign in_write_valid = in_write_valid_reg;
	assign out_in_data = out_in_data_reg;
	assign out_read_valid = out_read_valid_reg;
	assign out_write_valid = out_write_valid_reg;

	// Start debug wires and ports

	initial begin
	end





	// End debug wires and ports

	// Start Functional Units
	br_dummy br_unit();

	reg [31:0] raddr_ram_0_reg;
	reg [31:0] waddr_ram_0_reg;
	reg [31:0] wdata_ram_0_reg;
	reg [0:0] wen_ram_0_reg;
	wire [31:0] rdata_ram_0;
	register #(.WIDTH(32)) ram_0(.clk(clk), .raddr(raddr_ram_0_reg), .rdata(rdata_ram_0), .rst(rst), .waddr(waddr_ram_0_reg), .wdata(wdata_ram_0_reg), .wen(wen_ram_0_reg));

	wire [31:0] add_add13_in0;
	wire [31:0] add_add13_in1;
	wire [31:0] add_add13_out;
	add #(.WIDTH(32)) add_add13(.in0(add_add13_in0), .in1(add_add13_in1), .out(add_add13_out));

	wire [31:0] add_add15_in0;
	wire [31:0] add_add15_in1;
	wire [31:0] add_add15_out;
	add #(.WIDTH(32)) add_add15(.in0(add_add15_in0), .in1(add_add15_in1), .out(add_add15_out));

	wire [31:0] icmp_icmp16_in0;
	wire [31:0] icmp_icmp16_in1;
	wire [0:0] icmp_icmp16_out;
	eq #(.WIDTH(32)) icmp_icmp16(.in0(icmp_icmp16_in0), .in1(icmp_icmp16_in1), .out(icmp_icmp16_out));

	add call25();

	wire [63:0] phi_phi6_in;
	wire [31:0] phi_phi6_last_block;
	wire [63:0] phi_phi6_s;
	wire [31:0] phi_phi6_out;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_phi6(.in(phi_phi6_in), .last_block(phi_phi6_last_block), .out(phi_phi6_out), .s(phi_phi6_s));

	add alloca0();

	add bitcast1();

	add call2();

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] bb_0_active_in_state_1_in_data;
	wire [0:0] bb_0_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_1(.in_data(bb_0_active_in_state_1_in_data), .out_data(bb_0_active_in_state_1_out_data));

	reg [31:0] bb_0_predecessor_in_state_1_in_data;
	wire [31:0] bb_0_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_1(.in_data(bb_0_predecessor_in_state_1_in_data), .out_data(bb_0_predecessor_in_state_1_out_data));

	reg [0:0] br_0_happened_in_state_1_in_data;
	wire [0:0] br_0_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_1(.in_data(br_0_happened_in_state_1_in_data), .out_data(br_0_happened_in_state_1_out_data));

	reg [0:0] bb_8_active_in_state_1_in_data;
	wire [0:0] bb_8_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active_in_state_1(.in_data(bb_8_active_in_state_1_in_data), .out_data(bb_8_active_in_state_1_out_data));

	reg [31:0] bb_8_predecessor_in_state_1_in_data;
	wire [31:0] bb_8_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor_in_state_1(.in_data(bb_8_predecessor_in_state_1_in_data), .out_data(bb_8_predecessor_in_state_1_out_data));

	reg [0:0] br_8_happened_in_state_1_in_data;
	wire [0:0] br_8_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_8_happened_in_state_1(.in_data(br_8_happened_in_state_1_in_data), .out_data(br_8_happened_in_state_1_out_data));

	reg [0:0] bb_3_active_in_state_1_in_data;
	wire [0:0] bb_3_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_1(.in_data(bb_3_active_in_state_1_in_data), .out_data(bb_3_active_in_state_1_out_data));

	reg [31:0] bb_3_predecessor_in_state_1_in_data;
	wire [31:0] bb_3_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_1(.in_data(bb_3_predecessor_in_state_1_in_data), .out_data(bb_3_predecessor_in_state_1_out_data));

	reg [0:0] br_3_happened_in_state_1_in_data;
	wire [0:0] br_3_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_1(.in_data(br_3_happened_in_state_1_in_data), .out_data(br_3_happened_in_state_1_out_data));

	reg [0:0] bb_9_active_in_state_1_in_data;
	wire [0:0] bb_9_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_9_active_in_state_1(.in_data(bb_9_active_in_state_1_in_data), .out_data(bb_9_active_in_state_1_out_data));

	reg [31:0] bb_9_predecessor_in_state_1_in_data;
	wire [31:0] bb_9_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_9_predecessor_in_state_1(.in_data(bb_9_predecessor_in_state_1_in_data), .out_data(bb_9_predecessor_in_state_1_out_data));

	reg [0:0] br_9_happened_in_state_1_in_data;
	wire [0:0] br_9_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_9_happened_in_state_1(.in_data(br_9_happened_in_state_1_in_data), .out_data(br_9_happened_in_state_1_out_data));

	reg [0:0] bb_10_active_in_state_2_in_data;
	wire [0:0] bb_10_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_2(.in_data(bb_10_active_in_state_2_in_data), .out_data(bb_10_active_in_state_2_out_data));

	reg [31:0] bb_10_predecessor_in_state_2_in_data;
	wire [31:0] bb_10_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_2(.in_data(bb_10_predecessor_in_state_2_in_data), .out_data(bb_10_predecessor_in_state_2_out_data));

	reg [0:0] br_10_happened_in_state_2_in_data;
	wire [0:0] br_10_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_2(.in_data(br_10_happened_in_state_2_in_data), .out_data(br_10_happened_in_state_2_out_data));

	reg [0:0] bb_4_active_in_state_3_in_data;
	wire [0:0] bb_4_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_3(.in_data(bb_4_active_in_state_3_in_data), .out_data(bb_4_active_in_state_3_out_data));

	reg [31:0] bb_4_predecessor_in_state_3_in_data;
	wire [31:0] bb_4_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_3(.in_data(bb_4_predecessor_in_state_3_in_data), .out_data(bb_4_predecessor_in_state_3_out_data));

	reg [0:0] br_4_happened_in_state_3_in_data;
	wire [0:0] br_4_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_3(.in_data(br_4_happened_in_state_3_in_data), .out_data(br_4_happened_in_state_3_out_data));

	reg [0:0] bb_10_active_in_state_3_in_data;
	wire [0:0] bb_10_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_3(.in_data(bb_10_active_in_state_3_in_data), .out_data(bb_10_active_in_state_3_out_data));

	reg [31:0] bb_10_predecessor_in_state_3_in_data;
	wire [31:0] bb_10_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_3(.in_data(bb_10_predecessor_in_state_3_in_data), .out_data(bb_10_predecessor_in_state_3_out_data));

	reg [0:0] br_10_happened_in_state_3_in_data;
	wire [0:0] br_10_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_3(.in_data(br_10_happened_in_state_3_in_data), .out_data(br_10_happened_in_state_3_out_data));

	reg [0:0] bb_4_active_in_state_4_in_data;
	wire [0:0] bb_4_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_4(.in_data(bb_4_active_in_state_4_in_data), .out_data(bb_4_active_in_state_4_out_data));

	reg [31:0] bb_4_predecessor_in_state_4_in_data;
	wire [31:0] bb_4_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_4(.in_data(bb_4_predecessor_in_state_4_in_data), .out_data(bb_4_predecessor_in_state_4_out_data));

	reg [0:0] br_4_happened_in_state_4_in_data;
	wire [0:0] br_4_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_4(.in_data(br_4_happened_in_state_4_in_data), .out_data(br_4_happened_in_state_4_out_data));

	reg [0:0] bb_6_active_in_state_4_in_data;
	wire [0:0] bb_6_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_6_active_in_state_4(.in_data(bb_6_active_in_state_4_in_data), .out_data(bb_6_active_in_state_4_out_data));

	reg [31:0] bb_6_predecessor_in_state_4_in_data;
	wire [31:0] bb_6_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_6_predecessor_in_state_4(.in_data(bb_6_predecessor_in_state_4_in_data), .out_data(bb_6_predecessor_in_state_4_out_data));

	reg [0:0] br_6_happened_in_state_4_in_data;
	wire [0:0] br_6_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_6_happened_in_state_4(.in_data(br_6_happened_in_state_4_in_data), .out_data(br_6_happened_in_state_4_out_data));

	reg [0:0] bb_2_active_in_state_4_in_data;
	wire [0:0] bb_2_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_4(.in_data(bb_2_active_in_state_4_in_data), .out_data(bb_2_active_in_state_4_out_data));

	reg [31:0] bb_2_predecessor_in_state_4_in_data;
	wire [31:0] bb_2_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_4(.in_data(bb_2_predecessor_in_state_4_in_data), .out_data(bb_2_predecessor_in_state_4_out_data));

	reg [0:0] bb_5_active_in_state_4_in_data;
	wire [0:0] bb_5_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_5_active_in_state_4(.in_data(bb_5_active_in_state_4_in_data), .out_data(bb_5_active_in_state_4_out_data));

	reg [31:0] bb_5_predecessor_in_state_4_in_data;
	wire [31:0] bb_5_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_5_predecessor_in_state_4(.in_data(bb_5_predecessor_in_state_4_in_data), .out_data(bb_5_predecessor_in_state_4_out_data));

	reg [0:0] br_5_happened_in_state_4_in_data;
	wire [0:0] br_5_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_5_happened_in_state_4(.in_data(br_5_happened_in_state_4_in_data), .out_data(br_5_happened_in_state_4_out_data));

	reg [0:0] bb_7_active_in_state_4_in_data;
	wire [0:0] bb_7_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_7_active_in_state_4(.in_data(bb_7_active_in_state_4_in_data), .out_data(bb_7_active_in_state_4_out_data));

	reg [31:0] bb_7_predecessor_in_state_4_in_data;
	wire [31:0] bb_7_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_7_predecessor_in_state_4(.in_data(bb_7_predecessor_in_state_4_in_data), .out_data(bb_7_predecessor_in_state_4_out_data));

	reg [0:0] br_7_happened_in_state_4_in_data;
	wire [0:0] br_7_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_7_happened_in_state_4(.in_data(br_7_happened_in_state_4_in_data), .out_data(br_7_happened_in_state_4_out_data));

	reg [0:0] bb_1_active_in_state_4_in_data;
	wire [0:0] bb_1_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_4(.in_data(bb_1_active_in_state_4_in_data), .out_data(bb_1_active_in_state_4_out_data));

	reg [31:0] bb_1_predecessor_in_state_4_in_data;
	wire [31:0] bb_1_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_4(.in_data(bb_1_predecessor_in_state_4_in_data), .out_data(bb_1_predecessor_in_state_4_out_data));

	reg [0:0] br_1_happened_in_state_4_in_data;
	wire [0:0] br_1_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened_in_state_4(.in_data(br_1_happened_in_state_4_in_data), .out_data(br_1_happened_in_state_4_out_data));

	reg [31:0] data_in_0_1_in_data;
	wire [31:0] data_in_0_1_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_1(.in_data(data_in_0_1_in_data), .out_data(data_in_0_1_out_data));

	reg [31:0] data_in_0_3_in_data;
	wire [31:0] data_in_0_3_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_3(.in_data(data_in_0_3_in_data), .out_data(data_in_0_3_out_data));

	reg [31:0] data_in_1_5_in_data;
	wire [31:0] data_in_1_5_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_5(.in_data(data_in_1_5_in_data), .out_data(data_in_1_5_out_data));

	reg [31:0] data_in_1_7_in_data;
	wire [31:0] data_in_1_7_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_7(.in_data(data_in_1_7_in_data), .out_data(data_in_1_7_out_data));

	reg [31:0] data_in_2_9_in_data;
	wire [31:0] data_in_2_9_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_9(.in_data(data_in_2_9_in_data), .out_data(data_in_2_9_out_data));

	reg [31:0] data_in_3_13_in_data;
	wire [31:0] data_in_3_13_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_13(.in_data(data_in_3_13_in_data), .out_data(data_in_3_13_out_data));

	reg [31:0] data_in_4_15_in_data;
	wire [31:0] data_in_4_15_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_15(.in_data(data_in_4_15_in_data), .out_data(data_in_4_15_out_data));

	reg [0:0] data_in_4_17_in_data;
	wire [0:0] data_in_4_17_out_data;
	hls_wire #(.WIDTH(1)) data_in_4_17(.in_data(data_in_4_17_in_data), .out_data(data_in_4_17_out_data));

	reg [31:0] data_in_4_19_in_data;
	wire [31:0] data_in_4_19_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_19(.in_data(data_in_4_19_in_data), .out_data(data_in_4_19_out_data));

	wire [0:0] andOp_20_in0;
	wire [0:0] andOp_20_in1;
	wire [0:0] andOp_20_out;
	andOp #(.WIDTH(1)) andOp_20(.in0(andOp_20_in0), .in1(andOp_20_in1), .out(andOp_20_out));

	wire [0:0] notOp_21_in0;
	wire [0:0] notOp_21_out;
	notOp #(.WIDTH(1)) notOp_21(.in(notOp_21_in0), .out(notOp_21_out));

	wire [0:0] andOp_22_in0;
	wire [0:0] andOp_22_in1;
	wire [0:0] andOp_22_out;
	andOp #(.WIDTH(1)) andOp_22(.in0(andOp_22_in0), .in1(andOp_22_in1), .out(andOp_22_out));

	wire [0:0] notOp_23_in0;
	wire [0:0] notOp_23_out;
	notOp #(.WIDTH(1)) notOp_23(.in(notOp_23_in0), .out(notOp_23_out));

	wire [0:0] andOp_24_in0;
	wire [0:0] andOp_24_in1;
	wire [0:0] andOp_24_out;
	andOp #(.WIDTH(1)) andOp_24(.in0(andOp_24_in0), .in1(andOp_24_in1), .out(andOp_24_out));

	wire [0:0] notOp_25_in0;
	wire [0:0] notOp_25_out;
	notOp #(.WIDTH(1)) notOp_25(.in(notOp_25_in0), .out(notOp_25_out));

	wire [0:0] andOp_26_in0;
	wire [0:0] andOp_26_in1;
	wire [0:0] andOp_26_out;
	andOp #(.WIDTH(1)) andOp_26(.in0(andOp_26_in0), .in1(andOp_26_in1), .out(andOp_26_out));

	wire [0:0] notOp_27_in0;
	wire [0:0] notOp_27_out;
	notOp #(.WIDTH(1)) notOp_27(.in(notOp_27_in0), .out(notOp_27_out));

	wire [0:0] andOp_28_in0;
	wire [0:0] andOp_28_in1;
	wire [0:0] andOp_28_out;
	andOp #(.WIDTH(1)) andOp_28(.in0(andOp_28_in0), .in1(andOp_28_in1), .out(andOp_28_out));

	wire [0:0] notOp_29_in0;
	wire [0:0] notOp_29_out;
	notOp #(.WIDTH(1)) notOp_29(.in(notOp_29_in0), .out(notOp_29_out));

	wire [0:0] andOp_30_in0;
	wire [0:0] andOp_30_in1;
	wire [0:0] andOp_30_out;
	andOp #(.WIDTH(1)) andOp_30(.in0(andOp_30_in0), .in1(andOp_30_in1), .out(andOp_30_out));

	wire [0:0] notOp_31_in0;
	wire [0:0] notOp_31_out;
	notOp #(.WIDTH(1)) notOp_31(.in(notOp_31_in0), .out(notOp_31_out));

	wire [0:0] andOp_32_in0;
	wire [0:0] andOp_32_in1;
	wire [0:0] andOp_32_out;
	andOp #(.WIDTH(1)) andOp_32(.in0(andOp_32_in0), .in1(andOp_32_in1), .out(andOp_32_out));

	wire [0:0] andOp_33_in0;
	wire [0:0] andOp_33_in1;
	wire [0:0] andOp_33_out;
	andOp #(.WIDTH(1)) andOp_33(.in0(andOp_33_in0), .in1(andOp_33_in1), .out(andOp_33_out));

	wire [0:0] notOp_34_in0;
	wire [0:0] notOp_34_out;
	notOp #(.WIDTH(1)) notOp_34(.in(notOp_34_in0), .out(notOp_34_out));

	wire [0:0] andOp_35_in0;
	wire [0:0] andOp_35_in1;
	wire [0:0] andOp_35_out;
	andOp #(.WIDTH(1)) andOp_35(.in0(andOp_35_in0), .in1(andOp_35_in1), .out(andOp_35_out));

	wire [0:0] notOp_36_in0;
	wire [0:0] notOp_36_out;
	notOp #(.WIDTH(1)) notOp_36(.in(notOp_36_in0), .out(notOp_36_out));

	wire [0:0] andOp_37_in0;
	wire [0:0] andOp_37_in1;
	wire [0:0] andOp_37_out;
	andOp #(.WIDTH(1)) andOp_37(.in0(andOp_37_in0), .in1(andOp_37_in1), .out(andOp_37_out));

	wire [0:0] notOp_38_in0;
	wire [0:0] notOp_38_out;
	notOp #(.WIDTH(1)) notOp_38(.in(notOp_38_in0), .out(notOp_38_out));

	wire [0:0] andOp_39_in0;
	wire [0:0] andOp_39_in1;
	wire [0:0] andOp_39_out;
	andOp #(.WIDTH(1)) andOp_39(.in0(andOp_39_in0), .in1(andOp_39_in1), .out(andOp_39_out));

	wire [0:0] andOp_40_in0;
	wire [0:0] andOp_40_in1;
	wire [0:0] andOp_40_out;
	andOp #(.WIDTH(1)) andOp_40(.in0(andOp_40_in0), .in1(andOp_40_in1), .out(andOp_40_out));

	wire [0:0] notOp_41_in0;
	wire [0:0] notOp_41_out;
	notOp #(.WIDTH(1)) notOp_41(.in(notOp_41_in0), .out(notOp_41_out));

	wire [0:0] andOp_42_in0;
	wire [0:0] andOp_42_in1;
	wire [0:0] andOp_42_out;
	andOp #(.WIDTH(1)) andOp_42(.in0(andOp_42_in0), .in1(andOp_42_in1), .out(andOp_42_out));

	wire [0:0] notOp_43_in0;
	wire [0:0] notOp_43_out;
	notOp #(.WIDTH(1)) notOp_43(.in(notOp_43_in0), .out(notOp_43_out));

	wire [0:0] andOp_44_in0;
	wire [0:0] andOp_44_in1;
	wire [0:0] andOp_44_out;
	andOp #(.WIDTH(1)) andOp_44(.in0(andOp_44_in0), .in1(andOp_44_in1), .out(andOp_44_out));

	wire [0:0] notOp_45_in0;
	wire [0:0] notOp_45_out;
	notOp #(.WIDTH(1)) notOp_45(.in(notOp_45_in0), .out(notOp_45_out));

	wire [0:0] andOp_46_in0;
	wire [0:0] andOp_46_in1;
	wire [0:0] andOp_46_out;
	andOp #(.WIDTH(1)) andOp_46(.in0(andOp_46_in0), .in1(andOp_46_in1), .out(andOp_46_out));

	wire [0:0] andOp_47_in0;
	wire [0:0] andOp_47_in1;
	wire [0:0] andOp_47_out;
	andOp #(.WIDTH(1)) andOp_47(.in0(andOp_47_in0), .in1(andOp_47_in1), .out(andOp_47_out));

	wire [0:0] notOp_48_in0;
	wire [0:0] notOp_48_out;
	notOp #(.WIDTH(1)) notOp_48(.in(notOp_48_in0), .out(notOp_48_out));

	wire [0:0] andOp_49_in0;
	wire [0:0] andOp_49_in1;
	wire [0:0] andOp_49_out;
	andOp #(.WIDTH(1)) andOp_49(.in0(andOp_49_in0), .in1(andOp_49_in1), .out(andOp_49_out));

	wire [0:0] notOp_50_in0;
	wire [0:0] notOp_50_out;
	notOp #(.WIDTH(1)) notOp_50(.in(notOp_50_in0), .out(notOp_50_out));

	wire [0:0] andOp_51_in0;
	wire [0:0] andOp_51_in1;
	wire [0:0] andOp_51_out;
	andOp #(.WIDTH(1)) andOp_51(.in0(andOp_51_in0), .in1(andOp_51_in1), .out(andOp_51_out));

	wire [0:0] andOp_52_in0;
	wire [0:0] andOp_52_in1;
	wire [0:0] andOp_52_out;
	andOp #(.WIDTH(1)) andOp_52(.in0(andOp_52_in0), .in1(andOp_52_in1), .out(andOp_52_out));

	wire [0:0] notOp_53_in0;
	wire [0:0] notOp_53_out;
	notOp #(.WIDTH(1)) notOp_53(.in(notOp_53_in0), .out(notOp_53_out));

	wire [0:0] andOp_54_in0;
	wire [0:0] andOp_54_in1;
	wire [0:0] andOp_54_out;
	andOp #(.WIDTH(1)) andOp_54(.in0(andOp_54_in0), .in1(andOp_54_in1), .out(andOp_54_out));

	wire [0:0] notOp_55_in0;
	wire [0:0] notOp_55_out;
	notOp #(.WIDTH(1)) notOp_55(.in(notOp_55_in0), .out(notOp_55_out));

	wire [0:0] andOp_56_in0;
	wire [0:0] andOp_56_in1;
	wire [0:0] andOp_56_out;
	andOp #(.WIDTH(1)) andOp_56(.in0(andOp_56_in0), .in1(andOp_56_in1), .out(andOp_56_out));

	wire [0:0] notOp_57_in0;
	wire [0:0] notOp_57_out;
	notOp #(.WIDTH(1)) notOp_57(.in(notOp_57_in0), .out(notOp_57_out));

	wire [31:0] eq_58_in0;
	wire [31:0] eq_58_in1;
	wire [0:0] eq_58_out;
	eq #(.WIDTH(32)) eq_58(.in0(eq_58_in0), .in1(eq_58_in1), .out(eq_58_out));

	wire [31:0] eq_59_in0;
	wire [31:0] eq_59_in1;
	wire [0:0] eq_59_out;
	eq #(.WIDTH(32)) eq_59(.in0(eq_59_in0), .in1(eq_59_in1), .out(eq_59_out));

	wire [31:0] eq_60_in0;
	wire [31:0] eq_60_in1;
	wire [0:0] eq_60_out;
	eq #(.WIDTH(32)) eq_60(.in0(eq_60_in0), .in1(eq_60_in1), .out(eq_60_out));

	wire [0:0] orOp_61_in0;
	wire [0:0] orOp_61_in1;
	wire [0:0] orOp_61_out;
	orOp #(.WIDTH(1)) orOp_61(.in0(orOp_61_in0), .in1(orOp_61_in1), .out(orOp_61_out));

	wire [31:0] eq_62_in0;
	wire [31:0] eq_62_in1;
	wire [0:0] eq_62_out;
	eq #(.WIDTH(32)) eq_62(.in0(eq_62_in0), .in1(eq_62_in1), .out(eq_62_out));

	wire [0:0] orOp_63_in0;
	wire [0:0] orOp_63_in1;
	wire [0:0] orOp_63_out;
	orOp #(.WIDTH(1)) orOp_63(.in0(orOp_63_in0), .in1(orOp_63_in1), .out(orOp_63_out));

	wire [31:0] eq_64_in0;
	wire [31:0] eq_64_in1;
	wire [0:0] eq_64_out;
	eq #(.WIDTH(32)) eq_64(.in0(eq_64_in0), .in1(eq_64_in1), .out(eq_64_out));

	wire [0:0] orOp_65_in0;
	wire [0:0] orOp_65_in1;
	wire [0:0] orOp_65_out;
	orOp #(.WIDTH(1)) orOp_65(.in0(orOp_65_in0), .in1(orOp_65_in1), .out(orOp_65_out));

	wire [31:0] eq_66_in0;
	wire [31:0] eq_66_in1;
	wire [0:0] eq_66_out;
	eq #(.WIDTH(32)) eq_66(.in0(eq_66_in0), .in1(eq_66_in1), .out(eq_66_out));

	wire [31:0] eq_67_in0;
	wire [31:0] eq_67_in1;
	wire [0:0] eq_67_out;
	eq #(.WIDTH(32)) eq_67(.in0(eq_67_in0), .in1(eq_67_in1), .out(eq_67_out));

	wire [0:0] orOp_68_in0;
	wire [0:0] orOp_68_in1;
	wire [0:0] orOp_68_out;
	orOp #(.WIDTH(1)) orOp_68(.in0(orOp_68_in0), .in1(orOp_68_in1), .out(orOp_68_out));

	wire [31:0] eq_69_in0;
	wire [31:0] eq_69_in1;
	wire [0:0] eq_69_out;
	eq #(.WIDTH(32)) eq_69(.in0(eq_69_in0), .in1(eq_69_in1), .out(eq_69_out));

	wire [31:0] eq_70_in0;
	wire [31:0] eq_70_in1;
	wire [0:0] eq_70_out;
	eq #(.WIDTH(32)) eq_70(.in0(eq_70_in0), .in1(eq_70_in1), .out(eq_70_out));

	wire [31:0] eq_71_in0;
	wire [31:0] eq_71_in1;
	wire [0:0] eq_71_out;
	eq #(.WIDTH(32)) eq_71(.in0(eq_71_in0), .in1(eq_71_in1), .out(eq_71_out));

	wire [0:0] orOp_72_in0;
	wire [0:0] orOp_72_in1;
	wire [0:0] orOp_72_out;
	orOp #(.WIDTH(1)) orOp_72(.in0(orOp_72_in0), .in1(orOp_72_in1), .out(orOp_72_out));

	wire [31:0] eq_73_in0;
	wire [31:0] eq_73_in1;
	wire [0:0] eq_73_out;
	eq #(.WIDTH(32)) eq_73(.in0(eq_73_in0), .in1(eq_73_in1), .out(eq_73_out));

	wire [0:0] orOp_74_in0;
	wire [0:0] orOp_74_in1;
	wire [0:0] orOp_74_out;
	orOp #(.WIDTH(1)) orOp_74(.in0(orOp_74_in0), .in1(orOp_74_in1), .out(orOp_74_out));

	wire [31:0] eq_75_in0;
	wire [31:0] eq_75_in1;
	wire [0:0] eq_75_out;
	eq #(.WIDTH(32)) eq_75(.in0(eq_75_in0), .in1(eq_75_in1), .out(eq_75_out));

	wire [0:0] orOp_76_in0;
	wire [0:0] orOp_76_in1;
	wire [0:0] orOp_76_out;
	orOp #(.WIDTH(1)) orOp_76(.in0(orOp_76_in0), .in1(orOp_76_in1), .out(orOp_76_out));

	wire [31:0] eq_77_in0;
	wire [31:0] eq_77_in1;
	wire [0:0] eq_77_out;
	eq #(.WIDTH(32)) eq_77(.in0(eq_77_in0), .in1(eq_77_in1), .out(eq_77_out));

	wire [0:0] orOp_78_in0;
	wire [0:0] orOp_78_in1;
	wire [0:0] orOp_78_out;
	orOp #(.WIDTH(1)) orOp_78(.in0(orOp_78_in0), .in1(orOp_78_in1), .out(orOp_78_out));

	wire [31:0] eq_79_in0;
	wire [31:0] eq_79_in1;
	wire [0:0] eq_79_out;
	eq #(.WIDTH(32)) eq_79(.in0(eq_79_in0), .in1(eq_79_in1), .out(eq_79_out));

	wire [0:0] orOp_80_in0;
	wire [0:0] orOp_80_in1;
	wire [0:0] orOp_80_out;
	orOp #(.WIDTH(1)) orOp_80(.in0(orOp_80_in0), .in1(orOp_80_in1), .out(orOp_80_out));

	wire [31:0] eq_81_in0;
	wire [31:0] eq_81_in1;
	wire [0:0] eq_81_out;
	eq #(.WIDTH(32)) eq_81(.in0(eq_81_in0), .in1(eq_81_in1), .out(eq_81_out));

	wire [31:0] eq_82_in0;
	wire [31:0] eq_82_in1;
	wire [0:0] eq_82_out;
	eq #(.WIDTH(32)) eq_82(.in0(eq_82_in0), .in1(eq_82_in1), .out(eq_82_out));

	wire [31:0] eq_83_in0;
	wire [31:0] eq_83_in1;
	wire [0:0] eq_83_out;
	eq #(.WIDTH(32)) eq_83(.in0(eq_83_in0), .in1(eq_83_in1), .out(eq_83_out));

	wire [0:0] notOp_84_in0;
	wire [0:0] notOp_84_out;
	notOp #(.WIDTH(1)) notOp_84(.in(notOp_84_in0), .out(notOp_84_out));

	wire [0:0] andOp_85_in0;
	wire [0:0] andOp_85_in1;
	wire [0:0] andOp_85_out;
	andOp #(.WIDTH(1)) andOp_85(.in0(andOp_85_in0), .in1(andOp_85_in1), .out(andOp_85_out));

	wire [31:0] eq_86_in0;
	wire [31:0] eq_86_in1;
	wire [0:0] eq_86_out;
	eq #(.WIDTH(32)) eq_86(.in0(eq_86_in0), .in1(eq_86_in1), .out(eq_86_out));

	wire [0:0] notOp_87_in0;
	wire [0:0] notOp_87_out;
	notOp #(.WIDTH(1)) notOp_87(.in(notOp_87_in0), .out(notOp_87_out));

	wire [0:0] andOp_88_in0;
	wire [0:0] andOp_88_in1;
	wire [0:0] andOp_88_out;
	andOp #(.WIDTH(1)) andOp_88(.in0(andOp_88_in0), .in1(andOp_88_in1), .out(andOp_88_out));

	wire [31:0] eq_89_in0;
	wire [31:0] eq_89_in1;
	wire [0:0] eq_89_out;
	eq #(.WIDTH(32)) eq_89(.in0(eq_89_in0), .in1(eq_89_in1), .out(eq_89_out));

	wire [0:0] notOp_90_in0;
	wire [0:0] notOp_90_out;
	notOp #(.WIDTH(1)) notOp_90(.in(notOp_90_in0), .out(notOp_90_out));

	wire [0:0] andOp_91_in0;
	wire [0:0] andOp_91_in1;
	wire [0:0] andOp_91_out;
	andOp #(.WIDTH(1)) andOp_91(.in0(andOp_91_in0), .in1(andOp_91_in1), .out(andOp_91_out));

	wire [31:0] eq_92_in0;
	wire [31:0] eq_92_in1;
	wire [0:0] eq_92_out;
	eq #(.WIDTH(32)) eq_92(.in0(eq_92_in0), .in1(eq_92_in1), .out(eq_92_out));

	wire [31:0] eq_93_in0;
	wire [31:0] eq_93_in1;
	wire [0:0] eq_93_out;
	eq #(.WIDTH(32)) eq_93(.in0(eq_93_in0), .in1(eq_93_in1), .out(eq_93_out));

	wire [0:0] notOp_94_in0;
	wire [0:0] notOp_94_out;
	notOp #(.WIDTH(1)) notOp_94(.in(notOp_94_in0), .out(notOp_94_out));

	wire [0:0] andOp_95_in0;
	wire [0:0] andOp_95_in1;
	wire [0:0] andOp_95_out;
	andOp #(.WIDTH(1)) andOp_95(.in0(andOp_95_in0), .in1(andOp_95_in1), .out(andOp_95_out));

	wire [31:0] eq_96_in0;
	wire [31:0] eq_96_in1;
	wire [0:0] eq_96_out;
	eq #(.WIDTH(32)) eq_96(.in0(eq_96_in0), .in1(eq_96_in1), .out(eq_96_out));

	wire [31:0] eq_97_in0;
	wire [31:0] eq_97_in1;
	wire [0:0] eq_97_out;
	eq #(.WIDTH(32)) eq_97(.in0(eq_97_in0), .in1(eq_97_in1), .out(eq_97_out));

	wire [31:0] eq_98_in0;
	wire [31:0] eq_98_in1;
	wire [0:0] eq_98_out;
	eq #(.WIDTH(32)) eq_98(.in0(eq_98_in0), .in1(eq_98_in1), .out(eq_98_out));

	wire [0:0] notOp_99_in0;
	wire [0:0] notOp_99_out;
	notOp #(.WIDTH(1)) notOp_99(.in(notOp_99_in0), .out(notOp_99_out));

	wire [0:0] andOp_100_in0;
	wire [0:0] andOp_100_in1;
	wire [0:0] andOp_100_out;
	andOp #(.WIDTH(1)) andOp_100(.in0(andOp_100_in0), .in1(andOp_100_in1), .out(andOp_100_out));

	wire [31:0] eq_101_in0;
	wire [31:0] eq_101_in1;
	wire [0:0] eq_101_out;
	eq #(.WIDTH(32)) eq_101(.in0(eq_101_in0), .in1(eq_101_in1), .out(eq_101_out));

	wire [0:0] notOp_102_in0;
	wire [0:0] notOp_102_out;
	notOp #(.WIDTH(1)) notOp_102(.in(notOp_102_in0), .out(notOp_102_out));

	wire [0:0] andOp_103_in0;
	wire [0:0] andOp_103_in1;
	wire [0:0] andOp_103_out;
	andOp #(.WIDTH(1)) andOp_103(.in0(andOp_103_in0), .in1(andOp_103_in1), .out(andOp_103_out));

	wire [31:0] eq_104_in0;
	wire [31:0] eq_104_in1;
	wire [0:0] eq_104_out;
	eq #(.WIDTH(32)) eq_104(.in0(eq_104_in0), .in1(eq_104_in1), .out(eq_104_out));

	wire [0:0] notOp_105_in0;
	wire [0:0] notOp_105_out;
	notOp #(.WIDTH(1)) notOp_105(.in(notOp_105_in0), .out(notOp_105_out));

	wire [0:0] andOp_106_in0;
	wire [0:0] andOp_106_in1;
	wire [0:0] andOp_106_out;
	andOp #(.WIDTH(1)) andOp_106(.in0(andOp_106_in0), .in1(andOp_106_in1), .out(andOp_106_out));

	wire [31:0] eq_107_in0;
	wire [31:0] eq_107_in1;
	wire [0:0] eq_107_out;
	eq #(.WIDTH(32)) eq_107(.in0(eq_107_in0), .in1(eq_107_in1), .out(eq_107_out));

	wire [0:0] notOp_108_in0;
	wire [0:0] notOp_108_out;
	notOp #(.WIDTH(1)) notOp_108(.in(notOp_108_in0), .out(notOp_108_out));

	wire [0:0] andOp_109_in0;
	wire [0:0] andOp_109_in1;
	wire [0:0] andOp_109_out;
	andOp #(.WIDTH(1)) andOp_109(.in0(andOp_109_in0), .in1(andOp_109_in1), .out(andOp_109_out));

	wire [31:0] eq_110_in0;
	wire [31:0] eq_110_in1;
	wire [0:0] eq_110_out;
	eq #(.WIDTH(32)) eq_110(.in0(eq_110_in0), .in1(eq_110_in1), .out(eq_110_out));

	wire [0:0] notOp_111_in0;
	wire [0:0] notOp_111_out;
	notOp #(.WIDTH(1)) notOp_111(.in(notOp_111_in0), .out(notOp_111_out));

	wire [0:0] andOp_112_in0;
	wire [0:0] andOp_112_in1;
	wire [0:0] andOp_112_out;
	andOp #(.WIDTH(1)) andOp_112(.in0(andOp_112_in0), .in1(andOp_112_in1), .out(andOp_112_out));

	wire [0:0] andOp_113_in0;
	wire [0:0] andOp_113_in1;
	wire [0:0] andOp_113_out;
	andOp #(.WIDTH(1)) andOp_113(.in0(andOp_113_in0), .in1(andOp_113_in1), .out(andOp_113_out));

	wire [0:0] andOp_114_in0;
	wire [0:0] andOp_114_in1;
	wire [0:0] andOp_114_out;
	andOp #(.WIDTH(1)) andOp_114(.in0(andOp_114_in0), .in1(andOp_114_in1), .out(andOp_114_out));

	wire [0:0] andOp_115_in0;
	wire [0:0] andOp_115_in1;
	wire [0:0] andOp_115_out;
	andOp #(.WIDTH(1)) andOp_115(.in0(andOp_115_in0), .in1(andOp_115_in1), .out(andOp_115_out));

	wire [0:0] andOp_116_in0;
	wire [0:0] andOp_116_in1;
	wire [0:0] andOp_116_out;
	andOp #(.WIDTH(1)) andOp_116(.in0(andOp_116_in0), .in1(andOp_116_in1), .out(andOp_116_out));

	wire [0:0] andOp_117_in0;
	wire [0:0] andOp_117_in1;
	wire [0:0] andOp_117_out;
	andOp #(.WIDTH(1)) andOp_117(.in0(andOp_117_in0), .in1(andOp_117_in1), .out(andOp_117_out));

	wire [0:0] andOp_118_in0;
	wire [0:0] andOp_118_in1;
	wire [0:0] andOp_118_out;
	andOp #(.WIDTH(1)) andOp_118(.in0(andOp_118_in0), .in1(andOp_118_in1), .out(andOp_118_out));

	wire [0:0] andOp_119_in0;
	wire [0:0] andOp_119_in1;
	wire [0:0] andOp_119_out;
	andOp #(.WIDTH(1)) andOp_119(.in0(andOp_119_in0), .in1(andOp_119_in1), .out(andOp_119_out));

	wire [0:0] andOp_120_in0;
	wire [0:0] andOp_120_in1;
	wire [0:0] andOp_120_out;
	andOp #(.WIDTH(1)) andOp_120(.in0(andOp_120_in0), .in1(andOp_120_in1), .out(andOp_120_out));

	wire [31:0] concat_121_in0;
	wire [31:0] concat_121_in1;
	wire [63:0] concat_121_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_121(.in0(concat_121_in0), .in1(concat_121_in1), .out(concat_121_out));

	wire [31:0] concat_122_in0;
	wire [31:0] concat_122_in1;
	wire [63:0] concat_122_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_122(.in0(concat_122_in0), .in1(concat_122_in1), .out(concat_122_out));

	wire [0:0] andOp_123_in0;
	wire [0:0] andOp_123_in1;
	wire [0:0] andOp_123_out;
	andOp #(.WIDTH(1)) andOp_123(.in0(andOp_123_in0), .in1(andOp_123_in1), .out(andOp_123_out));

	wire [0:0] andOp_124_in0;
	wire [0:0] andOp_124_in1;
	wire [0:0] andOp_124_out;
	andOp #(.WIDTH(1)) andOp_124(.in0(andOp_124_in0), .in1(andOp_124_in1), .out(andOp_124_out));

	wire [0:0] andOp_125_in0;
	wire [0:0] andOp_125_in1;
	wire [0:0] andOp_125_out;
	andOp #(.WIDTH(1)) andOp_125(.in0(andOp_125_in0), .in1(andOp_125_in1), .out(andOp_125_out));

	wire [0:0] andOp_126_in0;
	wire [0:0] andOp_126_in1;
	wire [0:0] andOp_126_out;
	andOp #(.WIDTH(1)) andOp_126(.in0(andOp_126_in0), .in1(andOp_126_in1), .out(andOp_126_out));

	reg [31:0] tmp_output_127_in_data;
	wire [31:0] tmp_output_127_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_127(.in_data(tmp_output_127_in_data), .out_data(tmp_output_127_out_data));

	wire [31:0] eq_128_in0;
	wire [31:0] eq_128_in1;
	wire [0:0] eq_128_out;
	eq #(.WIDTH(32)) eq_128(.in0(eq_128_in0), .in1(eq_128_in1), .out(eq_128_out));

	wire [0:0] andOp_129_in0;
	wire [0:0] andOp_129_in1;
	wire [0:0] andOp_129_out;
	andOp #(.WIDTH(1)) andOp_129(.in0(andOp_129_in0), .in1(andOp_129_in1), .out(andOp_129_out));

	wire [0:0] andOp_130_in0;
	wire [0:0] andOp_130_in1;
	wire [0:0] andOp_130_out;
	andOp #(.WIDTH(1)) andOp_130(.in0(andOp_130_in0), .in1(andOp_130_in1), .out(andOp_130_out));

	wire [0:0] andOp_131_in0;
	wire [0:0] andOp_131_in1;
	wire [0:0] andOp_131_out;
	andOp #(.WIDTH(1)) andOp_131(.in0(andOp_131_in0), .in1(andOp_131_in1), .out(andOp_131_out));

	wire [0:0] andOp_132_in0;
	wire [0:0] andOp_132_in1;
	wire [0:0] andOp_132_out;
	andOp #(.WIDTH(1)) andOp_132(.in0(andOp_132_in0), .in1(andOp_132_in1), .out(andOp_132_out));

	wire [0:0] andOp_133_in0;
	wire [0:0] andOp_133_in1;
	wire [0:0] andOp_133_out;
	andOp #(.WIDTH(1)) andOp_133(.in0(andOp_133_in0), .in1(andOp_133_in1), .out(andOp_133_out));

	wire [0:0] andOp_134_in0;
	wire [0:0] andOp_134_in1;
	wire [0:0] andOp_134_out;
	andOp #(.WIDTH(1)) andOp_134(.in0(andOp_134_in0), .in1(andOp_134_in1), .out(andOp_134_out));

	wire [0:0] andOp_135_in0;
	wire [0:0] andOp_135_in1;
	wire [0:0] andOp_135_out;
	andOp #(.WIDTH(1)) andOp_135(.in0(andOp_135_in0), .in1(andOp_135_in1), .out(andOp_135_out));

	wire [0:0] andOp_136_in0;
	wire [0:0] andOp_136_in1;
	wire [0:0] andOp_136_out;
	andOp #(.WIDTH(1)) andOp_136(.in0(andOp_136_in0), .in1(andOp_136_in1), .out(andOp_136_out));

	wire [0:0] andOp_137_in0;
	wire [0:0] andOp_137_in1;
	wire [0:0] andOp_137_out;
	andOp #(.WIDTH(1)) andOp_137(.in0(andOp_137_in0), .in1(andOp_137_in1), .out(andOp_137_out));

	wire [0:0] andOp_138_in0;
	wire [0:0] andOp_138_in1;
	wire [0:0] andOp_138_out;
	andOp #(.WIDTH(1)) andOp_138(.in0(andOp_138_in0), .in1(andOp_138_in1), .out(andOp_138_out));

	wire [0:0] andOp_139_in0;
	wire [0:0] andOp_139_in1;
	wire [0:0] andOp_139_out;
	andOp #(.WIDTH(1)) andOp_139(.in0(andOp_139_in0), .in1(andOp_139_in1), .out(andOp_139_out));

	wire [0:0] notOp_140_in0;
	wire [0:0] notOp_140_out;
	notOp #(.WIDTH(1)) notOp_140(.in(notOp_140_in0), .out(notOp_140_out));

	wire [0:0] andOp_141_in0;
	wire [0:0] andOp_141_in1;
	wire [0:0] andOp_141_out;
	andOp #(.WIDTH(1)) andOp_141(.in0(andOp_141_in0), .in1(andOp_141_in1), .out(andOp_141_out));

	wire [0:0] notOp_142_in0;
	wire [0:0] notOp_142_out;
	notOp #(.WIDTH(1)) notOp_142(.in(notOp_142_in0), .out(notOp_142_out));

	wire [0:0] andOp_143_in0;
	wire [0:0] andOp_143_in1;
	wire [0:0] andOp_143_out;
	andOp #(.WIDTH(1)) andOp_143(.in0(andOp_143_in0), .in1(andOp_143_in1), .out(andOp_143_out));

	wire [0:0] notOp_144_in0;
	wire [0:0] notOp_144_out;
	notOp #(.WIDTH(1)) notOp_144(.in(notOp_144_in0), .out(notOp_144_out));

	wire [0:0] andOp_145_in0;
	wire [0:0] andOp_145_in1;
	wire [0:0] andOp_145_out;
	andOp #(.WIDTH(1)) andOp_145(.in0(andOp_145_in0), .in1(andOp_145_in1), .out(andOp_145_out));

	wire [0:0] notOp_146_in0;
	wire [0:0] notOp_146_out;
	notOp #(.WIDTH(1)) notOp_146(.in(notOp_146_in0), .out(notOp_146_out));

	wire [0:0] andOp_147_in0;
	wire [0:0] andOp_147_in1;
	wire [0:0] andOp_147_out;
	andOp #(.WIDTH(1)) andOp_147(.in0(andOp_147_in0), .in1(andOp_147_in1), .out(andOp_147_out));

	wire [0:0] notOp_148_in0;
	wire [0:0] notOp_148_out;
	notOp #(.WIDTH(1)) notOp_148(.in(notOp_148_in0), .out(notOp_148_out));

	wire [0:0] andOp_149_in0;
	wire [0:0] andOp_149_in1;
	wire [0:0] andOp_149_out;
	andOp #(.WIDTH(1)) andOp_149(.in0(andOp_149_in0), .in1(andOp_149_in1), .out(andOp_149_out));

	wire [0:0] notOp_150_in0;
	wire [0:0] notOp_150_out;
	notOp #(.WIDTH(1)) notOp_150(.in(notOp_150_in0), .out(notOp_150_out));

	wire [0:0] andOp_151_in0;
	wire [0:0] andOp_151_in1;
	wire [0:0] andOp_151_out;
	andOp #(.WIDTH(1)) andOp_151(.in0(andOp_151_in0), .in1(andOp_151_in1), .out(andOp_151_out));

	wire [0:0] notOp_152_in0;
	wire [0:0] notOp_152_out;
	notOp #(.WIDTH(1)) notOp_152(.in(notOp_152_in0), .out(notOp_152_out));

	wire [0:0] andOp_153_in0;
	wire [0:0] andOp_153_in1;
	wire [0:0] andOp_153_out;
	andOp #(.WIDTH(1)) andOp_153(.in0(andOp_153_in0), .in1(andOp_153_in1), .out(andOp_153_out));

	wire [0:0] notOp_154_in0;
	wire [0:0] notOp_154_out;
	notOp #(.WIDTH(1)) notOp_154(.in(notOp_154_in0), .out(notOp_154_out));

	wire [0:0] andOp_155_in0;
	wire [0:0] andOp_155_in1;
	wire [0:0] andOp_155_out;
	andOp #(.WIDTH(1)) andOp_155(.in0(andOp_155_in0), .in1(andOp_155_in1), .out(andOp_155_out));

	wire [31:0] eq_156_in0;
	wire [31:0] eq_156_in1;
	wire [0:0] eq_156_out;
	eq #(.WIDTH(32)) eq_156(.in0(eq_156_in0), .in1(eq_156_in1), .out(eq_156_out));

	wire [31:0] eq_157_in0;
	wire [31:0] eq_157_in1;
	wire [0:0] eq_157_out;
	eq #(.WIDTH(32)) eq_157(.in0(eq_157_in0), .in1(eq_157_in1), .out(eq_157_out));

	wire [31:0] eq_158_in0;
	wire [31:0] eq_158_in1;
	wire [0:0] eq_158_out;
	eq #(.WIDTH(32)) eq_158(.in0(eq_158_in0), .in1(eq_158_in1), .out(eq_158_out));

	wire [31:0] eq_159_in0;
	wire [31:0] eq_159_in1;
	wire [0:0] eq_159_out;
	eq #(.WIDTH(32)) eq_159(.in0(eq_159_in0), .in1(eq_159_in1), .out(eq_159_out));

	wire [0:0] andOp_160_in0;
	wire [0:0] andOp_160_in1;
	wire [0:0] andOp_160_out;
	andOp #(.WIDTH(1)) andOp_160(.in0(andOp_160_in0), .in1(andOp_160_in1), .out(andOp_160_out));

	wire [31:0] eq_161_in0;
	wire [31:0] eq_161_in1;
	wire [0:0] eq_161_out;
	eq #(.WIDTH(32)) eq_161(.in0(eq_161_in0), .in1(eq_161_in1), .out(eq_161_out));

	wire [31:0] eq_162_in0;
	wire [31:0] eq_162_in1;
	wire [0:0] eq_162_out;
	eq #(.WIDTH(32)) eq_162(.in0(eq_162_in0), .in1(eq_162_in1), .out(eq_162_out));

	wire [31:0] eq_163_in0;
	wire [31:0] eq_163_in1;
	wire [0:0] eq_163_out;
	eq #(.WIDTH(32)) eq_163(.in0(eq_163_in0), .in1(eq_163_in1), .out(eq_163_out));

	wire [31:0] eq_164_in0;
	wire [31:0] eq_164_in1;
	wire [0:0] eq_164_out;
	eq #(.WIDTH(32)) eq_164(.in0(eq_164_in0), .in1(eq_164_in1), .out(eq_164_out));

	wire [0:0] andOp_165_in0;
	wire [0:0] andOp_165_in1;
	wire [0:0] andOp_165_out;
	andOp #(.WIDTH(1)) andOp_165(.in0(andOp_165_in0), .in1(andOp_165_in1), .out(andOp_165_out));

	wire [0:0] andOp_166_in0;
	wire [0:0] andOp_166_in1;
	wire [0:0] andOp_166_out;
	andOp #(.WIDTH(1)) andOp_166(.in0(andOp_166_in0), .in1(andOp_166_in1), .out(andOp_166_out));

	wire [31:0] eq_167_in0;
	wire [31:0] eq_167_in1;
	wire [0:0] eq_167_out;
	eq #(.WIDTH(32)) eq_167(.in0(eq_167_in0), .in1(eq_167_in1), .out(eq_167_out));

	wire [31:0] eq_168_in0;
	wire [31:0] eq_168_in1;
	wire [0:0] eq_168_out;
	eq #(.WIDTH(32)) eq_168(.in0(eq_168_in0), .in1(eq_168_in1), .out(eq_168_out));

	// End Functional Units

	reg [31:0] data_store_0_0;
	reg [31:0] data_store_0_2;
	reg [31:0] data_store_1_4;
	reg [31:0] data_store_1_6;
	reg [31:0] data_store_2_8;
	reg [31:0] data_store_3_10;
	reg [0:0] data_store_3_11;
	reg [31:0] data_store_3_12;
	reg [31:0] data_store_4_14;
	reg [0:0] data_store_4_16;
	reg [31:0] data_store_4_18;
	reg [31:0] global_state;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_3_last_state;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;
	reg [31:0] state_4_last_state;

	// controller for add_add13.add_add13_in0
	// controller for add_add13.add_add13_in1
	// Insensitive connections
	assign add_add13_in0 = rdata_ram_0;
	assign add_add13_in1 = tmp_output_127_out_data;
	// controller for add_add15.add_add15_in0
	// controller for add_add15.add_add15_in1
	// Insensitive connections
	assign add_add15_in0 = data_in_3_13_out_data;
	assign add_add15_in1 = 32'd1;
	// controller for andOp_100.andOp_100_in0
	// controller for andOp_100.andOp_100_in1
	// Insensitive connections
	assign andOp_100_in0 = notOp_99_out;
	assign andOp_100_in1 = andOp_52_out;
	// controller for andOp_103.andOp_103_in0
	// controller for andOp_103.andOp_103_in1
	// Insensitive connections
	assign andOp_103_in0 = notOp_102_out;
	assign andOp_103_in1 = andOp_54_out;
	// controller for andOp_106.andOp_106_in0
	// controller for andOp_106.andOp_106_in1
	// Insensitive connections
	assign andOp_106_in0 = notOp_105_out;
	assign andOp_106_in1 = andOp_56_out;
	// controller for andOp_109.andOp_109_in0
	// controller for andOp_109.andOp_109_in1
	// Insensitive connections
	assign andOp_109_in0 = notOp_108_out;
	assign andOp_109_in1 = andOp_49_out;
	// controller for andOp_112.andOp_112_in0
	// controller for andOp_112.andOp_112_in1
	// Insensitive connections
	assign andOp_112_in0 = notOp_111_out;
	assign andOp_112_in1 = andOp_37_out;
	// controller for andOp_113.andOp_113_in0
	// controller for andOp_113.andOp_113_in1
	// Insensitive connections
	assign andOp_113_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_113_in1 = state_0_is_active;
	// controller for andOp_114.andOp_114_in0
	// controller for andOp_114.andOp_114_in1
	// Insensitive connections
	assign andOp_114_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_114_in1 = state_0_is_active;
	// controller for andOp_115.andOp_115_in0
	// controller for andOp_115.andOp_115_in1
	// Insensitive connections
	assign andOp_115_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_115_in1 = state_0_is_active;
	// controller for andOp_116.andOp_116_in0
	// controller for andOp_116.andOp_116_in1
	// Insensitive connections
	assign andOp_116_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_116_in1 = state_0_is_active;
	// controller for andOp_117.andOp_117_in0
	// controller for andOp_117.andOp_117_in1
	// Insensitive connections
	assign andOp_117_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_117_in1 = state_3_is_active;
	// controller for andOp_118.andOp_118_in0
	// controller for andOp_118.andOp_118_in1
	// Insensitive connections
	assign andOp_118_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_118_in1 = state_3_is_active;
	// controller for andOp_119.andOp_119_in0
	// controller for andOp_119.andOp_119_in1
	// Insensitive connections
	assign andOp_119_in0 = bb_7_active_in_state_4_out_data;
	assign andOp_119_in1 = state_4_is_active;
	// controller for andOp_120.andOp_120_in0
	// controller for andOp_120.andOp_120_in1
	// Insensitive connections
	assign andOp_120_in0 = bb_3_active_in_state_1_out_data;
	assign andOp_120_in1 = state_1_is_active;
	// controller for andOp_123.andOp_123_in0
	// controller for andOp_123.andOp_123_in1
	// Insensitive connections
	assign andOp_123_in0 = bb_9_active_in_state_1_out_data;
	assign andOp_123_in1 = state_1_is_active;
	// controller for andOp_124.andOp_124_in0
	// controller for andOp_124.andOp_124_in1
	// Insensitive connections
	assign andOp_124_in0 = bb_10_active_in_state_2_out_data;
	assign andOp_124_in1 = state_2_is_active;
	// controller for andOp_125.andOp_125_in0
	// controller for andOp_125.andOp_125_in1
	// Insensitive connections
	assign andOp_125_in0 = bb_10_active_in_state_3_out_data;
	assign andOp_125_in1 = state_3_is_active;
	// controller for andOp_126.andOp_126_in0
	// controller for andOp_126.andOp_126_in1
	// Insensitive connections
	assign andOp_126_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_126_in1 = state_3_is_active;
	// controller for andOp_129.andOp_129_in0
	// controller for andOp_129.andOp_129_in1
	// Insensitive connections
	assign andOp_129_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_129_in1 = state_3_is_active;
	// controller for andOp_130.andOp_130_in0
	// controller for andOp_130.andOp_130_in1
	// Insensitive connections
	assign andOp_130_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_130_in1 = state_3_is_active;
	// controller for andOp_131.andOp_131_in0
	// controller for andOp_131.andOp_131_in1
	// Insensitive connections
	assign andOp_131_in0 = bb_6_active_in_state_4_out_data;
	assign andOp_131_in1 = state_4_is_active;
	// controller for andOp_132.andOp_132_in0
	// controller for andOp_132.andOp_132_in1
	// Insensitive connections
	assign andOp_132_in0 = bb_7_active_in_state_4_out_data;
	assign andOp_132_in1 = state_4_is_active;
	// controller for andOp_133.andOp_133_in0
	// controller for andOp_133.andOp_133_in1
	// Insensitive connections
	assign andOp_133_in0 = bb_7_active_in_state_4_out_data;
	assign andOp_133_in1 = state_4_is_active;
	// controller for andOp_134.andOp_134_in0
	// controller for andOp_134.andOp_134_in1
	// Insensitive connections
	assign andOp_134_in0 = bb_2_active_in_state_4_out_data;
	assign andOp_134_in1 = state_4_is_active;
	// controller for andOp_135.andOp_135_in0
	// controller for andOp_135.andOp_135_in1
	// Insensitive connections
	assign andOp_135_in0 = bb_2_active_in_state_4_out_data;
	assign andOp_135_in1 = state_4_is_active;
	// controller for andOp_136.andOp_136_in0
	// controller for andOp_136.andOp_136_in1
	// Insensitive connections
	assign andOp_136_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_136_in1 = state_0_is_active;
	// controller for andOp_137.andOp_137_in0
	// controller for andOp_137.andOp_137_in1
	// Insensitive connections
	assign andOp_137_in0 = bb_10_active_in_state_2_out_data;
	assign andOp_137_in1 = state_2_is_active;
	// controller for andOp_138.andOp_138_in0
	// controller for andOp_138.andOp_138_in1
	// Insensitive connections
	assign andOp_138_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_138_in1 = state_3_is_active;
	// controller for andOp_139.andOp_139_in0
	// controller for andOp_139.andOp_139_in1
	// Insensitive connections
	assign andOp_139_in0 = bb_2_active_in_state_4_out_data;
	assign andOp_139_in1 = state_4_is_active;
	// controller for andOp_141.andOp_141_in0
	// controller for andOp_141.andOp_141_in1
	// Insensitive connections
	assign andOp_141_in0 = notOp_140_out;
	assign andOp_141_in1 = 1'd1;
	// controller for andOp_143.andOp_143_in0
	// controller for andOp_143.andOp_143_in1
	// Insensitive connections
	assign andOp_143_in0 = notOp_142_out;
	assign andOp_143_in1 = andOp_141_out;
	// controller for andOp_145.andOp_145_in0
	// controller for andOp_145.andOp_145_in1
	// Insensitive connections
	assign andOp_145_in0 = notOp_144_out;
	assign andOp_145_in1 = andOp_143_out;
	// controller for andOp_147.andOp_147_in0
	// controller for andOp_147.andOp_147_in1
	// Insensitive connections
	assign andOp_147_in0 = notOp_146_out;
	assign andOp_147_in1 = 1'd1;
	// controller for andOp_149.andOp_149_in0
	// controller for andOp_149.andOp_149_in1
	// Insensitive connections
	assign andOp_149_in0 = notOp_148_out;
	assign andOp_149_in1 = 1'd1;
	// controller for andOp_151.andOp_151_in0
	// controller for andOp_151.andOp_151_in1
	// Insensitive connections
	assign andOp_151_in0 = notOp_150_out;
	assign andOp_151_in1 = 1'd1;
	// controller for andOp_153.andOp_153_in0
	// controller for andOp_153.andOp_153_in1
	// Insensitive connections
	assign andOp_153_in0 = notOp_152_out;
	assign andOp_153_in1 = andOp_151_out;
	// controller for andOp_155.andOp_155_in0
	// controller for andOp_155.andOp_155_in1
	// Insensitive connections
	assign andOp_155_in0 = notOp_154_out;
	assign andOp_155_in1 = andOp_153_out;
	// controller for andOp_160.andOp_160_in0
	// controller for andOp_160.andOp_160_in1
	// Insensitive connections
	assign andOp_160_in0 = bb_3_active_in_state_1_out_data;
	assign andOp_160_in1 = state_1_is_active;
	// controller for andOp_165.andOp_165_in0
	// controller for andOp_165.andOp_165_in1
	// Insensitive connections
	assign andOp_165_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_165_in1 = state_3_is_active;
	// controller for andOp_166.andOp_166_in0
	// controller for andOp_166.andOp_166_in1
	// Insensitive connections
	assign andOp_166_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_166_in1 = state_3_is_active;
	// controller for andOp_20.andOp_20_in0
	// controller for andOp_20.andOp_20_in1
	// Insensitive connections
	assign andOp_20_in0 = bb_0_active_in_state_1_out_data;
	assign andOp_20_in1 = state_1_is_active;
	// controller for andOp_22.andOp_22_in0
	// controller for andOp_22.andOp_22_in1
	// Insensitive connections
	assign andOp_22_in0 = bb_0_active_in_state_1_out_data;
	assign andOp_22_in1 = state_1_is_active;
	// controller for andOp_24.andOp_24_in0
	// controller for andOp_24.andOp_24_in1
	// Insensitive connections
	assign andOp_24_in0 = bb_8_active_in_state_1_out_data;
	assign andOp_24_in1 = state_1_is_active;
	// controller for andOp_26.andOp_26_in0
	// controller for andOp_26.andOp_26_in1
	// Insensitive connections
	assign andOp_26_in0 = bb_3_active_in_state_1_out_data;
	assign andOp_26_in1 = state_1_is_active;
	// controller for andOp_28.andOp_28_in0
	// controller for andOp_28.andOp_28_in1
	// Insensitive connections
	assign andOp_28_in0 = bb_9_active_in_state_1_out_data;
	assign andOp_28_in1 = state_1_is_active;
	// controller for andOp_30.andOp_30_in0
	// controller for andOp_30.andOp_30_in1
	// Insensitive connections
	assign andOp_30_in0 = andOp_28_out;
	assign andOp_30_in1 = in_read_ready;
	// controller for andOp_32.andOp_32_in0
	// controller for andOp_32.andOp_32_in1
	// Insensitive connections
	assign andOp_32_in0 = andOp_28_out;
	assign andOp_32_in1 = notOp_31_out;
	// controller for andOp_33.andOp_33_in0
	// controller for andOp_33.andOp_33_in1
	// Insensitive connections
	assign andOp_33_in0 = bb_10_active_in_state_3_out_data;
	assign andOp_33_in1 = state_3_is_active;
	// controller for andOp_35.andOp_35_in0
	// controller for andOp_35.andOp_35_in1
	// Insensitive connections
	assign andOp_35_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_35_in1 = state_4_is_active;
	// controller for andOp_37.andOp_37_in0
	// controller for andOp_37.andOp_37_in1
	// Insensitive connections
	assign andOp_37_in0 = andOp_35_out;
	assign andOp_37_in1 = data_in_4_17_out_data;
	// controller for andOp_39.andOp_39_in0
	// controller for andOp_39.andOp_39_in1
	// Insensitive connections
	assign andOp_39_in0 = andOp_35_out;
	assign andOp_39_in1 = notOp_38_out;
	// controller for andOp_40.andOp_40_in0
	// controller for andOp_40.andOp_40_in1
	// Insensitive connections
	assign andOp_40_in0 = bb_10_active_in_state_3_out_data;
	assign andOp_40_in1 = state_3_is_active;
	// controller for andOp_42.andOp_42_in0
	// controller for andOp_42.andOp_42_in1
	// Insensitive connections
	assign andOp_42_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_42_in1 = state_4_is_active;
	// controller for andOp_44.andOp_44_in0
	// controller for andOp_44.andOp_44_in1
	// Insensitive connections
	assign andOp_44_in0 = andOp_42_out;
	assign andOp_44_in1 = data_in_4_17_out_data;
	// controller for andOp_46.andOp_46_in0
	// controller for andOp_46.andOp_46_in1
	// Insensitive connections
	assign andOp_46_in0 = andOp_42_out;
	assign andOp_46_in1 = notOp_45_out;
	// controller for andOp_47.andOp_47_in0
	// controller for andOp_47.andOp_47_in1
	// Insensitive connections
	assign andOp_47_in0 = bb_6_active_in_state_4_out_data;
	assign andOp_47_in1 = state_4_is_active;
	// controller for andOp_49.andOp_49_in0
	// controller for andOp_49.andOp_49_in1
	// Insensitive connections
	assign andOp_49_in0 = andOp_47_out;
	assign andOp_49_in1 = out_write_ready;
	// controller for andOp_51.andOp_51_in0
	// controller for andOp_51.andOp_51_in1
	// Insensitive connections
	assign andOp_51_in0 = andOp_47_out;
	assign andOp_51_in1 = notOp_50_out;
	// controller for andOp_52.andOp_52_in0
	// controller for andOp_52.andOp_52_in1
	// Insensitive connections
	assign andOp_52_in0 = bb_5_active_in_state_4_out_data;
	assign andOp_52_in1 = state_4_is_active;
	// controller for andOp_54.andOp_54_in0
	// controller for andOp_54.andOp_54_in1
	// Insensitive connections
	assign andOp_54_in0 = bb_7_active_in_state_4_out_data;
	assign andOp_54_in1 = state_4_is_active;
	// controller for andOp_56.andOp_56_in0
	// controller for andOp_56.andOp_56_in1
	// Insensitive connections
	assign andOp_56_in0 = bb_1_active_in_state_4_out_data;
	assign andOp_56_in1 = state_4_is_active;
	// controller for andOp_85.andOp_85_in0
	// controller for andOp_85.andOp_85_in1
	// Insensitive connections
	assign andOp_85_in0 = notOp_84_out;
	assign andOp_85_in1 = andOp_26_out;
	// controller for andOp_88.andOp_88_in0
	// controller for andOp_88.andOp_88_in1
	// Insensitive connections
	assign andOp_88_in0 = notOp_87_out;
	assign andOp_88_in1 = andOp_20_out;
	// controller for andOp_91.andOp_91_in0
	// controller for andOp_91.andOp_91_in1
	// Insensitive connections
	assign andOp_91_in0 = notOp_90_out;
	assign andOp_91_in1 = andOp_24_out;
	// controller for andOp_95.andOp_95_in0
	// controller for andOp_95.andOp_95_in1
	// Insensitive connections
	assign andOp_95_in0 = notOp_94_out;
	assign andOp_95_in1 = andOp_33_out;
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_58_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_active_in_state_1.bb_0_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_1_in_data = eq_59_out;
		end else begin
			bb_0_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_81_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_1.bb_0_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_82_out) begin 
			bb_0_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_2.bb_10_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_2_in_data = eq_66_out;
		end else begin
			bb_10_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_3.bb_10_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_3_in_data = eq_69_out;
		end else begin
			bb_10_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_2.bb_10_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_92_out) begin 
			bb_10_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_3.bb_10_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_96_out) begin 
			bb_10_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_4.bb_1_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_4_in_data = orOp_80_out;
		end else begin
			bb_1_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_4.bb_1_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_112_out) begin 
			bb_1_predecessor_in_state_4_in_data = 32'd4;
		end else if (eq_110_out) begin 
			bb_1_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_4.bb_2_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_4_in_data = orOp_74_out;
		end else begin
			bb_2_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_4.bb_2_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_103_out) begin 
			bb_2_predecessor_in_state_4_in_data = 32'd7;
		end else if (eq_101_out) begin 
			bb_2_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_1.bb_3_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_1_in_data = orOp_63_out;
		end else begin
			bb_3_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_1.bb_3_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_88_out) begin 
			bb_3_predecessor_in_state_1_in_data = 32'd0;
		end else if (eq_86_out) begin 
			bb_3_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_3.bb_4_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_3_in_data = orOp_68_out;
		end else begin
			bb_4_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_4.bb_4_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_4_in_data = eq_70_out;
		end else begin
			bb_4_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_3.bb_4_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_95_out) begin 
			bb_4_predecessor_in_state_3_in_data = 32'd10;
		end else if (eq_93_out) begin 
			bb_4_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_4.bb_4_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_97_out) begin 
			bb_4_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_5_active_in_state_4.bb_5_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_5_active_in_state_4_in_data = orOp_76_out;
		end else begin
			bb_5_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_5_predecessor_in_state_4.bb_5_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_106_out) begin 
			bb_5_predecessor_in_state_4_in_data = 32'd1;
		end else if (eq_104_out) begin 
			bb_5_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_5_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_6_active_in_state_4.bb_6_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_6_active_in_state_4_in_data = orOp_72_out;
		end else begin
			bb_6_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_6_predecessor_in_state_4.bb_6_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_100_out) begin 
			bb_6_predecessor_in_state_4_in_data = 32'd5;
		end else if (eq_98_out) begin 
			bb_6_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_6_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_7_active_in_state_4.bb_7_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_7_active_in_state_4_in_data = orOp_78_out;
		end else begin
			bb_7_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_7_predecessor_in_state_4.bb_7_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_109_out) begin 
			bb_7_predecessor_in_state_4_in_data = 32'd6;
		end else if (eq_107_out) begin 
			bb_7_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_7_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_8_active_in_state_1.bb_8_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_state_1_in_data = orOp_61_out;
		end else begin
			bb_8_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_8_predecessor_in_state_1.bb_8_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_85_out) begin 
			bb_8_predecessor_in_state_1_in_data = 32'd3;
		end else if (eq_83_out) begin 
			bb_8_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_8_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_9_active_in_state_1.bb_9_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_9_active_in_state_1_in_data = orOp_65_out;
		end else begin
			bb_9_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_9_predecessor_in_state_1.bb_9_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_91_out) begin 
			bb_9_predecessor_in_state_1_in_data = 32'd8;
		end else if (eq_89_out) begin 
			bb_9_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_9_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_20_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_21_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_1.br_0_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_22_out) begin 
			br_0_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_23_out) begin 
			br_0_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_2.br_10_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_33_out) begin 
			br_10_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_34_out) begin 
			br_10_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_3.br_10_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_40_out) begin 
			br_10_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_41_out) begin 
			br_10_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_1_happened_in_state_4.br_1_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_56_out) begin 
			br_1_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_57_out) begin 
			br_1_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_1_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_1.br_3_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_26_out) begin 
			br_3_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_27_out) begin 
			br_3_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_3.br_4_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_35_out) begin 
			br_4_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_36_out) begin 
			br_4_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_4.br_4_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_42_out) begin 
			br_4_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_43_out) begin 
			br_4_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_5_happened_in_state_4.br_5_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_52_out) begin 
			br_5_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_53_out) begin 
			br_5_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_5_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_6_happened_in_state_4.br_6_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_47_out) begin 
			br_6_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_48_out) begin 
			br_6_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_6_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_7_happened_in_state_4.br_7_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_54_out) begin 
			br_7_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_55_out) begin 
			br_7_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_7_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_8_happened_in_state_1.br_8_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_24_out) begin 
			br_8_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_25_out) begin 
			br_8_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_8_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_9_happened_in_state_1.br_9_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_28_out) begin 
			br_9_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_29_out) begin 
			br_9_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_9_happened_in_state_1_in_data = 0;
		end
	end
	// controller for concat_121.concat_121_in0
	// controller for concat_121.concat_121_in1
	// Insensitive connections
	assign concat_121_in0 = data_in_1_5_out_data;
	assign concat_121_in1 = 32'd0;
	// controller for concat_122.concat_122_in0
	// controller for concat_122.concat_122_in1
	// Insensitive connections
	assign concat_122_in0 = 32'd4;
	assign concat_122_in1 = 32'd0;
	// controller for data_in_0_1.data_in_0_1_in_data
	always @(*) begin
		if (eq_156_out) begin 
			data_in_0_1_in_data = data_store_0_0;
		end else begin
			data_in_0_1_in_data = 0;
		end
	end
	// controller for data_in_0_3.data_in_0_3_in_data
	always @(*) begin
		if (eq_156_out) begin 
			data_in_0_3_in_data = data_store_0_2;
		end else begin
			data_in_0_3_in_data = 0;
		end
	end
	// controller for data_in_1_5.data_in_1_5_in_data
	always @(*) begin
		if (eq_157_out) begin 
			data_in_1_5_in_data = data_store_0_0;
		end else if (eq_158_out) begin 
			data_in_1_5_in_data = data_store_1_4;
		end else if (eq_159_out) begin 
			data_in_1_5_in_data = data_store_4_14;
		end else begin
			data_in_1_5_in_data = 0;
		end
	end
	// controller for data_in_1_7.data_in_1_7_in_data
	always @(*) begin
		if (eq_157_out) begin 
			data_in_1_7_in_data = data_store_0_2;
		end else if (eq_158_out) begin 
			data_in_1_7_in_data = data_store_1_6;
		end else if (eq_159_out) begin 
			data_in_1_7_in_data = data_store_4_18;
		end else begin
			data_in_1_7_in_data = 0;
		end
	end
	// controller for data_in_2_9.data_in_2_9_in_data
	always @(*) begin
		if (eq_161_out) begin 
			data_in_2_9_in_data = data_store_1_6;
		end else if (eq_162_out) begin 
			data_in_2_9_in_data = data_store_2_8;
		end else begin
			data_in_2_9_in_data = 0;
		end
	end
	// controller for data_in_3_13.data_in_3_13_in_data
	always @(*) begin
		if (eq_163_out) begin 
			data_in_3_13_in_data = data_store_2_8;
		end else if (eq_164_out) begin 
			data_in_3_13_in_data = data_store_3_12;
		end else begin
			data_in_3_13_in_data = 0;
		end
	end
	// controller for data_in_4_15.data_in_4_15_in_data
	always @(*) begin
		if (eq_167_out) begin 
			data_in_4_15_in_data = data_store_3_10;
		end else if (eq_168_out) begin 
			data_in_4_15_in_data = data_store_4_14;
		end else begin
			data_in_4_15_in_data = 0;
		end
	end
	// controller for data_in_4_17.data_in_4_17_in_data
	always @(*) begin
		if (eq_167_out) begin 
			data_in_4_17_in_data = data_store_3_11;
		end else if (eq_168_out) begin 
			data_in_4_17_in_data = data_store_4_16;
		end else begin
			data_in_4_17_in_data = 0;
		end
	end
	// controller for data_in_4_19.data_in_4_19_in_data
	always @(*) begin
		if (eq_167_out) begin 
			data_in_4_19_in_data = data_store_3_12;
		end else if (eq_168_out) begin 
			data_in_4_19_in_data = data_store_4_18;
		end else begin
			data_in_4_19_in_data = 0;
		end
	end
	// controller for eq_101.eq_101_in0
	// controller for eq_101.eq_101_in1
	// Insensitive connections
	assign eq_101_in0 = 32'd2;
	assign eq_101_in1 = state_4_entry_BB_reg;
	// controller for eq_104.eq_104_in0
	// controller for eq_104.eq_104_in1
	// Insensitive connections
	assign eq_104_in0 = 32'd5;
	assign eq_104_in1 = state_4_entry_BB_reg;
	// controller for eq_107.eq_107_in0
	// controller for eq_107.eq_107_in1
	// Insensitive connections
	assign eq_107_in0 = 32'd7;
	assign eq_107_in1 = state_4_entry_BB_reg;
	// controller for eq_110.eq_110_in0
	// controller for eq_110.eq_110_in1
	// Insensitive connections
	assign eq_110_in0 = 32'd1;
	assign eq_110_in1 = state_4_entry_BB_reg;
	// controller for eq_128.eq_128_in0
	// controller for eq_128.eq_128_in1
	// Insensitive connections
	assign eq_128_in0 = 32'd10;
	assign eq_128_in1 = state_3_entry_BB_reg;
	// controller for eq_156.eq_156_in0
	// controller for eq_156.eq_156_in1
	// Insensitive connections
	assign eq_156_in0 = 32'd0;
	assign eq_156_in1 = state_0_last_state;
	// controller for eq_157.eq_157_in0
	// controller for eq_157.eq_157_in1
	// Insensitive connections
	assign eq_157_in0 = 32'd0;
	assign eq_157_in1 = state_1_last_state;
	// controller for eq_158.eq_158_in0
	// controller for eq_158.eq_158_in1
	// Insensitive connections
	assign eq_158_in0 = 32'd1;
	assign eq_158_in1 = state_1_last_state;
	// controller for eq_159.eq_159_in0
	// controller for eq_159.eq_159_in1
	// Insensitive connections
	assign eq_159_in0 = 32'd4;
	assign eq_159_in1 = state_1_last_state;
	// controller for eq_161.eq_161_in0
	// controller for eq_161.eq_161_in1
	// Insensitive connections
	assign eq_161_in0 = 32'd1;
	assign eq_161_in1 = state_2_last_state;
	// controller for eq_162.eq_162_in0
	// controller for eq_162.eq_162_in1
	// Insensitive connections
	assign eq_162_in0 = 32'd2;
	assign eq_162_in1 = state_2_last_state;
	// controller for eq_163.eq_163_in0
	// controller for eq_163.eq_163_in1
	// Insensitive connections
	assign eq_163_in0 = 32'd2;
	assign eq_163_in1 = state_3_last_state;
	// controller for eq_164.eq_164_in0
	// controller for eq_164.eq_164_in1
	// Insensitive connections
	assign eq_164_in0 = 32'd3;
	assign eq_164_in1 = state_3_last_state;
	// controller for eq_167.eq_167_in0
	// controller for eq_167.eq_167_in1
	// Insensitive connections
	assign eq_167_in0 = 32'd3;
	assign eq_167_in1 = state_4_last_state;
	// controller for eq_168.eq_168_in0
	// controller for eq_168.eq_168_in1
	// Insensitive connections
	assign eq_168_in0 = 32'd4;
	assign eq_168_in1 = state_4_last_state;
	// controller for eq_58.eq_58_in0
	// controller for eq_58.eq_58_in1
	// Insensitive connections
	assign eq_58_in0 = 32'd0;
	assign eq_58_in1 = state_0_entry_BB_reg;
	// controller for eq_59.eq_59_in0
	// controller for eq_59.eq_59_in1
	// Insensitive connections
	assign eq_59_in0 = 32'd0;
	assign eq_59_in1 = state_1_entry_BB_reg;
	// controller for eq_60.eq_60_in0
	// controller for eq_60.eq_60_in1
	// Insensitive connections
	assign eq_60_in0 = 32'd8;
	assign eq_60_in1 = state_1_entry_BB_reg;
	// controller for eq_62.eq_62_in0
	// controller for eq_62.eq_62_in1
	// Insensitive connections
	assign eq_62_in0 = 32'd3;
	assign eq_62_in1 = state_1_entry_BB_reg;
	// controller for eq_64.eq_64_in0
	// controller for eq_64.eq_64_in1
	// Insensitive connections
	assign eq_64_in0 = 32'd9;
	assign eq_64_in1 = state_1_entry_BB_reg;
	// controller for eq_66.eq_66_in0
	// controller for eq_66.eq_66_in1
	// Insensitive connections
	assign eq_66_in0 = 32'd10;
	assign eq_66_in1 = state_2_entry_BB_reg;
	// controller for eq_67.eq_67_in0
	// controller for eq_67.eq_67_in1
	// Insensitive connections
	assign eq_67_in0 = 32'd4;
	assign eq_67_in1 = state_3_entry_BB_reg;
	// controller for eq_69.eq_69_in0
	// controller for eq_69.eq_69_in1
	// Insensitive connections
	assign eq_69_in0 = 32'd10;
	assign eq_69_in1 = state_3_entry_BB_reg;
	// controller for eq_70.eq_70_in0
	// controller for eq_70.eq_70_in1
	// Insensitive connections
	assign eq_70_in0 = 32'd4;
	assign eq_70_in1 = state_4_entry_BB_reg;
	// controller for eq_71.eq_71_in0
	// controller for eq_71.eq_71_in1
	// Insensitive connections
	assign eq_71_in0 = 32'd6;
	assign eq_71_in1 = state_4_entry_BB_reg;
	// controller for eq_73.eq_73_in0
	// controller for eq_73.eq_73_in1
	// Insensitive connections
	assign eq_73_in0 = 32'd2;
	assign eq_73_in1 = state_4_entry_BB_reg;
	// controller for eq_75.eq_75_in0
	// controller for eq_75.eq_75_in1
	// Insensitive connections
	assign eq_75_in0 = 32'd5;
	assign eq_75_in1 = state_4_entry_BB_reg;
	// controller for eq_77.eq_77_in0
	// controller for eq_77.eq_77_in1
	// Insensitive connections
	assign eq_77_in0 = 32'd7;
	assign eq_77_in1 = state_4_entry_BB_reg;
	// controller for eq_79.eq_79_in0
	// controller for eq_79.eq_79_in1
	// Insensitive connections
	assign eq_79_in0 = 32'd1;
	assign eq_79_in1 = state_4_entry_BB_reg;
	// controller for eq_81.eq_81_in0
	// controller for eq_81.eq_81_in1
	// Insensitive connections
	assign eq_81_in0 = 32'd0;
	assign eq_81_in1 = state_0_entry_BB_reg;
	// controller for eq_82.eq_82_in0
	// controller for eq_82.eq_82_in1
	// Insensitive connections
	assign eq_82_in0 = 32'd0;
	assign eq_82_in1 = state_1_entry_BB_reg;
	// controller for eq_83.eq_83_in0
	// controller for eq_83.eq_83_in1
	// Insensitive connections
	assign eq_83_in0 = 32'd8;
	assign eq_83_in1 = state_1_entry_BB_reg;
	// controller for eq_86.eq_86_in0
	// controller for eq_86.eq_86_in1
	// Insensitive connections
	assign eq_86_in0 = 32'd3;
	assign eq_86_in1 = state_1_entry_BB_reg;
	// controller for eq_89.eq_89_in0
	// controller for eq_89.eq_89_in1
	// Insensitive connections
	assign eq_89_in0 = 32'd9;
	assign eq_89_in1 = state_1_entry_BB_reg;
	// controller for eq_92.eq_92_in0
	// controller for eq_92.eq_92_in1
	// Insensitive connections
	assign eq_92_in0 = 32'd10;
	assign eq_92_in1 = state_2_entry_BB_reg;
	// controller for eq_93.eq_93_in0
	// controller for eq_93.eq_93_in1
	// Insensitive connections
	assign eq_93_in0 = 32'd4;
	assign eq_93_in1 = state_3_entry_BB_reg;
	// controller for eq_96.eq_96_in0
	// controller for eq_96.eq_96_in1
	// Insensitive connections
	assign eq_96_in0 = 32'd10;
	assign eq_96_in1 = state_3_entry_BB_reg;
	// controller for eq_97.eq_97_in0
	// controller for eq_97.eq_97_in1
	// Insensitive connections
	assign eq_97_in0 = 32'd4;
	assign eq_97_in1 = state_4_entry_BB_reg;
	// controller for eq_98.eq_98_in0
	// controller for eq_98.eq_98_in1
	// Insensitive connections
	assign eq_98_in0 = 32'd6;
	assign eq_98_in1 = state_4_entry_BB_reg;
	// controller for icmp_icmp16.icmp_icmp16_in0
	// controller for icmp_icmp16.icmp_icmp16_in1
	// Insensitive connections
	assign icmp_icmp16_in0 = add_add15_out;
	assign icmp_icmp16_in1 = 32'd4;
	// controller for in.in_read_valid_reg
	always @(*) begin
		if (andOp_124_out) begin 
			in_read_valid_reg = -(1'd1);
		end else begin
			in_read_valid_reg = 0;
		end
	end
	// controller for notOp_102.notOp_102_in0
	// Insensitive connections
	assign notOp_102_in0 = eq_101_out;
	// controller for notOp_105.notOp_105_in0
	// Insensitive connections
	assign notOp_105_in0 = eq_104_out;
	// controller for notOp_108.notOp_108_in0
	// Insensitive connections
	assign notOp_108_in0 = eq_107_out;
	// controller for notOp_111.notOp_111_in0
	// Insensitive connections
	assign notOp_111_in0 = eq_110_out;
	// controller for notOp_140.notOp_140_in0
	// Insensitive connections
	assign notOp_140_in0 = andOp_136_out;
	// controller for notOp_142.notOp_142_in0
	// Insensitive connections
	assign notOp_142_in0 = andOp_32_out;
	// controller for notOp_144.notOp_144_in0
	// Insensitive connections
	assign notOp_144_in0 = andOp_39_out;
	// controller for notOp_146.notOp_146_in0
	// Insensitive connections
	assign notOp_146_in0 = andOp_30_out;
	// controller for notOp_148.notOp_148_in0
	// Insensitive connections
	assign notOp_148_in0 = andOp_137_out;
	// controller for notOp_150.notOp_150_in0
	// Insensitive connections
	assign notOp_150_in0 = andOp_138_out;
	// controller for notOp_152.notOp_152_in0
	// Insensitive connections
	assign notOp_152_in0 = andOp_139_out;
	// controller for notOp_154.notOp_154_in0
	// Insensitive connections
	assign notOp_154_in0 = andOp_51_out;
	// controller for notOp_21.notOp_21_in0
	// Insensitive connections
	assign notOp_21_in0 = andOp_20_out;
	// controller for notOp_23.notOp_23_in0
	// Insensitive connections
	assign notOp_23_in0 = andOp_22_out;
	// controller for notOp_25.notOp_25_in0
	// Insensitive connections
	assign notOp_25_in0 = andOp_24_out;
	// controller for notOp_27.notOp_27_in0
	// Insensitive connections
	assign notOp_27_in0 = andOp_26_out;
	// controller for notOp_29.notOp_29_in0
	// Insensitive connections
	assign notOp_29_in0 = andOp_28_out;
	// controller for notOp_31.notOp_31_in0
	// Insensitive connections
	assign notOp_31_in0 = in_read_ready;
	// controller for notOp_34.notOp_34_in0
	// Insensitive connections
	assign notOp_34_in0 = andOp_33_out;
	// controller for notOp_36.notOp_36_in0
	// Insensitive connections
	assign notOp_36_in0 = andOp_35_out;
	// controller for notOp_38.notOp_38_in0
	// Insensitive connections
	assign notOp_38_in0 = data_in_4_17_out_data;
	// controller for notOp_41.notOp_41_in0
	// Insensitive connections
	assign notOp_41_in0 = andOp_40_out;
	// controller for notOp_43.notOp_43_in0
	// Insensitive connections
	assign notOp_43_in0 = andOp_42_out;
	// controller for notOp_45.notOp_45_in0
	// Insensitive connections
	assign notOp_45_in0 = data_in_4_17_out_data;
	// controller for notOp_48.notOp_48_in0
	// Insensitive connections
	assign notOp_48_in0 = andOp_47_out;
	// controller for notOp_50.notOp_50_in0
	// Insensitive connections
	assign notOp_50_in0 = out_write_ready;
	// controller for notOp_53.notOp_53_in0
	// Insensitive connections
	assign notOp_53_in0 = andOp_52_out;
	// controller for notOp_55.notOp_55_in0
	// Insensitive connections
	assign notOp_55_in0 = andOp_54_out;
	// controller for notOp_57.notOp_57_in0
	// Insensitive connections
	assign notOp_57_in0 = andOp_56_out;
	// controller for notOp_84.notOp_84_in0
	// Insensitive connections
	assign notOp_84_in0 = eq_83_out;
	// controller for notOp_87.notOp_87_in0
	// Insensitive connections
	assign notOp_87_in0 = eq_86_out;
	// controller for notOp_90.notOp_90_in0
	// Insensitive connections
	assign notOp_90_in0 = eq_89_out;
	// controller for notOp_94.notOp_94_in0
	// Insensitive connections
	assign notOp_94_in0 = eq_93_out;
	// controller for notOp_99.notOp_99_in0
	// Insensitive connections
	assign notOp_99_in0 = eq_98_out;
	// controller for orOp_61.orOp_61_in0
	// controller for orOp_61.orOp_61_in1
	// Insensitive connections
	assign orOp_61_in0 = eq_60_out;
	assign orOp_61_in1 = andOp_26_out;
	// controller for orOp_63.orOp_63_in0
	// controller for orOp_63.orOp_63_in1
	// Insensitive connections
	assign orOp_63_in0 = eq_62_out;
	assign orOp_63_in1 = andOp_20_out;
	// controller for orOp_65.orOp_65_in0
	// controller for orOp_65.orOp_65_in1
	// Insensitive connections
	assign orOp_65_in0 = eq_64_out;
	assign orOp_65_in1 = andOp_24_out;
	// controller for orOp_68.orOp_68_in0
	// controller for orOp_68.orOp_68_in1
	// Insensitive connections
	assign orOp_68_in0 = eq_67_out;
	assign orOp_68_in1 = andOp_33_out;
	// controller for orOp_72.orOp_72_in0
	// controller for orOp_72.orOp_72_in1
	// Insensitive connections
	assign orOp_72_in0 = eq_71_out;
	assign orOp_72_in1 = andOp_52_out;
	// controller for orOp_74.orOp_74_in0
	// controller for orOp_74.orOp_74_in1
	// Insensitive connections
	assign orOp_74_in0 = eq_73_out;
	assign orOp_74_in1 = andOp_54_out;
	// controller for orOp_76.orOp_76_in0
	// controller for orOp_76.orOp_76_in1
	// Insensitive connections
	assign orOp_76_in0 = eq_75_out;
	assign orOp_76_in1 = andOp_56_out;
	// controller for orOp_78.orOp_78_in0
	// controller for orOp_78.orOp_78_in1
	// Insensitive connections
	assign orOp_78_in0 = eq_77_out;
	assign orOp_78_in1 = andOp_49_out;
	// controller for orOp_80.orOp_80_in0
	// controller for orOp_80.orOp_80_in1
	// Insensitive connections
	assign orOp_80_in0 = eq_79_out;
	assign orOp_80_in1 = andOp_37_out;
	// controller for out.out_in_data_reg
	always @(*) begin
		if (andOp_132_out) begin 
			out_in_data_reg = rdata_ram_0;
		end else begin
			out_in_data_reg = 0;
		end
	end
	// controller for out.out_write_valid_reg
	always @(*) begin
		if (andOp_133_out) begin 
			out_write_valid_reg = -(1'd1);
		end else begin
			out_write_valid_reg = 0;
		end
	end
	// controller for phi_phi6.phi_phi6_in
	// controller for phi_phi6.phi_phi6_last_block
	// controller for phi_phi6.phi_phi6_s
	// Insensitive connections
	assign phi_phi6_in = concat_121_out;
	assign phi_phi6_last_block = bb_3_predecessor_in_state_1_out_data;
	assign phi_phi6_s = concat_122_out;
	// controller for ram_0.raddr_ram_0_reg
	always @(*) begin
		if (andOp_117_out) begin 
			raddr_ram_0_reg = 32'd0;
		end else if (andOp_119_out) begin 
			raddr_ram_0_reg = 32'd0;
		end else begin
			raddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.waddr_ram_0_reg
	always @(*) begin
		if (andOp_116_out) begin 
			waddr_ram_0_reg = 32'd0;
		end else if (andOp_118_out) begin 
			waddr_ram_0_reg = 32'd0;
		end else begin
			waddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wdata_ram_0_reg
	always @(*) begin
		if (andOp_116_out) begin 
			wdata_ram_0_reg = 32'd0;
		end else if (andOp_118_out) begin 
			wdata_ram_0_reg = add_add13_out;
		end else begin
			wdata_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wen_ram_0_reg
	always @(*) begin
		if (andOp_116_out) begin 
			wen_ram_0_reg = 1'd1;
		end else if (andOp_118_out) begin 
			wen_ram_0_reg = 1'd1;
		end else begin
			wen_ram_0_reg = 0;
		end
	end
	// controller for ret26.valid_reg
	always @(*) begin
		if (andOp_135_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// controller for tmp_output_127.tmp_output_127_in_data
	always @(*) begin
		if (eq_128_out) begin 
			tmp_output_127_in_data = in_out_data;
		end else begin
			tmp_output_127_in_data = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			data_store_0_0 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_0 <= data_in_0_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_2 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_2 <= data_in_0_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_4 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_4 <= data_in_1_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_6 <= 0;
		end else begin
			if (andOp_160_out) begin
				data_store_1_6 <= phi_phi6_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_8 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_8 <= data_in_2_9_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_10 <= 0;
		end else begin
			if (andOp_165_out) begin
				data_store_3_10 <= add_add15_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_11 <= 0;
		end else begin
			if (andOp_166_out) begin
				data_store_3_11 <= icmp_icmp16_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_12 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_12 <= data_in_3_13_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_14 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_14 <= data_in_4_15_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_16 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_16 <= data_in_4_17_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_18 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_18 <= data_in_4_19_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_136_out) begin
				global_state <= 32'd1;
			end
			if (andOp_137_out) begin
				global_state <= 32'd3;
			end
			if (andOp_138_out) begin
				global_state <= 32'd4;
			end
			if (andOp_139_out) begin
				global_state <= 32'd4;
			end
			if (andOp_30_out) begin
				global_state <= 32'd2;
			end
			if (andOp_32_out) begin
				global_state <= 32'd1;
			end
			if (andOp_39_out) begin
				global_state <= 32'd1;
			end
			if (andOp_51_out) begin
				global_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (1'd1) begin
				state_0_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_136_out) begin
				state_1_entry_BB_reg <= 32'd0;
			end
			if (andOp_32_out) begin
				state_1_entry_BB_reg <= 32'd9;
			end
			if (andOp_39_out) begin
				state_1_entry_BB_reg <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_136_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_145_out) begin
				state_1_is_active <= 1'd0;
			end
			if (andOp_32_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_39_out) begin
				state_1_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_136_out) begin
				state_1_last_BB_reg <= bb_0_predecessor_in_state_0_out_data;
			end
			if (andOp_32_out) begin
				state_1_last_BB_reg <= 32'd9;
			end
			if (andOp_39_out) begin
				state_1_last_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_136_out) begin
				state_1_last_state <= 32'd0;
			end
			if (andOp_32_out) begin
				state_1_last_state <= 32'd1;
			end
			if (andOp_39_out) begin
				state_1_last_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_30_out) begin
				state_2_entry_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_147_out) begin
				state_2_is_active <= 1'd0;
			end
			if (andOp_30_out) begin
				state_2_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_30_out) begin
				state_2_last_BB_reg <= 32'd9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_30_out) begin
				state_2_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_137_out) begin
				state_3_entry_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_137_out) begin
				state_3_is_active <= 1'd1;
			end
			if (andOp_149_out) begin
				state_3_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_137_out) begin
				state_3_last_BB_reg <= bb_10_predecessor_in_state_2_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_state <= 0;
		end else begin
			if (andOp_137_out) begin
				state_3_last_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_138_out) begin
				state_4_entry_BB_reg <= 32'd4;
			end
			if (andOp_139_out) begin
				state_4_entry_BB_reg <= 32'd2;
			end
			if (andOp_51_out) begin
				state_4_entry_BB_reg <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_138_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_139_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_155_out) begin
				state_4_is_active <= 1'd0;
			end
			if (andOp_51_out) begin
				state_4_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_138_out) begin
				state_4_last_BB_reg <= bb_4_predecessor_in_state_3_out_data;
			end
			if (andOp_139_out) begin
				state_4_last_BB_reg <= bb_2_predecessor_in_state_4_out_data;
			end
			if (andOp_51_out) begin
				state_4_last_BB_reg <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_state <= 0;
		end else begin
			if (andOp_138_out) begin
				state_4_last_state <= 32'd3;
			end
			if (andOp_139_out) begin
				state_4_last_state <= 32'd4;
			end
			if (andOp_51_out) begin
				state_4_last_state <= 32'd4;
			end
		end
	end

endmodule

