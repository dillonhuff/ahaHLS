
//------> /hd/cad/mentor/2016.9/Mgc_home/pkgs/siflibs/mgc_in_wire_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_in_wire_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  output [width-1:0] d;
  output             lz;
  input              vz;
  input  [width-1:0] z;

  wire               vd;
  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;
  assign vd = vz;

endmodule


//------> /hd/cad/mentor/2016.9/Mgc_home/pkgs/siflibs/mgc_out_stdreg_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_stdreg_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  input  [width-1:0] d;
  output             lz;
  input              vz;
  output [width-1:0] z;

  wire               vd;
  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;
  assign vd = vz;

endmodule



//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0/263344 Production Release
//  HLS Date:       Sun Jul  3 19:13:39 PDT 2016
// 
//  Generated by:   dhuff@kiwi
//  Generated date: Mon Feb 18 17:38:21 2019
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    dct_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module dct_core_core_fsm (
  dillons_clk, rst, core_wen, fsm_output, for_C_0_tr0
);
  input dillons_clk;
  input rst;
  input core_wen;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;
  input for_C_0_tr0;


  // FSM State Type Declaration for dct_core_core_fsm_1
  parameter
    main_C_0 = 2'd0,
    for_C_0 = 2'd1,
    main_C_1 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : dct_core_core_fsm_1
    case (state_var)
      for_C_0 : begin
        fsm_output = 3'b10;
        if ( for_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 3'b100;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 3'b1;
        state_var_NS = for_C_0;
      end
    endcase
  end

  always @(posedge dillons_clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    dct_core_staller
// ------------------------------------------------------------------


module dct_core_staller (
  dillons_clk, rst, core_wen, in_rsci_wen_comp, core_wten, out_rsci_wen_comp
);
  input dillons_clk;
  input rst;
  output core_wen;
  input in_rsci_wen_comp;
  output core_wten;
  reg core_wten;
  input out_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = in_rsci_wen_comp & out_rsci_wen_comp;
  always @(posedge dillons_clk) begin
    if ( rst ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    dct_core_out_rsci_out_wait_dp
// ------------------------------------------------------------------


module dct_core_out_rsci_out_wait_dp (
  dillons_clk, rst, out_rsci_oswt, out_rsci_wen_comp, out_rsci_biwt, out_rsci_bdwt
);
  input dillons_clk;
  input rst;
  input out_rsci_oswt;
  output out_rsci_wen_comp;
  input out_rsci_biwt;
  input out_rsci_bdwt;


  // Interconnect Declarations
  reg out_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign out_rsci_wen_comp = (~ out_rsci_oswt) | out_rsci_biwt | out_rsci_bcwt;
  always @(posedge dillons_clk) begin
    if ( rst ) begin
      out_rsci_bcwt <= 1'b0;
    end
    else begin
      out_rsci_bcwt <= ~((~(out_rsci_bcwt | out_rsci_biwt)) | out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    dct_core_out_rsci_out_wait_ctrl
// ------------------------------------------------------------------


module dct_core_out_rsci_out_wait_ctrl (
  dillons_clk, rst, core_wen, core_wten, out_rsci_oswt, out_rsci_biwt, out_rsci_bdwt,
      out_rsci_ld_core_sct, out_rsci_vd
);
  input dillons_clk;
  input rst;
  input core_wen;
  input core_wten;
  input out_rsci_oswt;
  output out_rsci_biwt;
  output out_rsci_bdwt;
  output out_rsci_ld_core_sct;
  input out_rsci_vd;


  // Interconnect Declarations
  wire out_rsci_ogwt;
  wire out_rsci_pdswt0;
  reg out_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign out_rsci_pdswt0 = (~ core_wten) & out_rsci_oswt;
  assign out_rsci_biwt = out_rsci_ogwt & out_rsci_vd;
  assign out_rsci_ogwt = out_rsci_pdswt0 | out_rsci_icwt;
  assign out_rsci_bdwt = out_rsci_oswt & core_wen;
  assign out_rsci_ld_core_sct = out_rsci_oswt & out_rsci_ogwt;
  always @(posedge dillons_clk) begin
    if ( rst ) begin
      out_rsci_icwt <= 1'b0;
    end
    else begin
      out_rsci_icwt <= ~((~(out_rsci_icwt | out_rsci_pdswt0)) | out_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    dct_core_in_rsci_in_wait_dp
// ------------------------------------------------------------------


module dct_core_in_rsci_in_wait_dp (
  dillons_clk, rst, in_rsci_oswt, in_rsci_wen_comp, in_rsci_d_mxwt, in_rsci_biwt,
      in_rsci_bdwt, in_rsci_d
);
  input dillons_clk;
  input rst;
  input in_rsci_oswt;
  output in_rsci_wen_comp;
  output [31:0] in_rsci_d_mxwt;
  input in_rsci_biwt;
  input in_rsci_bdwt;
  input [31:0] in_rsci_d;


  // Interconnect Declarations
  reg in_rsci_bcwt;
  reg [31:0] in_rsci_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign in_rsci_wen_comp = (~ in_rsci_oswt) | in_rsci_biwt | in_rsci_bcwt;
  assign in_rsci_d_mxwt = MUX_v_32_2_2(in_rsci_d, in_rsci_d_bfwt, in_rsci_bcwt);
  always @(posedge dillons_clk) begin
    if ( rst ) begin
      in_rsci_bcwt <= 1'b0;
      in_rsci_d_bfwt <= 32'b0;
    end
    else begin
      in_rsci_bcwt <= ~((~(in_rsci_bcwt | in_rsci_biwt)) | in_rsci_bdwt);
      in_rsci_d_bfwt <= in_rsci_d_mxwt;
    end
  end

  function [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    dct_core_in_rsci_in_wait_ctrl
// ------------------------------------------------------------------


module dct_core_in_rsci_in_wait_ctrl (
  dillons_clk, rst, core_wen, in_rsci_oswt, core_wten, in_rsci_biwt, in_rsci_bdwt,
      in_rsci_ld_core_sct, in_rsci_vd
);
  input dillons_clk;
  input rst;
  input core_wen;
  input in_rsci_oswt;
  input core_wten;
  output in_rsci_biwt;
  output in_rsci_bdwt;
  output in_rsci_ld_core_sct;
  input in_rsci_vd;


  // Interconnect Declarations
  wire in_rsci_ogwt;
  wire in_rsci_pdswt0;
  reg in_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign in_rsci_pdswt0 = (~ core_wten) & in_rsci_oswt;
  assign in_rsci_biwt = in_rsci_ogwt & in_rsci_vd;
  assign in_rsci_ogwt = in_rsci_pdswt0 | in_rsci_icwt;
  assign in_rsci_bdwt = in_rsci_oswt & core_wen;
  assign in_rsci_ld_core_sct = in_rsci_oswt & in_rsci_ogwt;
  always @(posedge dillons_clk) begin
    if ( rst ) begin
      in_rsci_icwt <= 1'b0;
    end
    else begin
      in_rsci_icwt <= ~((~(in_rsci_icwt | in_rsci_pdswt0)) | in_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    dct_core_out_rsci
// ------------------------------------------------------------------


module dct_core_out_rsci (
  dillons_clk, rst, out_rsc_z, out_rsc_vz, out_rsc_lz, core_wen, core_wten, out_rsci_oswt,
      out_rsci_wen_comp, out_rsci_d
);
  input dillons_clk;
  input rst;
  output [31:0] out_rsc_z;
  input out_rsc_vz;
  output out_rsc_lz;
  input core_wen;
  input core_wten;
  input out_rsci_oswt;
  output out_rsci_wen_comp;
  input [31:0] out_rsci_d;


  // Interconnect Declarations
  wire out_rsci_biwt;
  wire out_rsci_bdwt;
  wire out_rsci_ld_core_sct;
  wire out_rsci_vd;


  // Interconnect Declarations for Component Instantiations 
  mgc_out_stdreg_wait_v1 #(.rscid(32'sd2),
  .width(32'sd32)) out_rsci (
      .ld(out_rsci_ld_core_sct),
      .vd(out_rsci_vd),
      .d(out_rsci_d),
      .lz(out_rsc_lz),
      .vz(out_rsc_vz),
      .z(out_rsc_z)
    );
  dct_core_out_rsci_out_wait_ctrl dct_core_out_rsci_out_wait_ctrl_inst (
      .dillons_clk(dillons_clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .out_rsci_oswt(out_rsci_oswt),
      .out_rsci_biwt(out_rsci_biwt),
      .out_rsci_bdwt(out_rsci_bdwt),
      .out_rsci_ld_core_sct(out_rsci_ld_core_sct),
      .out_rsci_vd(out_rsci_vd)
    );
  dct_core_out_rsci_out_wait_dp dct_core_out_rsci_out_wait_dp_inst (
      .dillons_clk(dillons_clk),
      .rst(rst),
      .out_rsci_oswt(out_rsci_oswt),
      .out_rsci_wen_comp(out_rsci_wen_comp),
      .out_rsci_biwt(out_rsci_biwt),
      .out_rsci_bdwt(out_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    dct_core_in_rsci
// ------------------------------------------------------------------


module dct_core_in_rsci (
  dillons_clk, rst, in_rsc_z, in_rsc_vz, in_rsc_lz, core_wen, in_rsci_oswt, in_rsci_wen_comp,
      in_rsci_d_mxwt, core_wten
);
  input dillons_clk;
  input rst;
  input [31:0] in_rsc_z;
  input in_rsc_vz;
  output in_rsc_lz;
  input core_wen;
  input in_rsci_oswt;
  output in_rsci_wen_comp;
  output [31:0] in_rsci_d_mxwt;
  input core_wten;


  // Interconnect Declarations
  wire in_rsci_biwt;
  wire in_rsci_bdwt;
  wire in_rsci_ld_core_sct;
  wire in_rsci_vd;
  wire [31:0] in_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_wire_wait_v1 #(.rscid(32'sd1),
  .width(32'sd32)) in_rsci (
      .ld(in_rsci_ld_core_sct),
      .vd(in_rsci_vd),
      .d(in_rsci_d),
      .lz(in_rsc_lz),
      .vz(in_rsc_vz),
      .z(in_rsc_z)
    );
  dct_core_in_rsci_in_wait_ctrl dct_core_in_rsci_in_wait_ctrl_inst (
      .dillons_clk(dillons_clk),
      .rst(rst),
      .core_wen(core_wen),
      .in_rsci_oswt(in_rsci_oswt),
      .core_wten(core_wten),
      .in_rsci_biwt(in_rsci_biwt),
      .in_rsci_bdwt(in_rsci_bdwt),
      .in_rsci_ld_core_sct(in_rsci_ld_core_sct),
      .in_rsci_vd(in_rsci_vd)
    );
  dct_core_in_rsci_in_wait_dp dct_core_in_rsci_in_wait_dp_inst (
      .dillons_clk(dillons_clk),
      .rst(rst),
      .in_rsci_oswt(in_rsci_oswt),
      .in_rsci_wen_comp(in_rsci_wen_comp),
      .in_rsci_d_mxwt(in_rsci_d_mxwt),
      .in_rsci_biwt(in_rsci_biwt),
      .in_rsci_bdwt(in_rsci_bdwt),
      .in_rsci_d(in_rsci_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    dct_core
// ------------------------------------------------------------------


module dct_core (
  dillons_clk, rst, in_rsc_z, in_rsc_vz, in_rsc_lz, out_rsc_z, out_rsc_vz, out_rsc_lz
);
  input dillons_clk;
  input rst;
  input [31:0] in_rsc_z;
  input in_rsc_vz;
  output in_rsc_lz;
  output [31:0] out_rsc_z;
  input out_rsc_vz;
  output out_rsc_lz;


  // Interconnect Declarations
  wire core_wen;
  wire in_rsci_wen_comp;
  wire [31:0] in_rsci_d_mxwt;
  wire core_wten;
  wire out_rsci_wen_comp;
  reg [31:0] out_rsci_d;
  wire [2:0] fsm_output;
  reg [31:0] sum_sva;
  reg [1:0] for_i_2_0_sva_1_0_1;
  wire and_6_cse;
  wire [2:0] for_i_2_0_sva_1;
  wire [3:0] nl_for_i_2_0_sva_1;
  reg reg_out_rsci_ld_core_psct_cse;
  reg reg_in_rsci_ld_core_psct_cse;
  wire [31:0] sum_sva_1;
  wire [32:0] nl_sum_sva_1;


  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_dct_core_core_fsm_inst_for_C_0_tr0;
  assign nl_dct_core_core_fsm_inst_for_C_0_tr0 = for_i_2_0_sva_1[2];
  dct_core_in_rsci dct_core_in_rsci_inst (
      .dillons_clk(dillons_clk),
      .rst(rst),
      .in_rsc_z(in_rsc_z),
      .in_rsc_vz(in_rsc_vz),
      .in_rsc_lz(in_rsc_lz),
      .core_wen(core_wen),
      .in_rsci_oswt(reg_in_rsci_ld_core_psct_cse),
      .in_rsci_wen_comp(in_rsci_wen_comp),
      .in_rsci_d_mxwt(in_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  dct_core_out_rsci dct_core_out_rsci_inst (
      .dillons_clk(dillons_clk),
      .rst(rst),
      .out_rsc_z(out_rsc_z),
      .out_rsc_vz(out_rsc_vz),
      .out_rsc_lz(out_rsc_lz),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .out_rsci_oswt(reg_out_rsci_ld_core_psct_cse),
      .out_rsci_wen_comp(out_rsci_wen_comp),
      .out_rsci_d(out_rsci_d)
    );
  dct_core_staller dct_core_staller_inst (
      .dillons_clk(dillons_clk),
      .rst(rst),
      .core_wen(core_wen),
      .in_rsci_wen_comp(in_rsci_wen_comp),
      .core_wten(core_wten),
      .out_rsci_wen_comp(out_rsci_wen_comp)
    );
  dct_core_core_fsm dct_core_core_fsm_inst (
      .dillons_clk(dillons_clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output),
      .for_C_0_tr0(nl_dct_core_core_fsm_inst_for_C_0_tr0[0:0])
    );
  assign nl_sum_sva_1 = sum_sva + in_rsci_d_mxwt;
  assign sum_sva_1 = nl_sum_sva_1[31:0];
  assign nl_for_i_2_0_sva_1 = conv_u2u_2_3(for_i_2_0_sva_1_0_1) + 3'b1;
  assign for_i_2_0_sva_1 = nl_for_i_2_0_sva_1[2:0];
  assign and_6_cse = (for_i_2_0_sva_1[2]) & (fsm_output[1]);
  always @(posedge dillons_clk) begin
    if ( rst ) begin
      for_i_2_0_sva_1_0_1 <= 2'b0;
      sum_sva <= 32'b0;
      reg_out_rsci_ld_core_psct_cse <= 1'b0;
      reg_in_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen ) begin
      for_i_2_0_sva_1_0_1 <= MUX_v_2_2_2(2'b00, (for_i_2_0_sva_1[1:0]), (fsm_output[1]));
      sum_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000, sum_sva_1, (fsm_output[1]));
      reg_out_rsci_ld_core_psct_cse <= and_6_cse;
      reg_in_rsci_ld_core_psct_cse <= ~(and_6_cse | (fsm_output[2]));
    end
  end
  always @(posedge dillons_clk) begin
    if ( rst ) begin
      out_rsci_d <= 32'b0;
    end
    else if ( core_wen & (for_i_2_0_sva_1[2]) & (fsm_output[1]) ) begin
      out_rsci_d <= sum_sva_1;
    end
  end

  function [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function  [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    dct
// ------------------------------------------------------------------


module dct (
  dillons_clk, rst, in_rsc_z, in_rsc_vz, in_rsc_lz, out_rsc_z, out_rsc_vz, out_rsc_lz
);
  input dillons_clk;
  input rst;
  input [31:0] in_rsc_z;
  input in_rsc_vz;
  output in_rsc_lz;
  output [31:0] out_rsc_z;
  input out_rsc_vz;
  output out_rsc_lz;



  // Interconnect Declarations for Component Instantiations 
  dct_core dct_core_inst (
      .dillons_clk(dillons_clk),
      .rst(rst),
      .in_rsc_z(in_rsc_z),
      .in_rsc_vz(in_rsc_vz),
      .in_rsc_lz(in_rsc_lz),
      .out_rsc_z(out_rsc_z),
      .out_rsc_vz(out_rsc_vz),
      .out_rsc_lz(out_rsc_lz)
    );
endmodule



