module axi_wb(input [0:0] clk, input [0:0] rst, output [7:0] arg_1_raddr, output [7:0] arg_1_waddr, output [7:0] arg_1_wdata, output [0:0] arg_1_wen, input [7:0] arg_1_rdata, output [15:0] arg_2_raddr, output [15:0] arg_2_waddr, output [15:0] arg_2_wdata, output [0:0] arg_2_wen, input [15:0] arg_2_rdata, output [0:0] valid, output [15:0] arg_3_s_axi_araddr, output [1:0] arg_3_s_axi_arburst, output [7:0] arg_3_s_axi_arlen, output [2:0] arg_3_s_axi_arsize, output [0:0] arg_3_s_axi_arvalid, output [15:0] arg_3_s_axi_awaddr, output [1:0] arg_3_s_axi_awburst, output [7:0] arg_3_s_axi_awlen, output [2:0] arg_3_s_axi_awsize, output [0:0] arg_3_s_axi_awvalid, output [0:0] arg_3_s_axi_bready, output [0:0] arg_3_s_axi_rready, output [31:0] arg_3_s_axi_wdata, output [3:0] arg_3_s_axi_wstrb, output [0:0] arg_3_s_axi_wvalid, input [0:0] arg_3_s_axi_arready, input [0:0] arg_3_s_axi_awready, input [0:0] arg_3_s_axi_bvalid, input [31:0] arg_3_s_axi_rdata, input [0:0] arg_3_s_axi_rvalid, input [0:0] arg_3_s_axi_wready, output [31:0] arg_0_in_data, output [0:0] arg_0_read_valid, output [0:0] arg_0_write_valid, input [31:0] arg_0_out_data, input [0:0] arg_0_read_ready, input [0:0] arg_0_write_ready);

	reg [7:0] arg_1_raddr_reg;
	reg [7:0] arg_1_waddr_reg;
	reg [7:0] arg_1_wdata_reg;
	reg [0:0] arg_1_wen_reg;
	reg [15:0] arg_2_raddr_reg;
	reg [15:0] arg_2_waddr_reg;
	reg [15:0] arg_2_wdata_reg;
	reg [0:0] arg_2_wen_reg;
	reg [0:0] valid_reg;
	reg [15:0] arg_3_s_axi_araddr_reg;
	reg [1:0] arg_3_s_axi_arburst_reg;
	reg [7:0] arg_3_s_axi_arlen_reg;
	reg [2:0] arg_3_s_axi_arsize_reg;
	reg [0:0] arg_3_s_axi_arvalid_reg;
	reg [15:0] arg_3_s_axi_awaddr_reg;
	reg [1:0] arg_3_s_axi_awburst_reg;
	reg [7:0] arg_3_s_axi_awlen_reg;
	reg [2:0] arg_3_s_axi_awsize_reg;
	reg [0:0] arg_3_s_axi_awvalid_reg;
	reg [0:0] arg_3_s_axi_bready_reg;
	reg [0:0] arg_3_s_axi_rready_reg;
	reg [31:0] arg_3_s_axi_wdata_reg;
	reg [3:0] arg_3_s_axi_wstrb_reg;
	reg [0:0] arg_3_s_axi_wvalid_reg;
	reg [31:0] arg_0_in_data_reg;
	reg [0:0] arg_0_read_valid_reg;
	reg [0:0] arg_0_write_valid_reg;

	assign arg_1_raddr = arg_1_raddr_reg;
	assign arg_1_waddr = arg_1_waddr_reg;
	assign arg_1_wdata = arg_1_wdata_reg;
	assign arg_1_wen = arg_1_wen_reg;
	assign arg_2_raddr = arg_2_raddr_reg;
	assign arg_2_waddr = arg_2_waddr_reg;
	assign arg_2_wdata = arg_2_wdata_reg;
	assign arg_2_wen = arg_2_wen_reg;
	assign valid = valid_reg;
	assign arg_3_s_axi_araddr = arg_3_s_axi_araddr_reg;
	assign arg_3_s_axi_arburst = arg_3_s_axi_arburst_reg;
	assign arg_3_s_axi_arlen = arg_3_s_axi_arlen_reg;
	assign arg_3_s_axi_arsize = arg_3_s_axi_arsize_reg;
	assign arg_3_s_axi_arvalid = arg_3_s_axi_arvalid_reg;
	assign arg_3_s_axi_awaddr = arg_3_s_axi_awaddr_reg;
	assign arg_3_s_axi_awburst = arg_3_s_axi_awburst_reg;
	assign arg_3_s_axi_awlen = arg_3_s_axi_awlen_reg;
	assign arg_3_s_axi_awsize = arg_3_s_axi_awsize_reg;
	assign arg_3_s_axi_awvalid = arg_3_s_axi_awvalid_reg;
	assign arg_3_s_axi_bready = arg_3_s_axi_bready_reg;
	assign arg_3_s_axi_rready = arg_3_s_axi_rready_reg;
	assign arg_3_s_axi_wdata = arg_3_s_axi_wdata_reg;
	assign arg_3_s_axi_wstrb = arg_3_s_axi_wstrb_reg;
	assign arg_3_s_axi_wvalid = arg_3_s_axi_wvalid_reg;
	assign arg_0_in_data = arg_0_in_data_reg;
	assign arg_0_read_valid = arg_0_read_valid_reg;
	assign arg_0_write_valid = arg_0_write_valid_reg;

	// Start debug wires and ports

	initial begin
	end





	// End debug wires and ports

	// Start Functional Units
	br_dummy br_unit();

	wire [31:0] sgt_in0_sext_21;
	wire [63:0] sgt_out_sext_21;
	sext sext_21(.in(sgt_in0_sext_21), .out(sgt_out_sext_21));

	wire [31:0] add_in0_add_22;
	wire [31:0] add_in1_add_22;
	wire [31:0] add_out_add_22;
	add #(.WIDTH(32)) add_add_22(.in0(add_in0_add_22), .in1(add_in1_add_22), .out(add_out_add_22));

	wire [7:0] cmp_in0_icmp_33;
	wire [7:0] cmp_in1_icmp_33;
	wire [0:0] cmp_out_icmp_33;
	slt #(.WIDTH(8)) icmp_33(.in0(cmp_in0_icmp_33), .in1(cmp_in1_icmp_33), .out(cmp_out_icmp_33));

	wire [31:0] trunc_in_trunc_23;
	wire [7:0] trunc_out_trunc_23;
	trunc #(.IN_WIDTH(32), .OUT_WIDTH(8)) trunc_23(.in(trunc_in_trunc_23), .out(trunc_out_trunc_23));

	wire [15:0] phi_in_phi_5;
	wire [31:0] phi_last_block_phi_5;
	wire [63:0] phi_s_phi_5;
	wire [31:0] phi_out_phi_5;
	phi #(.NB_PAIR(2), .WIDTH(8)) phi_5(.in(phi_in_phi_5), .last_block(phi_last_block_phi_5), .out(phi_out_phi_5), .s(phi_s_phi_5));

	wire [31:0] sgt_in0_sext_8;
	wire [63:0] sgt_out_sext_8;
	sext sext_8(.in(sgt_in0_sext_8), .out(sgt_out_sext_8));

	wire [31:0] sgt_in0_sext_12;
	wire [63:0] sgt_out_sext_12;
	sext sext_12(.in(sgt_in0_sext_12), .out(sgt_out_sext_12));

	wire [31:0] cmp_in0_icmp_13;
	wire [31:0] cmp_in1_icmp_13;
	wire [0:0] cmp_out_icmp_13;
	eq #(.WIDTH(32)) icmp_13(.in0(cmp_in0_icmp_13), .in1(cmp_in1_icmp_13), .out(cmp_out_icmp_13));

	wire [31:0] cmp_in0_icmp_15;
	wire [31:0] cmp_in1_icmp_15;
	wire [0:0] cmp_out_icmp_15;
	eq #(.WIDTH(32)) icmp_15(.in0(cmp_in0_icmp_15), .in1(cmp_in1_icmp_15), .out(cmp_out_icmp_15));

	add call_35();

	wire [31:0] sgt_in0_sext_30;
	wire [63:0] sgt_out_sext_30;
	sext sext_30(.in(sgt_in0_sext_30), .out(sgt_out_sext_30));

	wire [31:0] cmp_in0_icmp_31;
	wire [31:0] cmp_in1_icmp_31;
	wire [0:0] cmp_out_icmp_31;
	eq #(.WIDTH(32)) icmp_31(.in0(cmp_in0_icmp_31), .in1(cmp_in1_icmp_31), .out(cmp_out_icmp_31));

	reg [7:0] data_in_0_1_in_data;
	wire [7:0] data_in_0_1_out_data;
	hls_wire #(.WIDTH(8)) data_in_0_1(.in_data(data_in_0_1_in_data), .out_data(data_in_0_1_out_data));

	reg [15:0] data_in_0_3_in_data;
	wire [15:0] data_in_0_3_out_data;
	hls_wire #(.WIDTH(16)) data_in_0_3(.in_data(data_in_0_3_in_data), .out_data(data_in_0_3_out_data));

	reg [7:0] data_in_0_5_in_data;
	wire [7:0] data_in_0_5_out_data;
	hls_wire #(.WIDTH(8)) data_in_0_5(.in_data(data_in_0_5_in_data), .out_data(data_in_0_5_out_data));

	reg [7:0] data_in_0_7_in_data;
	wire [7:0] data_in_0_7_out_data;
	hls_wire #(.WIDTH(8)) data_in_0_7(.in_data(data_in_0_7_in_data), .out_data(data_in_0_7_out_data));

	reg [31:0] data_in_0_9_in_data;
	wire [31:0] data_in_0_9_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_9(.in_data(data_in_0_9_in_data), .out_data(data_in_0_9_out_data));

	reg [7:0] data_in_1_11_in_data;
	wire [7:0] data_in_1_11_out_data;
	hls_wire #(.WIDTH(8)) data_in_1_11(.in_data(data_in_1_11_in_data), .out_data(data_in_1_11_out_data));

	reg [15:0] data_in_1_13_in_data;
	wire [15:0] data_in_1_13_out_data;
	hls_wire #(.WIDTH(16)) data_in_1_13(.in_data(data_in_1_13_in_data), .out_data(data_in_1_13_out_data));

	reg [7:0] data_in_1_15_in_data;
	wire [7:0] data_in_1_15_out_data;
	hls_wire #(.WIDTH(8)) data_in_1_15(.in_data(data_in_1_15_in_data), .out_data(data_in_1_15_out_data));

	reg [7:0] data_in_1_17_in_data;
	wire [7:0] data_in_1_17_out_data;
	hls_wire #(.WIDTH(8)) data_in_1_17(.in_data(data_in_1_17_in_data), .out_data(data_in_1_17_out_data));

	reg [31:0] data_in_1_19_in_data;
	wire [31:0] data_in_1_19_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_19(.in_data(data_in_1_19_in_data), .out_data(data_in_1_19_out_data));

	reg [7:0] data_in_2_21_in_data;
	wire [7:0] data_in_2_21_out_data;
	hls_wire #(.WIDTH(8)) data_in_2_21(.in_data(data_in_2_21_in_data), .out_data(data_in_2_21_out_data));

	reg [15:0] data_in_2_23_in_data;
	wire [15:0] data_in_2_23_out_data;
	hls_wire #(.WIDTH(16)) data_in_2_23(.in_data(data_in_2_23_in_data), .out_data(data_in_2_23_out_data));

	reg [7:0] data_in_2_25_in_data;
	wire [7:0] data_in_2_25_out_data;
	hls_wire #(.WIDTH(8)) data_in_2_25(.in_data(data_in_2_25_in_data), .out_data(data_in_2_25_out_data));

	reg [7:0] data_in_2_27_in_data;
	wire [7:0] data_in_2_27_out_data;
	hls_wire #(.WIDTH(8)) data_in_2_27(.in_data(data_in_2_27_in_data), .out_data(data_in_2_27_out_data));

	reg [31:0] data_in_2_29_in_data;
	wire [31:0] data_in_2_29_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_29(.in_data(data_in_2_29_in_data), .out_data(data_in_2_29_out_data));

	reg [7:0] data_in_3_31_in_data;
	wire [7:0] data_in_3_31_out_data;
	hls_wire #(.WIDTH(8)) data_in_3_31(.in_data(data_in_3_31_in_data), .out_data(data_in_3_31_out_data));

	reg [15:0] data_in_3_33_in_data;
	wire [15:0] data_in_3_33_out_data;
	hls_wire #(.WIDTH(16)) data_in_3_33(.in_data(data_in_3_33_in_data), .out_data(data_in_3_33_out_data));

	reg [7:0] data_in_3_35_in_data;
	wire [7:0] data_in_3_35_out_data;
	hls_wire #(.WIDTH(8)) data_in_3_35(.in_data(data_in_3_35_in_data), .out_data(data_in_3_35_out_data));

	reg [7:0] data_in_3_37_in_data;
	wire [7:0] data_in_3_37_out_data;
	hls_wire #(.WIDTH(8)) data_in_3_37(.in_data(data_in_3_37_in_data), .out_data(data_in_3_37_out_data));

	reg [31:0] data_in_3_39_in_data;
	wire [31:0] data_in_3_39_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_39(.in_data(data_in_3_39_in_data), .out_data(data_in_3_39_out_data));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] bb_1_active_in_state_0_in_data;
	wire [0:0] bb_1_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_0(.in_data(bb_1_active_in_state_0_in_data), .out_data(bb_1_active_in_state_0_out_data));

	reg [31:0] bb_1_predecessor_in_state_0_in_data;
	wire [31:0] bb_1_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_0(.in_data(bb_1_predecessor_in_state_0_in_data), .out_data(bb_1_predecessor_in_state_0_out_data));

	reg [0:0] bb_3_active_in_state_0_in_data;
	wire [0:0] bb_3_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_0(.in_data(bb_3_active_in_state_0_in_data), .out_data(bb_3_active_in_state_0_out_data));

	reg [31:0] bb_3_predecessor_in_state_0_in_data;
	wire [31:0] bb_3_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_0(.in_data(bb_3_predecessor_in_state_0_in_data), .out_data(bb_3_predecessor_in_state_0_out_data));

	reg [0:0] bb_4_active_in_state_0_in_data;
	wire [0:0] bb_4_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_0(.in_data(bb_4_active_in_state_0_in_data), .out_data(bb_4_active_in_state_0_out_data));

	reg [31:0] bb_4_predecessor_in_state_0_in_data;
	wire [31:0] bb_4_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_0(.in_data(bb_4_predecessor_in_state_0_in_data), .out_data(bb_4_predecessor_in_state_0_out_data));

	reg [0:0] bb_5_active_in_state_0_in_data;
	wire [0:0] bb_5_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_5_active_in_state_0(.in_data(bb_5_active_in_state_0_in_data), .out_data(bb_5_active_in_state_0_out_data));

	reg [31:0] bb_5_predecessor_in_state_0_in_data;
	wire [31:0] bb_5_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_5_predecessor_in_state_0(.in_data(bb_5_predecessor_in_state_0_in_data), .out_data(bb_5_predecessor_in_state_0_out_data));

	reg [0:0] bb_6_active_in_state_1_in_data;
	wire [0:0] bb_6_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_6_active_in_state_1(.in_data(bb_6_active_in_state_1_in_data), .out_data(bb_6_active_in_state_1_out_data));

	reg [31:0] bb_6_predecessor_in_state_1_in_data;
	wire [31:0] bb_6_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_6_predecessor_in_state_1(.in_data(bb_6_predecessor_in_state_1_in_data), .out_data(bb_6_predecessor_in_state_1_out_data));

	reg [0:0] bb_6_active_in_state_2_in_data;
	wire [0:0] bb_6_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_6_active_in_state_2(.in_data(bb_6_active_in_state_2_in_data), .out_data(bb_6_active_in_state_2_out_data));

	reg [31:0] bb_6_predecessor_in_state_2_in_data;
	wire [31:0] bb_6_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_6_predecessor_in_state_2(.in_data(bb_6_predecessor_in_state_2_in_data), .out_data(bb_6_predecessor_in_state_2_out_data));

	reg [0:0] bb_7_active_in_state_2_in_data;
	wire [0:0] bb_7_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_7_active_in_state_2(.in_data(bb_7_active_in_state_2_in_data), .out_data(bb_7_active_in_state_2_out_data));

	reg [31:0] bb_7_predecessor_in_state_2_in_data;
	wire [31:0] bb_7_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_7_predecessor_in_state_2(.in_data(bb_7_predecessor_in_state_2_in_data), .out_data(bb_7_predecessor_in_state_2_out_data));

	reg [0:0] bb_8_active_in_state_2_in_data;
	wire [0:0] bb_8_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active_in_state_2(.in_data(bb_8_active_in_state_2_in_data), .out_data(bb_8_active_in_state_2_out_data));

	reg [31:0] bb_8_predecessor_in_state_2_in_data;
	wire [31:0] bb_8_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor_in_state_2(.in_data(bb_8_predecessor_in_state_2_in_data), .out_data(bb_8_predecessor_in_state_2_out_data));

	reg [0:0] bb_2_active_in_state_3_in_data;
	wire [0:0] bb_2_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_3(.in_data(bb_2_active_in_state_3_in_data), .out_data(bb_2_active_in_state_3_out_data));

	reg [31:0] bb_2_predecessor_in_state_3_in_data;
	wire [31:0] bb_2_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_3(.in_data(bb_2_predecessor_in_state_3_in_data), .out_data(bb_2_predecessor_in_state_3_out_data));

	reg [0:0] bb_8_active_in_state_3_in_data;
	wire [0:0] bb_8_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active_in_state_3(.in_data(bb_8_active_in_state_3_in_data), .out_data(bb_8_active_in_state_3_out_data));

	reg [31:0] bb_8_predecessor_in_state_3_in_data;
	wire [31:0] bb_8_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor_in_state_3(.in_data(bb_8_predecessor_in_state_3_in_data), .out_data(bb_8_predecessor_in_state_3_out_data));

	reg [0:0] bb_2_active_in_state_4_in_data;
	wire [0:0] bb_2_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_4(.in_data(bb_2_active_in_state_4_in_data), .out_data(bb_2_active_in_state_4_out_data));

	reg [31:0] bb_2_predecessor_in_state_4_in_data;
	wire [31:0] bb_2_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_4(.in_data(bb_2_predecessor_in_state_4_in_data), .out_data(bb_2_predecessor_in_state_4_out_data));

	reg [0:0] bb_2_active_in_state_5_in_data;
	wire [0:0] bb_2_active_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_5(.in_data(bb_2_active_in_state_5_in_data), .out_data(bb_2_active_in_state_5_out_data));

	reg [31:0] bb_2_predecessor_in_state_5_in_data;
	wire [31:0] bb_2_predecessor_in_state_5_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_5(.in_data(bb_2_predecessor_in_state_5_in_data), .out_data(bb_2_predecessor_in_state_5_out_data));

	wire [0:0] andOp_40_in0;
	wire [0:0] andOp_40_in1;
	wire [0:0] andOp_40_out;
	andOp #(.WIDTH(1)) andOp_40(.in0(andOp_40_in0), .in1(andOp_40_in1), .out(andOp_40_out));

	wire [0:0] andOp_41_in0;
	wire [0:0] andOp_41_in1;
	wire [0:0] andOp_41_out;
	andOp #(.WIDTH(1)) andOp_41(.in0(andOp_41_in0), .in1(andOp_41_in1), .out(andOp_41_out));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	wire [0:0] notOp_42_in0;
	wire [0:0] notOp_42_out;
	notOp #(.WIDTH(1)) notOp_42(.in(notOp_42_in0), .out(notOp_42_out));

	wire [0:0] andOp_43_in0;
	wire [0:0] andOp_43_in1;
	wire [0:0] andOp_43_out;
	andOp #(.WIDTH(1)) andOp_43(.in0(andOp_43_in0), .in1(andOp_43_in1), .out(andOp_43_out));

	wire [0:0] andOp_44_in0;
	wire [0:0] andOp_44_in1;
	wire [0:0] andOp_44_out;
	andOp #(.WIDTH(1)) andOp_44(.in0(andOp_44_in0), .in1(andOp_44_in1), .out(andOp_44_out));

	reg [0:0] br_1_happened_in_state_0_in_data;
	wire [0:0] br_1_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened_in_state_0(.in_data(br_1_happened_in_state_0_in_data), .out_data(br_1_happened_in_state_0_out_data));

	wire [0:0] notOp_45_in0;
	wire [0:0] notOp_45_out;
	notOp #(.WIDTH(1)) notOp_45(.in(notOp_45_in0), .out(notOp_45_out));

	wire [0:0] andOp_46_in0;
	wire [0:0] andOp_46_in1;
	wire [0:0] andOp_46_out;
	andOp #(.WIDTH(1)) andOp_46(.in0(andOp_46_in0), .in1(andOp_46_in1), .out(andOp_46_out));

	wire [0:0] andOp_47_in0;
	wire [0:0] andOp_47_in1;
	wire [0:0] andOp_47_out;
	andOp #(.WIDTH(1)) andOp_47(.in0(andOp_47_in0), .in1(andOp_47_in1), .out(andOp_47_out));

	reg [0:0] br_3_happened_in_state_0_in_data;
	wire [0:0] br_3_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_0(.in_data(br_3_happened_in_state_0_in_data), .out_data(br_3_happened_in_state_0_out_data));

	wire [0:0] notOp_48_in0;
	wire [0:0] notOp_48_out;
	notOp #(.WIDTH(1)) notOp_48(.in(notOp_48_in0), .out(notOp_48_out));

	wire [0:0] andOp_49_in0;
	wire [0:0] andOp_49_in1;
	wire [0:0] andOp_49_out;
	andOp #(.WIDTH(1)) andOp_49(.in0(andOp_49_in0), .in1(andOp_49_in1), .out(andOp_49_out));

	wire [0:0] notOp_50_in0;
	wire [0:0] notOp_50_out;
	notOp #(.WIDTH(1)) notOp_50(.in(notOp_50_in0), .out(notOp_50_out));

	wire [0:0] andOp_51_in0;
	wire [0:0] andOp_51_in1;
	wire [0:0] andOp_51_out;
	andOp #(.WIDTH(1)) andOp_51(.in0(andOp_51_in0), .in1(andOp_51_in1), .out(andOp_51_out));

	wire [0:0] andOp_52_in0;
	wire [0:0] andOp_52_in1;
	wire [0:0] andOp_52_out;
	andOp #(.WIDTH(1)) andOp_52(.in0(andOp_52_in0), .in1(andOp_52_in1), .out(andOp_52_out));

	wire [0:0] andOp_53_in0;
	wire [0:0] andOp_53_in1;
	wire [0:0] andOp_53_out;
	andOp #(.WIDTH(1)) andOp_53(.in0(andOp_53_in0), .in1(andOp_53_in1), .out(andOp_53_out));

	reg [0:0] br_4_happened_in_state_0_in_data;
	wire [0:0] br_4_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_0(.in_data(br_4_happened_in_state_0_in_data), .out_data(br_4_happened_in_state_0_out_data));

	wire [0:0] notOp_54_in0;
	wire [0:0] notOp_54_out;
	notOp #(.WIDTH(1)) notOp_54(.in(notOp_54_in0), .out(notOp_54_out));

	wire [0:0] andOp_55_in0;
	wire [0:0] andOp_55_in1;
	wire [0:0] andOp_55_out;
	andOp #(.WIDTH(1)) andOp_55(.in0(andOp_55_in0), .in1(andOp_55_in1), .out(andOp_55_out));

	wire [0:0] andOp_56_in0;
	wire [0:0] andOp_56_in1;
	wire [0:0] andOp_56_out;
	andOp #(.WIDTH(1)) andOp_56(.in0(andOp_56_in0), .in1(andOp_56_in1), .out(andOp_56_out));

	reg [0:0] br_5_happened_in_state_0_in_data;
	wire [0:0] br_5_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_5_happened_in_state_0(.in_data(br_5_happened_in_state_0_in_data), .out_data(br_5_happened_in_state_0_out_data));

	wire [0:0] notOp_57_in0;
	wire [0:0] notOp_57_out;
	notOp #(.WIDTH(1)) notOp_57(.in(notOp_57_in0), .out(notOp_57_out));

	wire [0:0] andOp_58_in0;
	wire [0:0] andOp_58_in1;
	wire [0:0] andOp_58_out;
	andOp #(.WIDTH(1)) andOp_58(.in0(andOp_58_in0), .in1(andOp_58_in1), .out(andOp_58_out));

	wire [0:0] notOp_59_in0;
	wire [0:0] notOp_59_out;
	notOp #(.WIDTH(1)) notOp_59(.in(notOp_59_in0), .out(notOp_59_out));

	wire [0:0] andOp_60_in0;
	wire [0:0] andOp_60_in1;
	wire [0:0] andOp_60_out;
	andOp #(.WIDTH(1)) andOp_60(.in0(andOp_60_in0), .in1(andOp_60_in1), .out(andOp_60_out));

	wire [0:0] andOp_61_in0;
	wire [0:0] andOp_61_in1;
	wire [0:0] andOp_61_out;
	andOp #(.WIDTH(1)) andOp_61(.in0(andOp_61_in0), .in1(andOp_61_in1), .out(andOp_61_out));

	wire [0:0] andOp_62_in0;
	wire [0:0] andOp_62_in1;
	wire [0:0] andOp_62_out;
	andOp #(.WIDTH(1)) andOp_62(.in0(andOp_62_in0), .in1(andOp_62_in1), .out(andOp_62_out));

	reg [0:0] br_6_happened_in_state_1_in_data;
	wire [0:0] br_6_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_6_happened_in_state_1(.in_data(br_6_happened_in_state_1_in_data), .out_data(br_6_happened_in_state_1_out_data));

	wire [0:0] notOp_63_in0;
	wire [0:0] notOp_63_out;
	notOp #(.WIDTH(1)) notOp_63(.in(notOp_63_in0), .out(notOp_63_out));

	wire [0:0] andOp_64_in0;
	wire [0:0] andOp_64_in1;
	wire [0:0] andOp_64_out;
	andOp #(.WIDTH(1)) andOp_64(.in0(andOp_64_in0), .in1(andOp_64_in1), .out(andOp_64_out));

	wire [0:0] andOp_65_in0;
	wire [0:0] andOp_65_in1;
	wire [0:0] andOp_65_out;
	andOp #(.WIDTH(1)) andOp_65(.in0(andOp_65_in0), .in1(andOp_65_in1), .out(andOp_65_out));

	reg [0:0] br_6_happened_in_state_2_in_data;
	wire [0:0] br_6_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_6_happened_in_state_2(.in_data(br_6_happened_in_state_2_in_data), .out_data(br_6_happened_in_state_2_out_data));

	wire [0:0] notOp_66_in0;
	wire [0:0] notOp_66_out;
	notOp #(.WIDTH(1)) notOp_66(.in(notOp_66_in0), .out(notOp_66_out));

	wire [0:0] andOp_67_in0;
	wire [0:0] andOp_67_in1;
	wire [0:0] andOp_67_out;
	andOp #(.WIDTH(1)) andOp_67(.in0(andOp_67_in0), .in1(andOp_67_in1), .out(andOp_67_out));

	wire [0:0] andOp_68_in0;
	wire [0:0] andOp_68_in1;
	wire [0:0] andOp_68_out;
	andOp #(.WIDTH(1)) andOp_68(.in0(andOp_68_in0), .in1(andOp_68_in1), .out(andOp_68_out));

	reg [0:0] br_7_happened_in_state_2_in_data;
	wire [0:0] br_7_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_7_happened_in_state_2(.in_data(br_7_happened_in_state_2_in_data), .out_data(br_7_happened_in_state_2_out_data));

	wire [0:0] notOp_69_in0;
	wire [0:0] notOp_69_out;
	notOp #(.WIDTH(1)) notOp_69(.in(notOp_69_in0), .out(notOp_69_out));

	wire [0:0] andOp_70_in0;
	wire [0:0] andOp_70_in1;
	wire [0:0] andOp_70_out;
	andOp #(.WIDTH(1)) andOp_70(.in0(andOp_70_in0), .in1(andOp_70_in1), .out(andOp_70_out));

	wire [0:0] notOp_71_in0;
	wire [0:0] notOp_71_out;
	notOp #(.WIDTH(1)) notOp_71(.in(notOp_71_in0), .out(notOp_71_out));

	wire [0:0] andOp_72_in0;
	wire [0:0] andOp_72_in1;
	wire [0:0] andOp_72_out;
	andOp #(.WIDTH(1)) andOp_72(.in0(andOp_72_in0), .in1(andOp_72_in1), .out(andOp_72_out));

	wire [0:0] andOp_73_in0;
	wire [0:0] andOp_73_in1;
	wire [0:0] andOp_73_out;
	andOp #(.WIDTH(1)) andOp_73(.in0(andOp_73_in0), .in1(andOp_73_in1), .out(andOp_73_out));

	wire [0:0] andOp_74_in0;
	wire [0:0] andOp_74_in1;
	wire [0:0] andOp_74_out;
	andOp #(.WIDTH(1)) andOp_74(.in0(andOp_74_in0), .in1(andOp_74_in1), .out(andOp_74_out));

	reg [0:0] br_8_happened_in_state_2_in_data;
	wire [0:0] br_8_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_8_happened_in_state_2(.in_data(br_8_happened_in_state_2_in_data), .out_data(br_8_happened_in_state_2_out_data));

	wire [0:0] notOp_75_in0;
	wire [0:0] notOp_75_out;
	notOp #(.WIDTH(1)) notOp_75(.in(notOp_75_in0), .out(notOp_75_out));

	wire [0:0] andOp_76_in0;
	wire [0:0] andOp_76_in1;
	wire [0:0] andOp_76_out;
	andOp #(.WIDTH(1)) andOp_76(.in0(andOp_76_in0), .in1(andOp_76_in1), .out(andOp_76_out));

	wire [0:0] notOp_77_in0;
	wire [0:0] notOp_77_out;
	notOp #(.WIDTH(1)) notOp_77(.in(notOp_77_in0), .out(notOp_77_out));

	wire [0:0] andOp_78_in0;
	wire [0:0] andOp_78_in1;
	wire [0:0] andOp_78_out;
	andOp #(.WIDTH(1)) andOp_78(.in0(andOp_78_in0), .in1(andOp_78_in1), .out(andOp_78_out));

	wire [0:0] andOp_79_in0;
	wire [0:0] andOp_79_in1;
	wire [0:0] andOp_79_out;
	andOp #(.WIDTH(1)) andOp_79(.in0(andOp_79_in0), .in1(andOp_79_in1), .out(andOp_79_out));

	wire [0:0] andOp_80_in0;
	wire [0:0] andOp_80_in1;
	wire [0:0] andOp_80_out;
	andOp #(.WIDTH(1)) andOp_80(.in0(andOp_80_in0), .in1(andOp_80_in1), .out(andOp_80_out));

	reg [0:0] br_8_happened_in_state_3_in_data;
	wire [0:0] br_8_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_8_happened_in_state_3(.in_data(br_8_happened_in_state_3_in_data), .out_data(br_8_happened_in_state_3_out_data));

	wire [0:0] notOp_81_in0;
	wire [0:0] notOp_81_out;
	notOp #(.WIDTH(1)) notOp_81(.in(notOp_81_in0), .out(notOp_81_out));

	wire [0:0] andOp_82_in0;
	wire [0:0] andOp_82_in1;
	wire [0:0] andOp_82_out;
	andOp #(.WIDTH(1)) andOp_82(.in0(andOp_82_in0), .in1(andOp_82_in1), .out(andOp_82_out));

	wire [0:0] notOp_83_in0;
	wire [0:0] notOp_83_out;
	notOp #(.WIDTH(1)) notOp_83(.in(notOp_83_in0), .out(notOp_83_out));

	wire [0:0] andOp_84_in0;
	wire [0:0] andOp_84_in1;
	wire [0:0] andOp_84_out;
	andOp #(.WIDTH(1)) andOp_84(.in0(andOp_84_in0), .in1(andOp_84_in1), .out(andOp_84_out));

	wire [31:0] eq_85_in0;
	wire [31:0] eq_85_in1;
	wire [0:0] eq_85_out;
	eq #(.WIDTH(32)) eq_85(.in0(eq_85_in0), .in1(eq_85_in1), .out(eq_85_out));

	wire [31:0] eq_86_in0;
	wire [31:0] eq_86_in1;
	wire [0:0] eq_86_out;
	eq #(.WIDTH(32)) eq_86(.in0(eq_86_in0), .in1(eq_86_in1), .out(eq_86_out));

	wire [0:0] orOp_87_in0;
	wire [0:0] orOp_87_in1;
	wire [0:0] orOp_87_out;
	orOp #(.WIDTH(1)) orOp_87(.in0(orOp_87_in0), .in1(orOp_87_in1), .out(orOp_87_out));

	wire [31:0] eq_88_in0;
	wire [31:0] eq_88_in1;
	wire [0:0] eq_88_out;
	eq #(.WIDTH(32)) eq_88(.in0(eq_88_in0), .in1(eq_88_in1), .out(eq_88_out));

	wire [0:0] orOp_89_in0;
	wire [0:0] orOp_89_in1;
	wire [0:0] orOp_89_out;
	orOp #(.WIDTH(1)) orOp_89(.in0(orOp_89_in0), .in1(orOp_89_in1), .out(orOp_89_out));

	wire [31:0] eq_90_in0;
	wire [31:0] eq_90_in1;
	wire [0:0] eq_90_out;
	eq #(.WIDTH(32)) eq_90(.in0(eq_90_in0), .in1(eq_90_in1), .out(eq_90_out));

	wire [0:0] orOp_91_in0;
	wire [0:0] orOp_91_in1;
	wire [0:0] orOp_91_out;
	orOp #(.WIDTH(1)) orOp_91(.in0(orOp_91_in0), .in1(orOp_91_in1), .out(orOp_91_out));

	wire [31:0] eq_92_in0;
	wire [31:0] eq_92_in1;
	wire [0:0] eq_92_out;
	eq #(.WIDTH(32)) eq_92(.in0(eq_92_in0), .in1(eq_92_in1), .out(eq_92_out));

	wire [0:0] orOp_93_in0;
	wire [0:0] orOp_93_in1;
	wire [0:0] orOp_93_out;
	orOp #(.WIDTH(1)) orOp_93(.in0(orOp_93_in0), .in1(orOp_93_in1), .out(orOp_93_out));

	wire [31:0] eq_94_in0;
	wire [31:0] eq_94_in1;
	wire [0:0] eq_94_out;
	eq #(.WIDTH(32)) eq_94(.in0(eq_94_in0), .in1(eq_94_in1), .out(eq_94_out));

	wire [31:0] eq_95_in0;
	wire [31:0] eq_95_in1;
	wire [0:0] eq_95_out;
	eq #(.WIDTH(32)) eq_95(.in0(eq_95_in0), .in1(eq_95_in1), .out(eq_95_out));

	wire [31:0] eq_96_in0;
	wire [31:0] eq_96_in1;
	wire [0:0] eq_96_out;
	eq #(.WIDTH(32)) eq_96(.in0(eq_96_in0), .in1(eq_96_in1), .out(eq_96_out));

	wire [0:0] orOp_97_in0;
	wire [0:0] orOp_97_in1;
	wire [0:0] orOp_97_out;
	orOp #(.WIDTH(1)) orOp_97(.in0(orOp_97_in0), .in1(orOp_97_in1), .out(orOp_97_out));

	wire [31:0] eq_98_in0;
	wire [31:0] eq_98_in1;
	wire [0:0] eq_98_out;
	eq #(.WIDTH(32)) eq_98(.in0(eq_98_in0), .in1(eq_98_in1), .out(eq_98_out));

	wire [0:0] orOp_99_in0;
	wire [0:0] orOp_99_in1;
	wire [0:0] orOp_99_out;
	orOp #(.WIDTH(1)) orOp_99(.in0(orOp_99_in0), .in1(orOp_99_in1), .out(orOp_99_out));

	wire [31:0] eq_100_in0;
	wire [31:0] eq_100_in1;
	wire [0:0] eq_100_out;
	eq #(.WIDTH(32)) eq_100(.in0(eq_100_in0), .in1(eq_100_in1), .out(eq_100_out));

	wire [0:0] orOp_101_in0;
	wire [0:0] orOp_101_in1;
	wire [0:0] orOp_101_out;
	orOp #(.WIDTH(1)) orOp_101(.in0(orOp_101_in0), .in1(orOp_101_in1), .out(orOp_101_out));

	wire [31:0] eq_102_in0;
	wire [31:0] eq_102_in1;
	wire [0:0] eq_102_out;
	eq #(.WIDTH(32)) eq_102(.in0(eq_102_in0), .in1(eq_102_in1), .out(eq_102_out));

	wire [31:0] eq_103_in0;
	wire [31:0] eq_103_in1;
	wire [0:0] eq_103_out;
	eq #(.WIDTH(32)) eq_103(.in0(eq_103_in0), .in1(eq_103_in1), .out(eq_103_out));

	wire [31:0] eq_104_in0;
	wire [31:0] eq_104_in1;
	wire [0:0] eq_104_out;
	eq #(.WIDTH(32)) eq_104(.in0(eq_104_in0), .in1(eq_104_in1), .out(eq_104_out));

	wire [31:0] eq_105_in0;
	wire [31:0] eq_105_in1;
	wire [0:0] eq_105_out;
	eq #(.WIDTH(32)) eq_105(.in0(eq_105_in0), .in1(eq_105_in1), .out(eq_105_out));

	wire [31:0] eq_106_in0;
	wire [31:0] eq_106_in1;
	wire [0:0] eq_106_out;
	eq #(.WIDTH(32)) eq_106(.in0(eq_106_in0), .in1(eq_106_in1), .out(eq_106_out));

	wire [0:0] notOp_107_in0;
	wire [0:0] notOp_107_out;
	notOp #(.WIDTH(1)) notOp_107(.in(notOp_107_in0), .out(notOp_107_out));

	wire [0:0] andOp_108_in0;
	wire [0:0] andOp_108_in1;
	wire [0:0] andOp_108_out;
	andOp #(.WIDTH(1)) andOp_108(.in0(andOp_108_in0), .in1(andOp_108_in1), .out(andOp_108_out));

	wire [31:0] eq_109_in0;
	wire [31:0] eq_109_in1;
	wire [0:0] eq_109_out;
	eq #(.WIDTH(32)) eq_109(.in0(eq_109_in0), .in1(eq_109_in1), .out(eq_109_out));

	wire [0:0] notOp_110_in0;
	wire [0:0] notOp_110_out;
	notOp #(.WIDTH(1)) notOp_110(.in(notOp_110_in0), .out(notOp_110_out));

	wire [0:0] andOp_111_in0;
	wire [0:0] andOp_111_in1;
	wire [0:0] andOp_111_out;
	andOp #(.WIDTH(1)) andOp_111(.in0(andOp_111_in0), .in1(andOp_111_in1), .out(andOp_111_out));

	wire [31:0] eq_112_in0;
	wire [31:0] eq_112_in1;
	wire [0:0] eq_112_out;
	eq #(.WIDTH(32)) eq_112(.in0(eq_112_in0), .in1(eq_112_in1), .out(eq_112_out));

	wire [0:0] notOp_113_in0;
	wire [0:0] notOp_113_out;
	notOp #(.WIDTH(1)) notOp_113(.in(notOp_113_in0), .out(notOp_113_out));

	wire [0:0] andOp_114_in0;
	wire [0:0] andOp_114_in1;
	wire [0:0] andOp_114_out;
	andOp #(.WIDTH(1)) andOp_114(.in0(andOp_114_in0), .in1(andOp_114_in1), .out(andOp_114_out));

	wire [31:0] eq_115_in0;
	wire [31:0] eq_115_in1;
	wire [0:0] eq_115_out;
	eq #(.WIDTH(32)) eq_115(.in0(eq_115_in0), .in1(eq_115_in1), .out(eq_115_out));

	wire [0:0] notOp_116_in0;
	wire [0:0] notOp_116_out;
	notOp #(.WIDTH(1)) notOp_116(.in(notOp_116_in0), .out(notOp_116_out));

	wire [0:0] andOp_117_in0;
	wire [0:0] andOp_117_in1;
	wire [0:0] andOp_117_out;
	andOp #(.WIDTH(1)) andOp_117(.in0(andOp_117_in0), .in1(andOp_117_in1), .out(andOp_117_out));

	wire [31:0] eq_118_in0;
	wire [31:0] eq_118_in1;
	wire [0:0] eq_118_out;
	eq #(.WIDTH(32)) eq_118(.in0(eq_118_in0), .in1(eq_118_in1), .out(eq_118_out));

	wire [31:0] eq_119_in0;
	wire [31:0] eq_119_in1;
	wire [0:0] eq_119_out;
	eq #(.WIDTH(32)) eq_119(.in0(eq_119_in0), .in1(eq_119_in1), .out(eq_119_out));

	wire [31:0] eq_120_in0;
	wire [31:0] eq_120_in1;
	wire [0:0] eq_120_out;
	eq #(.WIDTH(32)) eq_120(.in0(eq_120_in0), .in1(eq_120_in1), .out(eq_120_out));

	wire [0:0] notOp_121_in0;
	wire [0:0] notOp_121_out;
	notOp #(.WIDTH(1)) notOp_121(.in(notOp_121_in0), .out(notOp_121_out));

	wire [0:0] andOp_122_in0;
	wire [0:0] andOp_122_in1;
	wire [0:0] andOp_122_out;
	andOp #(.WIDTH(1)) andOp_122(.in0(andOp_122_in0), .in1(andOp_122_in1), .out(andOp_122_out));

	wire [31:0] eq_123_in0;
	wire [31:0] eq_123_in1;
	wire [0:0] eq_123_out;
	eq #(.WIDTH(32)) eq_123(.in0(eq_123_in0), .in1(eq_123_in1), .out(eq_123_out));

	wire [0:0] notOp_124_in0;
	wire [0:0] notOp_124_out;
	notOp #(.WIDTH(1)) notOp_124(.in(notOp_124_in0), .out(notOp_124_out));

	wire [0:0] andOp_125_in0;
	wire [0:0] andOp_125_in1;
	wire [0:0] andOp_125_out;
	andOp #(.WIDTH(1)) andOp_125(.in0(andOp_125_in0), .in1(andOp_125_in1), .out(andOp_125_out));

	wire [31:0] eq_126_in0;
	wire [31:0] eq_126_in1;
	wire [0:0] eq_126_out;
	eq #(.WIDTH(32)) eq_126(.in0(eq_126_in0), .in1(eq_126_in1), .out(eq_126_out));

	wire [0:0] notOp_127_in0;
	wire [0:0] notOp_127_out;
	notOp #(.WIDTH(1)) notOp_127(.in(notOp_127_in0), .out(notOp_127_out));

	wire [0:0] andOp_128_in0;
	wire [0:0] andOp_128_in1;
	wire [0:0] andOp_128_out;
	andOp #(.WIDTH(1)) andOp_128(.in0(andOp_128_in0), .in1(andOp_128_in1), .out(andOp_128_out));

	wire [31:0] eq_129_in0;
	wire [31:0] eq_129_in1;
	wire [0:0] eq_129_out;
	eq #(.WIDTH(32)) eq_129(.in0(eq_129_in0), .in1(eq_129_in1), .out(eq_129_out));

	wire [31:0] eq_130_in0;
	wire [31:0] eq_130_in1;
	wire [0:0] eq_130_out;
	eq #(.WIDTH(32)) eq_130(.in0(eq_130_in0), .in1(eq_130_in1), .out(eq_130_out));

	wire [31:0] eq_131_in0;
	wire [31:0] eq_131_in1;
	wire [0:0] eq_131_out;
	eq #(.WIDTH(32)) eq_131(.in0(eq_131_in0), .in1(eq_131_in1), .out(eq_131_out));

	wire [0:0] andOp_132_in0;
	wire [0:0] andOp_132_in1;
	wire [0:0] andOp_132_out;
	andOp #(.WIDTH(1)) andOp_132(.in0(andOp_132_in0), .in1(andOp_132_in1), .out(andOp_132_out));

	wire [0:0] andOp_133_in0;
	wire [0:0] andOp_133_in1;
	wire [0:0] andOp_133_out;
	andOp #(.WIDTH(1)) andOp_133(.in0(andOp_133_in0), .in1(andOp_133_in1), .out(andOp_133_out));

	wire [0:0] andOp_134_in0;
	wire [0:0] andOp_134_in1;
	wire [0:0] andOp_134_out;
	andOp #(.WIDTH(1)) andOp_134(.in0(andOp_134_in0), .in1(andOp_134_in1), .out(andOp_134_out));

	wire [0:0] andOp_135_in0;
	wire [0:0] andOp_135_in1;
	wire [0:0] andOp_135_out;
	andOp #(.WIDTH(1)) andOp_135(.in0(andOp_135_in0), .in1(andOp_135_in1), .out(andOp_135_out));

	reg [7:0] tmp_output_136_in_data;
	wire [7:0] tmp_output_136_out_data;
	hls_wire #(.WIDTH(8)) tmp_output_136(.in_data(tmp_output_136_in_data), .out_data(tmp_output_136_out_data));

	wire [31:0] eq_137_in0;
	wire [31:0] eq_137_in1;
	wire [0:0] eq_137_out;
	eq #(.WIDTH(32)) eq_137(.in0(eq_137_in0), .in1(eq_137_in1), .out(eq_137_out));

	wire [31:0] eq_138_in0;
	wire [31:0] eq_138_in1;
	wire [0:0] eq_138_out;
	eq #(.WIDTH(32)) eq_138(.in0(eq_138_in0), .in1(eq_138_in1), .out(eq_138_out));

	wire [31:0] eq_139_in0;
	wire [31:0] eq_139_in1;
	wire [0:0] eq_139_out;
	eq #(.WIDTH(32)) eq_139(.in0(eq_139_in0), .in1(eq_139_in1), .out(eq_139_out));

	wire [31:0] eq_140_in0;
	wire [31:0] eq_140_in1;
	wire [0:0] eq_140_out;
	eq #(.WIDTH(32)) eq_140(.in0(eq_140_in0), .in1(eq_140_in1), .out(eq_140_out));

	wire [0:0] andOp_141_in0;
	wire [0:0] andOp_141_in1;
	wire [0:0] andOp_141_out;
	andOp #(.WIDTH(1)) andOp_141(.in0(andOp_141_in0), .in1(andOp_141_in1), .out(andOp_141_out));

	reg [15:0] tmp_output_142_in_data;
	wire [15:0] tmp_output_142_out_data;
	hls_wire #(.WIDTH(16)) tmp_output_142(.in_data(tmp_output_142_in_data), .out_data(tmp_output_142_out_data));

	wire [31:0] eq_143_in0;
	wire [31:0] eq_143_in1;
	wire [0:0] eq_143_out;
	eq #(.WIDTH(32)) eq_143(.in0(eq_143_in0), .in1(eq_143_in1), .out(eq_143_out));

	wire [31:0] eq_144_in0;
	wire [31:0] eq_144_in1;
	wire [0:0] eq_144_out;
	eq #(.WIDTH(32)) eq_144(.in0(eq_144_in0), .in1(eq_144_in1), .out(eq_144_out));

	wire [31:0] eq_145_in0;
	wire [31:0] eq_145_in1;
	wire [0:0] eq_145_out;
	eq #(.WIDTH(32)) eq_145(.in0(eq_145_in0), .in1(eq_145_in1), .out(eq_145_out));

	wire [31:0] eq_146_in0;
	wire [31:0] eq_146_in1;
	wire [0:0] eq_146_out;
	eq #(.WIDTH(32)) eq_146(.in0(eq_146_in0), .in1(eq_146_in1), .out(eq_146_out));

	wire [0:0] andOp_147_in0;
	wire [0:0] andOp_147_in1;
	wire [0:0] andOp_147_out;
	andOp #(.WIDTH(1)) andOp_147(.in0(andOp_147_in0), .in1(andOp_147_in1), .out(andOp_147_out));

	wire [0:0] andOp_148_in0;
	wire [0:0] andOp_148_in1;
	wire [0:0] andOp_148_out;
	andOp #(.WIDTH(1)) andOp_148(.in0(andOp_148_in0), .in1(andOp_148_in1), .out(andOp_148_out));

	wire [0:0] andOp_149_in0;
	wire [0:0] andOp_149_in1;
	wire [0:0] andOp_149_out;
	andOp #(.WIDTH(1)) andOp_149(.in0(andOp_149_in0), .in1(andOp_149_in1), .out(andOp_149_out));

	wire [0:0] andOp_150_in0;
	wire [0:0] andOp_150_in1;
	wire [0:0] andOp_150_out;
	andOp #(.WIDTH(1)) andOp_150(.in0(andOp_150_in0), .in1(andOp_150_in1), .out(andOp_150_out));

	wire [0:0] andOp_151_in0;
	wire [0:0] andOp_151_in1;
	wire [0:0] andOp_151_out;
	andOp #(.WIDTH(1)) andOp_151(.in0(andOp_151_in0), .in1(andOp_151_in1), .out(andOp_151_out));

	wire [0:0] andOp_152_in0;
	wire [0:0] andOp_152_in1;
	wire [0:0] andOp_152_out;
	andOp #(.WIDTH(1)) andOp_152(.in0(andOp_152_in0), .in1(andOp_152_in1), .out(andOp_152_out));

	wire [0:0] andOp_153_in0;
	wire [0:0] andOp_153_in1;
	wire [0:0] andOp_153_out;
	andOp #(.WIDTH(1)) andOp_153(.in0(andOp_153_in0), .in1(andOp_153_in1), .out(andOp_153_out));

	reg [31:0] tmp_output_154_in_data;
	wire [31:0] tmp_output_154_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_154(.in_data(tmp_output_154_in_data), .out_data(tmp_output_154_out_data));

	wire [31:0] eq_155_in0;
	wire [31:0] eq_155_in1;
	wire [0:0] eq_155_out;
	eq #(.WIDTH(32)) eq_155(.in0(eq_155_in0), .in1(eq_155_in1), .out(eq_155_out));

	wire [31:0] eq_156_in0;
	wire [31:0] eq_156_in1;
	wire [0:0] eq_156_out;
	eq #(.WIDTH(32)) eq_156(.in0(eq_156_in0), .in1(eq_156_in1), .out(eq_156_out));

	wire [0:0] andOp_157_in0;
	wire [0:0] andOp_157_in1;
	wire [0:0] andOp_157_out;
	andOp #(.WIDTH(1)) andOp_157(.in0(andOp_157_in0), .in1(andOp_157_in1), .out(andOp_157_out));

	wire [0:0] andOp_158_in0;
	wire [0:0] andOp_158_in1;
	wire [0:0] andOp_158_out;
	andOp #(.WIDTH(1)) andOp_158(.in0(andOp_158_in0), .in1(andOp_158_in1), .out(andOp_158_out));

	wire [0:0] andOp_159_in0;
	wire [0:0] andOp_159_in1;
	wire [0:0] andOp_159_out;
	andOp #(.WIDTH(1)) andOp_159(.in0(andOp_159_in0), .in1(andOp_159_in1), .out(andOp_159_out));

	wire [0:0] andOp_160_in0;
	wire [0:0] andOp_160_in1;
	wire [0:0] andOp_160_out;
	andOp #(.WIDTH(1)) andOp_160(.in0(andOp_160_in0), .in1(andOp_160_in1), .out(andOp_160_out));

	wire [0:0] andOp_161_in0;
	wire [0:0] andOp_161_in1;
	wire [0:0] andOp_161_out;
	andOp #(.WIDTH(1)) andOp_161(.in0(andOp_161_in0), .in1(andOp_161_in1), .out(andOp_161_out));

	wire [0:0] andOp_162_in0;
	wire [0:0] andOp_162_in1;
	wire [0:0] andOp_162_out;
	andOp #(.WIDTH(1)) andOp_162(.in0(andOp_162_in0), .in1(andOp_162_in1), .out(andOp_162_out));

	wire [7:0] concat_163_in0;
	wire [7:0] concat_163_in1;
	wire [15:0] concat_163_out;
	concat #(.IN0_WIDTH(8), .IN1_WIDTH(8)) concat_163(.in0(concat_163_in0), .in1(concat_163_in1), .out(concat_163_out));

	wire [31:0] concat_164_in0;
	wire [31:0] concat_164_in1;
	wire [63:0] concat_164_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_164(.in0(concat_164_in0), .in1(concat_164_in1), .out(concat_164_out));

	wire [0:0] andOp_165_in0;
	wire [0:0] andOp_165_in1;
	wire [0:0] andOp_165_out;
	andOp #(.WIDTH(1)) andOp_165(.in0(andOp_165_in0), .in1(andOp_165_in1), .out(andOp_165_out));

	wire [0:0] andOp_166_in0;
	wire [0:0] andOp_166_in1;
	wire [0:0] andOp_166_out;
	andOp #(.WIDTH(1)) andOp_166(.in0(andOp_166_in0), .in1(andOp_166_in1), .out(andOp_166_out));

	wire [0:0] andOp_167_in0;
	wire [0:0] andOp_167_in1;
	wire [0:0] andOp_167_out;
	andOp #(.WIDTH(1)) andOp_167(.in0(andOp_167_in0), .in1(andOp_167_in1), .out(andOp_167_out));

	wire [0:0] andOp_168_in0;
	wire [0:0] andOp_168_in1;
	wire [0:0] andOp_168_out;
	andOp #(.WIDTH(1)) andOp_168(.in0(andOp_168_in0), .in1(andOp_168_in1), .out(andOp_168_out));

	wire [0:0] andOp_169_in0;
	wire [0:0] andOp_169_in1;
	wire [0:0] andOp_169_out;
	andOp #(.WIDTH(1)) andOp_169(.in0(andOp_169_in0), .in1(andOp_169_in1), .out(andOp_169_out));

	wire [0:0] andOp_170_in0;
	wire [0:0] andOp_170_in1;
	wire [0:0] andOp_170_out;
	andOp #(.WIDTH(1)) andOp_170(.in0(andOp_170_in0), .in1(andOp_170_in1), .out(andOp_170_out));

	wire [0:0] andOp_171_in0;
	wire [0:0] andOp_171_in1;
	wire [0:0] andOp_171_out;
	andOp #(.WIDTH(1)) andOp_171(.in0(andOp_171_in0), .in1(andOp_171_in1), .out(andOp_171_out));

	wire [0:0] andOp_172_in0;
	wire [0:0] andOp_172_in1;
	wire [0:0] andOp_172_out;
	andOp #(.WIDTH(1)) andOp_172(.in0(andOp_172_in0), .in1(andOp_172_in1), .out(andOp_172_out));

	wire [0:0] andOp_173_in0;
	wire [0:0] andOp_173_in1;
	wire [0:0] andOp_173_out;
	andOp #(.WIDTH(1)) andOp_173(.in0(andOp_173_in0), .in1(andOp_173_in1), .out(andOp_173_out));

	wire [0:0] andOp_174_in0;
	wire [0:0] andOp_174_in1;
	wire [0:0] andOp_174_out;
	andOp #(.WIDTH(1)) andOp_174(.in0(andOp_174_in0), .in1(andOp_174_in1), .out(andOp_174_out));

	wire [0:0] andOp_175_in0;
	wire [0:0] andOp_175_in1;
	wire [0:0] andOp_175_out;
	andOp #(.WIDTH(1)) andOp_175(.in0(andOp_175_in0), .in1(andOp_175_in1), .out(andOp_175_out));

	wire [0:0] andOp_176_in0;
	wire [0:0] andOp_176_in1;
	wire [0:0] andOp_176_out;
	andOp #(.WIDTH(1)) andOp_176(.in0(andOp_176_in0), .in1(andOp_176_in1), .out(andOp_176_out));

	wire [0:0] andOp_177_in0;
	wire [0:0] andOp_177_in1;
	wire [0:0] andOp_177_out;
	andOp #(.WIDTH(1)) andOp_177(.in0(andOp_177_in0), .in1(andOp_177_in1), .out(andOp_177_out));

	wire [0:0] andOp_178_in0;
	wire [0:0] andOp_178_in1;
	wire [0:0] andOp_178_out;
	andOp #(.WIDTH(1)) andOp_178(.in0(andOp_178_in0), .in1(andOp_178_in1), .out(andOp_178_out));

	wire [0:0] andOp_179_in0;
	wire [0:0] andOp_179_in1;
	wire [0:0] andOp_179_out;
	andOp #(.WIDTH(1)) andOp_179(.in0(andOp_179_in0), .in1(andOp_179_in1), .out(andOp_179_out));

	wire [0:0] andOp_180_in0;
	wire [0:0] andOp_180_in1;
	wire [0:0] andOp_180_out;
	andOp #(.WIDTH(1)) andOp_180(.in0(andOp_180_in0), .in1(andOp_180_in1), .out(andOp_180_out));

	wire [0:0] andOp_181_in0;
	wire [0:0] andOp_181_in1;
	wire [0:0] andOp_181_out;
	andOp #(.WIDTH(1)) andOp_181(.in0(andOp_181_in0), .in1(andOp_181_in1), .out(andOp_181_out));

	wire [0:0] andOp_182_in0;
	wire [0:0] andOp_182_in1;
	wire [0:0] andOp_182_out;
	andOp #(.WIDTH(1)) andOp_182(.in0(andOp_182_in0), .in1(andOp_182_in1), .out(andOp_182_out));

	wire [0:0] andOp_183_in0;
	wire [0:0] andOp_183_in1;
	wire [0:0] andOp_183_out;
	andOp #(.WIDTH(1)) andOp_183(.in0(andOp_183_in0), .in1(andOp_183_in1), .out(andOp_183_out));

	wire [0:0] andOp_184_in0;
	wire [0:0] andOp_184_in1;
	wire [0:0] andOp_184_out;
	andOp #(.WIDTH(1)) andOp_184(.in0(andOp_184_in0), .in1(andOp_184_in1), .out(andOp_184_out));

	wire [0:0] notOp_185_in0;
	wire [0:0] notOp_185_out;
	notOp #(.WIDTH(1)) notOp_185(.in(notOp_185_in0), .out(notOp_185_out));

	wire [0:0] andOp_186_in0;
	wire [0:0] andOp_186_in1;
	wire [0:0] andOp_186_out;
	andOp #(.WIDTH(1)) andOp_186(.in0(andOp_186_in0), .in1(andOp_186_in1), .out(andOp_186_out));

	wire [0:0] notOp_187_in0;
	wire [0:0] notOp_187_out;
	notOp #(.WIDTH(1)) notOp_187(.in(notOp_187_in0), .out(notOp_187_out));

	wire [0:0] andOp_188_in0;
	wire [0:0] andOp_188_in1;
	wire [0:0] andOp_188_out;
	andOp #(.WIDTH(1)) andOp_188(.in0(andOp_188_in0), .in1(andOp_188_in1), .out(andOp_188_out));

	wire [0:0] notOp_189_in0;
	wire [0:0] notOp_189_out;
	notOp #(.WIDTH(1)) notOp_189(.in(notOp_189_in0), .out(notOp_189_out));

	wire [0:0] andOp_190_in0;
	wire [0:0] andOp_190_in1;
	wire [0:0] andOp_190_out;
	andOp #(.WIDTH(1)) andOp_190(.in0(andOp_190_in0), .in1(andOp_190_in1), .out(andOp_190_out));

	wire [0:0] notOp_191_in0;
	wire [0:0] notOp_191_out;
	notOp #(.WIDTH(1)) notOp_191(.in(notOp_191_in0), .out(notOp_191_out));

	wire [0:0] andOp_192_in0;
	wire [0:0] andOp_192_in1;
	wire [0:0] andOp_192_out;
	andOp #(.WIDTH(1)) andOp_192(.in0(andOp_192_in0), .in1(andOp_192_in1), .out(andOp_192_out));

	wire [0:0] notOp_193_in0;
	wire [0:0] notOp_193_out;
	notOp #(.WIDTH(1)) notOp_193(.in(notOp_193_in0), .out(notOp_193_out));

	wire [0:0] andOp_194_in0;
	wire [0:0] andOp_194_in1;
	wire [0:0] andOp_194_out;
	andOp #(.WIDTH(1)) andOp_194(.in0(andOp_194_in0), .in1(andOp_194_in1), .out(andOp_194_out));

	wire [0:0] notOp_195_in0;
	wire [0:0] notOp_195_out;
	notOp #(.WIDTH(1)) notOp_195(.in(notOp_195_in0), .out(notOp_195_out));

	wire [0:0] andOp_196_in0;
	wire [0:0] andOp_196_in1;
	wire [0:0] andOp_196_out;
	andOp #(.WIDTH(1)) andOp_196(.in0(andOp_196_in0), .in1(andOp_196_in1), .out(andOp_196_out));

	wire [0:0] notOp_197_in0;
	wire [0:0] notOp_197_out;
	notOp #(.WIDTH(1)) notOp_197(.in(notOp_197_in0), .out(notOp_197_out));

	wire [0:0] andOp_198_in0;
	wire [0:0] andOp_198_in1;
	wire [0:0] andOp_198_out;
	andOp #(.WIDTH(1)) andOp_198(.in0(andOp_198_in0), .in1(andOp_198_in1), .out(andOp_198_out));

	wire [0:0] notOp_199_in0;
	wire [0:0] notOp_199_out;
	notOp #(.WIDTH(1)) notOp_199(.in(notOp_199_in0), .out(notOp_199_out));

	wire [0:0] andOp_200_in0;
	wire [0:0] andOp_200_in1;
	wire [0:0] andOp_200_out;
	andOp #(.WIDTH(1)) andOp_200(.in0(andOp_200_in0), .in1(andOp_200_in1), .out(andOp_200_out));

	wire [0:0] notOp_201_in0;
	wire [0:0] notOp_201_out;
	notOp #(.WIDTH(1)) notOp_201(.in(notOp_201_in0), .out(notOp_201_out));

	wire [0:0] andOp_202_in0;
	wire [0:0] andOp_202_in1;
	wire [0:0] andOp_202_out;
	andOp #(.WIDTH(1)) andOp_202(.in0(andOp_202_in0), .in1(andOp_202_in1), .out(andOp_202_out));

	wire [0:0] notOp_203_in0;
	wire [0:0] notOp_203_out;
	notOp #(.WIDTH(1)) notOp_203(.in(notOp_203_in0), .out(notOp_203_out));

	wire [0:0] andOp_204_in0;
	wire [0:0] andOp_204_in1;
	wire [0:0] andOp_204_out;
	andOp #(.WIDTH(1)) andOp_204(.in0(andOp_204_in0), .in1(andOp_204_in1), .out(andOp_204_out));

	wire [31:0] eq_205_in0;
	wire [31:0] eq_205_in1;
	wire [0:0] eq_205_out;
	eq #(.WIDTH(32)) eq_205(.in0(eq_205_in0), .in1(eq_205_in1), .out(eq_205_out));

	wire [31:0] eq_206_in0;
	wire [31:0] eq_206_in1;
	wire [0:0] eq_206_out;
	eq #(.WIDTH(32)) eq_206(.in0(eq_206_in0), .in1(eq_206_in1), .out(eq_206_out));

	wire [0:0] andOp_207_in0;
	wire [0:0] andOp_207_in1;
	wire [0:0] andOp_207_out;
	andOp #(.WIDTH(1)) andOp_207(.in0(andOp_207_in0), .in1(andOp_207_in1), .out(andOp_207_out));

	wire [0:0] andOp_208_in0;
	wire [0:0] andOp_208_in1;
	wire [0:0] andOp_208_out;
	andOp #(.WIDTH(1)) andOp_208(.in0(andOp_208_in0), .in1(andOp_208_in1), .out(andOp_208_out));

	wire [0:0] andOp_209_in0;
	wire [0:0] andOp_209_in1;
	wire [0:0] andOp_209_out;
	andOp #(.WIDTH(1)) andOp_209(.in0(andOp_209_in0), .in1(andOp_209_in1), .out(andOp_209_out));

	wire [31:0] eq_210_in0;
	wire [31:0] eq_210_in1;
	wire [0:0] eq_210_out;
	eq #(.WIDTH(32)) eq_210(.in0(eq_210_in0), .in1(eq_210_in1), .out(eq_210_out));

	wire [31:0] eq_211_in0;
	wire [31:0] eq_211_in1;
	wire [0:0] eq_211_out;
	eq #(.WIDTH(32)) eq_211(.in0(eq_211_in0), .in1(eq_211_in1), .out(eq_211_out));

	wire [31:0] eq_212_in0;
	wire [31:0] eq_212_in1;
	wire [0:0] eq_212_out;
	eq #(.WIDTH(32)) eq_212(.in0(eq_212_in0), .in1(eq_212_in1), .out(eq_212_out));

	wire [31:0] eq_213_in0;
	wire [31:0] eq_213_in1;
	wire [0:0] eq_213_out;
	eq #(.WIDTH(32)) eq_213(.in0(eq_213_in0), .in1(eq_213_in1), .out(eq_213_out));

	wire [0:0] andOp_214_in0;
	wire [0:0] andOp_214_in1;
	wire [0:0] andOp_214_out;
	andOp #(.WIDTH(1)) andOp_214(.in0(andOp_214_in0), .in1(andOp_214_in1), .out(andOp_214_out));

	wire [0:0] andOp_215_in0;
	wire [0:0] andOp_215_in1;
	wire [0:0] andOp_215_out;
	andOp #(.WIDTH(1)) andOp_215(.in0(andOp_215_in0), .in1(andOp_215_in1), .out(andOp_215_out));

	wire [31:0] eq_216_in0;
	wire [31:0] eq_216_in1;
	wire [0:0] eq_216_out;
	eq #(.WIDTH(32)) eq_216(.in0(eq_216_in0), .in1(eq_216_in1), .out(eq_216_out));

	wire [31:0] eq_217_in0;
	wire [31:0] eq_217_in1;
	wire [0:0] eq_217_out;
	eq #(.WIDTH(32)) eq_217(.in0(eq_217_in0), .in1(eq_217_in1), .out(eq_217_out));

	wire [31:0] eq_218_in0;
	wire [31:0] eq_218_in1;
	wire [0:0] eq_218_out;
	eq #(.WIDTH(32)) eq_218(.in0(eq_218_in0), .in1(eq_218_in1), .out(eq_218_out));

	wire [31:0] eq_219_in0;
	wire [31:0] eq_219_in1;
	wire [0:0] eq_219_out;
	eq #(.WIDTH(32)) eq_219(.in0(eq_219_in0), .in1(eq_219_in1), .out(eq_219_out));

	wire [31:0] eq_220_in0;
	wire [31:0] eq_220_in1;
	wire [0:0] eq_220_out;
	eq #(.WIDTH(32)) eq_220(.in0(eq_220_in0), .in1(eq_220_in1), .out(eq_220_out));

	wire [31:0] eq_221_in0;
	wire [31:0] eq_221_in1;
	wire [0:0] eq_221_out;
	eq #(.WIDTH(32)) eq_221(.in0(eq_221_in0), .in1(eq_221_in1), .out(eq_221_out));

	// End Functional Units

	reg [7:0] data_store_0_0;
	reg [15:0] data_store_0_2;
	reg [7:0] data_store_0_4;
	reg [7:0] data_store_0_6;
	reg [31:0] data_store_0_8;
	reg [7:0] data_store_1_10;
	reg [15:0] data_store_1_12;
	reg [7:0] data_store_1_14;
	reg [7:0] data_store_1_16;
	reg [31:0] data_store_1_18;
	reg [7:0] data_store_2_20;
	reg [15:0] data_store_2_22;
	reg [7:0] data_store_2_24;
	reg [7:0] data_store_2_26;
	reg [31:0] data_store_2_28;
	reg [7:0] data_store_3_30;
	reg [15:0] data_store_3_32;
	reg [7:0] data_store_3_34;
	reg [7:0] data_store_3_36;
	reg [31:0] data_store_3_38;
	reg [31:0] global_state;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_3_last_state;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;
	reg [31:0] state_4_last_state;
	reg [31:0] state_5_entry_BB_reg;
	reg [0:0] state_5_is_active;
	reg [31:0] state_5_last_BB_reg;
	reg [31:0] state_5_last_state;

	// controller for add_add_22.add_in0_add_22
	// controller for add_add_22.add_in1_add_22
	// Insensitive connections
	assign add_in0_add_22 = sgt_out_sext_21;
	assign add_in1_add_22 = 32'd1;
	// controller for andOp_108.andOp_108_in0
	// controller for andOp_108.andOp_108_in1
	// Insensitive connections
	assign andOp_108_in0 = notOp_107_out;
	assign andOp_108_in1 = andOp_53_out;
	// controller for andOp_111.andOp_111_in0
	// controller for andOp_111.andOp_111_in1
	// Insensitive connections
	assign andOp_111_in0 = notOp_110_out;
	assign andOp_111_in1 = andOp_41_out;
	// controller for andOp_114.andOp_114_in0
	// controller for andOp_114.andOp_114_in1
	// Insensitive connections
	assign andOp_114_in0 = notOp_113_out;
	assign andOp_114_in1 = andOp_51_out;
	// controller for andOp_117.andOp_117_in0
	// controller for andOp_117.andOp_117_in1
	// Insensitive connections
	assign andOp_117_in0 = notOp_116_out;
	assign andOp_117_in1 = andOp_44_out;
	// controller for andOp_122.andOp_122_in0
	// controller for andOp_122.andOp_122_in1
	// Insensitive connections
	assign andOp_122_in0 = notOp_121_out;
	assign andOp_122_in1 = andOp_62_out;
	// controller for andOp_125.andOp_125_in0
	// controller for andOp_125.andOp_125_in1
	// Insensitive connections
	assign andOp_125_in0 = notOp_124_out;
	assign andOp_125_in1 = andOp_72_out;
	// controller for andOp_128.andOp_128_in0
	// controller for andOp_128.andOp_128_in1
	// Insensitive connections
	assign andOp_128_in0 = notOp_127_out;
	assign andOp_128_in1 = andOp_78_out;
	// controller for andOp_132.andOp_132_in0
	// controller for andOp_132.andOp_132_in1
	// Insensitive connections
	assign andOp_132_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_132_in1 = state_0_is_active;
	// controller for andOp_133.andOp_133_in0
	// controller for andOp_133.andOp_133_in1
	// Insensitive connections
	assign andOp_133_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_133_in1 = state_0_is_active;
	// controller for andOp_134.andOp_134_in0
	// controller for andOp_134.andOp_134_in1
	// Insensitive connections
	assign andOp_134_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_134_in1 = state_0_is_active;
	// controller for andOp_135.andOp_135_in0
	// controller for andOp_135.andOp_135_in1
	// Insensitive connections
	assign andOp_135_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_135_in1 = state_0_is_active;
	// controller for andOp_141.andOp_141_in0
	// controller for andOp_141.andOp_141_in1
	// Insensitive connections
	assign andOp_141_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_141_in1 = state_0_is_active;
	// controller for andOp_147.andOp_147_in0
	// controller for andOp_147.andOp_147_in1
	// Insensitive connections
	assign andOp_147_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_147_in1 = state_0_is_active;
	// controller for andOp_148.andOp_148_in0
	// controller for andOp_148.andOp_148_in1
	// Insensitive connections
	assign andOp_148_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_148_in1 = state_0_is_active;
	// controller for andOp_149.andOp_149_in0
	// controller for andOp_149.andOp_149_in1
	// Insensitive connections
	assign andOp_149_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_149_in1 = state_0_is_active;
	// controller for andOp_150.andOp_150_in0
	// controller for andOp_150.andOp_150_in1
	// Insensitive connections
	assign andOp_150_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_150_in1 = state_0_is_active;
	// controller for andOp_151.andOp_151_in0
	// controller for andOp_151.andOp_151_in1
	// Insensitive connections
	assign andOp_151_in0 = bb_7_active_in_state_2_out_data;
	assign andOp_151_in1 = state_2_is_active;
	// controller for andOp_152.andOp_152_in0
	// controller for andOp_152.andOp_152_in1
	// Insensitive connections
	assign andOp_152_in0 = bb_7_active_in_state_2_out_data;
	assign andOp_152_in1 = state_2_is_active;
	// controller for andOp_153.andOp_153_in0
	// controller for andOp_153.andOp_153_in1
	// Insensitive connections
	assign andOp_153_in0 = bb_7_active_in_state_2_out_data;
	assign andOp_153_in1 = state_2_is_active;
	// controller for andOp_157.andOp_157_in0
	// controller for andOp_157.andOp_157_in1
	// Insensitive connections
	assign andOp_157_in0 = bb_7_active_in_state_2_out_data;
	assign andOp_157_in1 = state_2_is_active;
	// controller for andOp_158.andOp_158_in0
	// controller for andOp_158.andOp_158_in1
	// Insensitive connections
	assign andOp_158_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_158_in1 = state_3_is_active;
	// controller for andOp_159.andOp_159_in0
	// controller for andOp_159.andOp_159_in1
	// Insensitive connections
	assign andOp_159_in0 = bb_2_active_in_state_4_out_data;
	assign andOp_159_in1 = state_4_is_active;
	// controller for andOp_160.andOp_160_in0
	// controller for andOp_160.andOp_160_in1
	// Insensitive connections
	assign andOp_160_in0 = bb_2_active_in_state_4_out_data;
	assign andOp_160_in1 = state_4_is_active;
	// controller for andOp_161.andOp_161_in0
	// controller for andOp_161.andOp_161_in1
	// Insensitive connections
	assign andOp_161_in0 = bb_2_active_in_state_4_out_data;
	assign andOp_161_in1 = state_4_is_active;
	// controller for andOp_162.andOp_162_in0
	// controller for andOp_162.andOp_162_in1
	// Insensitive connections
	assign andOp_162_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_162_in1 = state_0_is_active;
	// controller for andOp_165.andOp_165_in0
	// controller for andOp_165.andOp_165_in1
	// Insensitive connections
	assign andOp_165_in0 = bb_5_active_in_state_0_out_data;
	assign andOp_165_in1 = state_0_is_active;
	// controller for andOp_166.andOp_166_in0
	// controller for andOp_166.andOp_166_in1
	// Insensitive connections
	assign andOp_166_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_166_in1 = state_0_is_active;
	// controller for andOp_167.andOp_167_in0
	// controller for andOp_167.andOp_167_in1
	// Insensitive connections
	assign andOp_167_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_167_in1 = state_0_is_active;
	// controller for andOp_168.andOp_168_in0
	// controller for andOp_168.andOp_168_in1
	// Insensitive connections
	assign andOp_168_in0 = bb_5_active_in_state_0_out_data;
	assign andOp_168_in1 = state_0_is_active;
	// controller for andOp_169.andOp_169_in0
	// controller for andOp_169.andOp_169_in1
	// Insensitive connections
	assign andOp_169_in0 = bb_5_active_in_state_0_out_data;
	assign andOp_169_in1 = state_0_is_active;
	// controller for andOp_170.andOp_170_in0
	// controller for andOp_170.andOp_170_in1
	// Insensitive connections
	assign andOp_170_in0 = bb_6_active_in_state_1_out_data;
	assign andOp_170_in1 = state_1_is_active;
	// controller for andOp_171.andOp_171_in0
	// controller for andOp_171.andOp_171_in1
	// Insensitive connections
	assign andOp_171_in0 = bb_6_active_in_state_2_out_data;
	assign andOp_171_in1 = state_2_is_active;
	// controller for andOp_172.andOp_172_in0
	// controller for andOp_172.andOp_172_in1
	// Insensitive connections
	assign andOp_172_in0 = bb_8_active_in_state_2_out_data;
	assign andOp_172_in1 = state_2_is_active;
	// controller for andOp_173.andOp_173_in0
	// controller for andOp_173.andOp_173_in1
	// Insensitive connections
	assign andOp_173_in0 = bb_8_active_in_state_2_out_data;
	assign andOp_173_in1 = state_2_is_active;
	// controller for andOp_174.andOp_174_in0
	// controller for andOp_174.andOp_174_in1
	// Insensitive connections
	assign andOp_174_in0 = bb_8_active_in_state_2_out_data;
	assign andOp_174_in1 = state_2_is_active;
	// controller for andOp_175.andOp_175_in0
	// controller for andOp_175.andOp_175_in1
	// Insensitive connections
	assign andOp_175_in0 = bb_7_active_in_state_2_out_data;
	assign andOp_175_in1 = state_2_is_active;
	// controller for andOp_176.andOp_176_in0
	// controller for andOp_176.andOp_176_in1
	// Insensitive connections
	assign andOp_176_in0 = bb_7_active_in_state_2_out_data;
	assign andOp_176_in1 = state_2_is_active;
	// controller for andOp_177.andOp_177_in0
	// controller for andOp_177.andOp_177_in1
	// Insensitive connections
	assign andOp_177_in0 = bb_8_active_in_state_3_out_data;
	assign andOp_177_in1 = state_3_is_active;
	// controller for andOp_178.andOp_178_in0
	// controller for andOp_178.andOp_178_in1
	// Insensitive connections
	assign andOp_178_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_178_in1 = state_3_is_active;
	// controller for andOp_179.andOp_179_in0
	// controller for andOp_179.andOp_179_in1
	// Insensitive connections
	assign andOp_179_in0 = bb_2_active_in_state_5_out_data;
	assign andOp_179_in1 = state_5_is_active;
	// controller for andOp_180.andOp_180_in0
	// controller for andOp_180.andOp_180_in1
	// Insensitive connections
	assign andOp_180_in0 = bb_6_active_in_state_1_out_data;
	assign andOp_180_in1 = state_1_is_active;
	// controller for andOp_181.andOp_181_in0
	// controller for andOp_181.andOp_181_in1
	// Insensitive connections
	assign andOp_181_in0 = bb_8_active_in_state_2_out_data;
	assign andOp_181_in1 = state_2_is_active;
	// controller for andOp_182.andOp_182_in0
	// controller for andOp_182.andOp_182_in1
	// Insensitive connections
	assign andOp_182_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_182_in1 = state_3_is_active;
	// controller for andOp_183.andOp_183_in0
	// controller for andOp_183.andOp_183_in1
	// Insensitive connections
	assign andOp_183_in0 = bb_2_active_in_state_4_out_data;
	assign andOp_183_in1 = state_4_is_active;
	// controller for andOp_184.andOp_184_in0
	// controller for andOp_184.andOp_184_in1
	// Insensitive connections
	assign andOp_184_in0 = bb_2_active_in_state_5_out_data;
	assign andOp_184_in1 = state_5_is_active;
	// controller for andOp_186.andOp_186_in0
	// controller for andOp_186.andOp_186_in1
	// Insensitive connections
	assign andOp_186_in0 = notOp_185_out;
	assign andOp_186_in1 = 1'd1;
	// controller for andOp_188.andOp_188_in0
	// controller for andOp_188.andOp_188_in1
	// Insensitive connections
	assign andOp_188_in0 = notOp_187_out;
	assign andOp_188_in1 = andOp_186_out;
	// controller for andOp_190.andOp_190_in0
	// controller for andOp_190.andOp_190_in1
	// Insensitive connections
	assign andOp_190_in0 = notOp_189_out;
	assign andOp_190_in1 = andOp_188_out;
	// controller for andOp_192.andOp_192_in0
	// controller for andOp_192.andOp_192_in1
	// Insensitive connections
	assign andOp_192_in0 = notOp_191_out;
	assign andOp_192_in1 = 1'd1;
	// controller for andOp_194.andOp_194_in0
	// controller for andOp_194.andOp_194_in1
	// Insensitive connections
	assign andOp_194_in0 = notOp_193_out;
	assign andOp_194_in1 = 1'd1;
	// controller for andOp_196.andOp_196_in0
	// controller for andOp_196.andOp_196_in1
	// Insensitive connections
	assign andOp_196_in0 = notOp_195_out;
	assign andOp_196_in1 = andOp_194_out;
	// controller for andOp_198.andOp_198_in0
	// controller for andOp_198.andOp_198_in1
	// Insensitive connections
	assign andOp_198_in0 = notOp_197_out;
	assign andOp_198_in1 = 1'd1;
	// controller for andOp_200.andOp_200_in0
	// controller for andOp_200.andOp_200_in1
	// Insensitive connections
	assign andOp_200_in0 = notOp_199_out;
	assign andOp_200_in1 = 1'd1;
	// controller for andOp_202.andOp_202_in0
	// controller for andOp_202.andOp_202_in1
	// Insensitive connections
	assign andOp_202_in0 = notOp_201_out;
	assign andOp_202_in1 = 1'd1;
	// controller for andOp_204.andOp_204_in0
	// controller for andOp_204.andOp_204_in1
	// Insensitive connections
	assign andOp_204_in0 = notOp_203_out;
	assign andOp_204_in1 = andOp_202_out;
	// controller for andOp_207.andOp_207_in0
	// controller for andOp_207.andOp_207_in1
	// Insensitive connections
	assign andOp_207_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_207_in1 = state_0_is_active;
	// controller for andOp_208.andOp_208_in0
	// controller for andOp_208.andOp_208_in1
	// Insensitive connections
	assign andOp_208_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_208_in1 = state_0_is_active;
	// controller for andOp_209.andOp_209_in0
	// controller for andOp_209.andOp_209_in1
	// Insensitive connections
	assign andOp_209_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_209_in1 = state_0_is_active;
	// controller for andOp_214.andOp_214_in0
	// controller for andOp_214.andOp_214_in1
	// Insensitive connections
	assign andOp_214_in0 = bb_8_active_in_state_2_out_data;
	assign andOp_214_in1 = state_2_is_active;
	// controller for andOp_215.andOp_215_in0
	// controller for andOp_215.andOp_215_in1
	// Insensitive connections
	assign andOp_215_in0 = bb_6_active_in_state_2_out_data;
	assign andOp_215_in1 = state_2_is_active;
	// controller for andOp_40.andOp_40_in0
	// controller for andOp_40.andOp_40_in1
	// Insensitive connections
	assign andOp_40_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_40_in1 = state_0_is_active;
	// controller for andOp_41.andOp_41_in0
	// controller for andOp_41.andOp_41_in1
	// Insensitive connections
	assign andOp_41_in0 = andOp_40_out;
	assign andOp_41_in1 = 1'd1;
	// controller for andOp_43.andOp_43_in0
	// controller for andOp_43.andOp_43_in1
	// Insensitive connections
	assign andOp_43_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_43_in1 = state_0_is_active;
	// controller for andOp_44.andOp_44_in0
	// controller for andOp_44.andOp_44_in1
	// Insensitive connections
	assign andOp_44_in0 = andOp_43_out;
	assign andOp_44_in1 = 1'd1;
	// controller for andOp_46.andOp_46_in0
	// controller for andOp_46.andOp_46_in1
	// Insensitive connections
	assign andOp_46_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_46_in1 = state_0_is_active;
	// controller for andOp_47.andOp_47_in0
	// controller for andOp_47.andOp_47_in1
	// Insensitive connections
	assign andOp_47_in0 = andOp_46_out;
	assign andOp_47_in1 = 1'd1;
	// controller for andOp_49.andOp_49_in0
	// controller for andOp_49.andOp_49_in1
	// Insensitive connections
	assign andOp_49_in0 = andOp_47_out;
	assign andOp_49_in1 = cmp_out_icmp_13;
	// controller for andOp_51.andOp_51_in0
	// controller for andOp_51.andOp_51_in1
	// Insensitive connections
	assign andOp_51_in0 = andOp_47_out;
	assign andOp_51_in1 = notOp_50_out;
	// controller for andOp_52.andOp_52_in0
	// controller for andOp_52.andOp_52_in1
	// Insensitive connections
	assign andOp_52_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_52_in1 = state_0_is_active;
	// controller for andOp_53.andOp_53_in0
	// controller for andOp_53.andOp_53_in1
	// Insensitive connections
	assign andOp_53_in0 = andOp_52_out;
	assign andOp_53_in1 = 1'd1;
	// controller for andOp_55.andOp_55_in0
	// controller for andOp_55.andOp_55_in1
	// Insensitive connections
	assign andOp_55_in0 = bb_5_active_in_state_0_out_data;
	assign andOp_55_in1 = state_0_is_active;
	// controller for andOp_56.andOp_56_in0
	// controller for andOp_56.andOp_56_in1
	// Insensitive connections
	assign andOp_56_in0 = andOp_55_out;
	assign andOp_56_in1 = 1'd1;
	// controller for andOp_58.andOp_58_in0
	// controller for andOp_58.andOp_58_in1
	// Insensitive connections
	assign andOp_58_in0 = andOp_56_out;
	assign andOp_58_in1 = cmp_out_icmp_15;
	// controller for andOp_60.andOp_60_in0
	// controller for andOp_60.andOp_60_in1
	// Insensitive connections
	assign andOp_60_in0 = andOp_56_out;
	assign andOp_60_in1 = notOp_59_out;
	// controller for andOp_61.andOp_61_in0
	// controller for andOp_61.andOp_61_in1
	// Insensitive connections
	assign andOp_61_in0 = bb_6_active_in_state_2_out_data;
	assign andOp_61_in1 = state_2_is_active;
	// controller for andOp_62.andOp_62_in0
	// controller for andOp_62.andOp_62_in1
	// Insensitive connections
	assign andOp_62_in0 = andOp_61_out;
	assign andOp_62_in1 = 1'd1;
	// controller for andOp_64.andOp_64_in0
	// controller for andOp_64.andOp_64_in1
	// Insensitive connections
	assign andOp_64_in0 = bb_6_active_in_state_2_out_data;
	assign andOp_64_in1 = state_2_is_active;
	// controller for andOp_65.andOp_65_in0
	// controller for andOp_65.andOp_65_in1
	// Insensitive connections
	assign andOp_65_in0 = andOp_64_out;
	assign andOp_65_in1 = 1'd1;
	// controller for andOp_67.andOp_67_in0
	// controller for andOp_67.andOp_67_in1
	// Insensitive connections
	assign andOp_67_in0 = bb_7_active_in_state_2_out_data;
	assign andOp_67_in1 = state_2_is_active;
	// controller for andOp_68.andOp_68_in0
	// controller for andOp_68.andOp_68_in1
	// Insensitive connections
	assign andOp_68_in0 = andOp_67_out;
	assign andOp_68_in1 = 1'd1;
	// controller for andOp_70.andOp_70_in0
	// controller for andOp_70.andOp_70_in1
	// Insensitive connections
	assign andOp_70_in0 = andOp_68_out;
	assign andOp_70_in1 = cmp_out_icmp_31;
	// controller for andOp_72.andOp_72_in0
	// controller for andOp_72.andOp_72_in1
	// Insensitive connections
	assign andOp_72_in0 = andOp_68_out;
	assign andOp_72_in1 = notOp_71_out;
	// controller for andOp_73.andOp_73_in0
	// controller for andOp_73.andOp_73_in1
	// Insensitive connections
	assign andOp_73_in0 = bb_8_active_in_state_3_out_data;
	assign andOp_73_in1 = state_3_is_active;
	// controller for andOp_74.andOp_74_in0
	// controller for andOp_74.andOp_74_in1
	// Insensitive connections
	assign andOp_74_in0 = andOp_73_out;
	assign andOp_74_in1 = 1'd1;
	// controller for andOp_76.andOp_76_in0
	// controller for andOp_76.andOp_76_in1
	// Insensitive connections
	assign andOp_76_in0 = andOp_74_out;
	assign andOp_76_in1 = cmp_out_icmp_33;
	// controller for andOp_78.andOp_78_in0
	// controller for andOp_78.andOp_78_in1
	// Insensitive connections
	assign andOp_78_in0 = andOp_74_out;
	assign andOp_78_in1 = notOp_77_out;
	// controller for andOp_79.andOp_79_in0
	// controller for andOp_79.andOp_79_in1
	// Insensitive connections
	assign andOp_79_in0 = bb_8_active_in_state_3_out_data;
	assign andOp_79_in1 = state_3_is_active;
	// controller for andOp_80.andOp_80_in0
	// controller for andOp_80.andOp_80_in1
	// Insensitive connections
	assign andOp_80_in0 = andOp_79_out;
	assign andOp_80_in1 = 1'd1;
	// controller for andOp_82.andOp_82_in0
	// controller for andOp_82.andOp_82_in1
	// Insensitive connections
	assign andOp_82_in0 = andOp_80_out;
	assign andOp_82_in1 = cmp_out_icmp_33;
	// controller for andOp_84.andOp_84_in0
	// controller for andOp_84.andOp_84_in1
	// Insensitive connections
	assign andOp_84_in0 = andOp_80_out;
	assign andOp_84_in1 = notOp_83_out;
	// controller for arg_0.arg_0_read_valid_reg
	always @(*) begin
		if (andOp_170_out) begin 
			arg_0_read_valid_reg = 32'd1;
		end else begin
			arg_0_read_valid_reg = 0;
		end
	end
	// controller for arg_1.arg_1_raddr_reg
	always @(*) begin
		if (andOp_132_out) begin 
			arg_1_raddr_reg = arg_1_rdata;
		end else begin
			arg_1_raddr_reg = 0;
		end
	end
	// controller for arg_2.arg_2_raddr_reg
	always @(*) begin
		if (andOp_133_out) begin 
			arg_2_raddr_reg = arg_2_rdata;
		end else begin
			arg_2_raddr_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_awaddr_reg
	always @(*) begin
		if (andOp_141_out) begin 
			arg_3_s_axi_awaddr_reg = tmp_output_142_out_data;
		end else begin
			arg_3_s_axi_awaddr_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_awburst_reg
	always @(*) begin
		if (andOp_147_out) begin 
			arg_3_s_axi_awburst_reg = 2'd1;
		end else begin
			arg_3_s_axi_awburst_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_awlen_reg
	always @(*) begin
		if (andOp_135_out) begin 
			arg_3_s_axi_awlen_reg = tmp_output_136_out_data;
		end else begin
			arg_3_s_axi_awlen_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_awsize_reg
	always @(*) begin
		if (andOp_149_out) begin 
			arg_3_s_axi_awsize_reg = -(3'd3);
		end else begin
			arg_3_s_axi_awsize_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_awvalid_reg
	always @(*) begin
		if (andOp_150_out) begin 
			arg_3_s_axi_awvalid_reg = 32'd1;
		end else begin
			arg_3_s_axi_awvalid_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_wdata_reg
	always @(*) begin
		if (andOp_153_out) begin 
			arg_3_s_axi_wdata_reg = tmp_output_154_out_data;
		end else if (andOp_160_out) begin 
			arg_3_s_axi_wdata_reg = 32'd0;
		end else begin
			arg_3_s_axi_wdata_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_wstrb_reg
	always @(*) begin
		if (andOp_157_out) begin 
			arg_3_s_axi_wstrb_reg = -(4'd1);
		end else if (andOp_161_out) begin 
			arg_3_s_axi_wstrb_reg = 32'd0;
		end else begin
			arg_3_s_axi_wstrb_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_wvalid_reg
	always @(*) begin
		if (andOp_148_out) begin 
			arg_3_s_axi_wvalid_reg = 32'd1;
		end else if (andOp_152_out) begin 
			arg_3_s_axi_wvalid_reg = 32'd1;
		end else if (andOp_159_out) begin 
			arg_3_s_axi_wvalid_reg = 32'd1;
		end else begin
			arg_3_s_axi_wvalid_reg = 0;
		end
	end
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_85_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_105_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_0.bb_1_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_0_in_data = orOp_87_out;
		end else begin
			bb_1_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_0.bb_1_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_108_out) begin 
			bb_1_predecessor_in_state_0_in_data = 32'd4;
		end else if (eq_106_out) begin 
			bb_1_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_3.bb_2_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_3_in_data = orOp_101_out;
		end else begin
			bb_2_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_4.bb_2_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_4_in_data = eq_103_out;
		end else begin
			bb_2_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_5.bb_2_active_in_state_5_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_5_in_data = eq_104_out;
		end else begin
			bb_2_active_in_state_5_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_3.bb_2_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_128_out) begin 
			bb_2_predecessor_in_state_3_in_data = 32'd8;
		end else if (eq_126_out) begin 
			bb_2_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_4.bb_2_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_130_out) begin 
			bb_2_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_5.bb_2_predecessor_in_state_5_in_data
	always @(*) begin
		if (eq_131_out) begin 
			bb_2_predecessor_in_state_5_in_data = state_5_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_5_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_0.bb_3_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_0_in_data = orOp_89_out;
		end else begin
			bb_3_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_0.bb_3_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_111_out) begin 
			bb_3_predecessor_in_state_0_in_data = 32'd0;
		end else if (eq_109_out) begin 
			bb_3_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_0.bb_4_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_0_in_data = orOp_91_out;
		end else begin
			bb_4_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_0.bb_4_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_114_out) begin 
			bb_4_predecessor_in_state_0_in_data = 32'd3;
		end else if (eq_112_out) begin 
			bb_4_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_5_active_in_state_0.bb_5_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_5_active_in_state_0_in_data = orOp_93_out;
		end else begin
			bb_5_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_5_predecessor_in_state_0.bb_5_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_117_out) begin 
			bb_5_predecessor_in_state_0_in_data = 32'd1;
		end else if (eq_115_out) begin 
			bb_5_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_5_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_6_active_in_state_1.bb_6_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_6_active_in_state_1_in_data = eq_94_out;
		end else begin
			bb_6_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_6_active_in_state_2.bb_6_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_6_active_in_state_2_in_data = eq_95_out;
		end else begin
			bb_6_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_6_predecessor_in_state_1.bb_6_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_118_out) begin 
			bb_6_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_6_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_6_predecessor_in_state_2.bb_6_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_119_out) begin 
			bb_6_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_6_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_7_active_in_state_2.bb_7_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_7_active_in_state_2_in_data = orOp_97_out;
		end else begin
			bb_7_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_7_predecessor_in_state_2.bb_7_predecessor_in_state_2_in_data
	always @(*) begin
		if (andOp_122_out) begin 
			bb_7_predecessor_in_state_2_in_data = 32'd6;
		end else if (eq_120_out) begin 
			bb_7_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_7_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_8_active_in_state_2.bb_8_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_state_2_in_data = orOp_99_out;
		end else begin
			bb_8_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_8_active_in_state_3.bb_8_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_state_3_in_data = eq_102_out;
		end else begin
			bb_8_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_8_predecessor_in_state_2.bb_8_predecessor_in_state_2_in_data
	always @(*) begin
		if (andOp_125_out) begin 
			bb_8_predecessor_in_state_2_in_data = 32'd7;
		end else if (eq_123_out) begin 
			bb_8_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_8_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_8_predecessor_in_state_3.bb_8_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_129_out) begin 
			bb_8_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_8_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_41_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_42_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_1_happened_in_state_0.br_1_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_44_out) begin 
			br_1_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_45_out) begin 
			br_1_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_1_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_0.br_3_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_47_out) begin 
			br_3_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_48_out) begin 
			br_3_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_0.br_4_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_53_out) begin 
			br_4_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_54_out) begin 
			br_4_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_5_happened_in_state_0.br_5_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_56_out) begin 
			br_5_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_57_out) begin 
			br_5_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_5_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_6_happened_in_state_1.br_6_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_62_out) begin 
			br_6_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_63_out) begin 
			br_6_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_6_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_6_happened_in_state_2.br_6_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_65_out) begin 
			br_6_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_66_out) begin 
			br_6_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_6_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_7_happened_in_state_2.br_7_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_68_out) begin 
			br_7_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_69_out) begin 
			br_7_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_7_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_8_happened_in_state_2.br_8_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_74_out) begin 
			br_8_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_75_out) begin 
			br_8_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_8_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_8_happened_in_state_3.br_8_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_80_out) begin 
			br_8_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_81_out) begin 
			br_8_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_8_happened_in_state_3_in_data = 0;
		end
	end
	// controller for concat_163.concat_163_in0
	// controller for concat_163.concat_163_in1
	// Insensitive connections
	assign concat_163_in0 = 8'd0;
	assign concat_163_in1 = data_in_0_5_out_data;
	// controller for concat_164.concat_164_in0
	// controller for concat_164.concat_164_in1
	// Insensitive connections
	assign concat_164_in0 = 32'd4;
	assign concat_164_in1 = 32'd8;
	// controller for data_in_0_1.data_in_0_1_in_data
	always @(*) begin
		if (eq_205_out) begin 
			data_in_0_1_in_data = data_store_0_0;
		end else if (eq_206_out) begin 
			data_in_0_1_in_data = data_store_3_30;
		end else begin
			data_in_0_1_in_data = 0;
		end
	end
	// controller for data_in_0_3.data_in_0_3_in_data
	always @(*) begin
		if (eq_205_out) begin 
			data_in_0_3_in_data = data_store_0_2;
		end else if (eq_206_out) begin 
			data_in_0_3_in_data = data_store_3_32;
		end else begin
			data_in_0_3_in_data = 0;
		end
	end
	// controller for data_in_0_5.data_in_0_5_in_data
	always @(*) begin
		if (eq_205_out) begin 
			data_in_0_5_in_data = data_store_0_4;
		end else if (eq_206_out) begin 
			data_in_0_5_in_data = data_store_3_34;
		end else begin
			data_in_0_5_in_data = 0;
		end
	end
	// controller for data_in_0_7.data_in_0_7_in_data
	always @(*) begin
		if (eq_205_out) begin 
			data_in_0_7_in_data = data_store_0_6;
		end else if (eq_206_out) begin 
			data_in_0_7_in_data = data_store_3_36;
		end else begin
			data_in_0_7_in_data = 0;
		end
	end
	// controller for data_in_0_9.data_in_0_9_in_data
	always @(*) begin
		if (eq_205_out) begin 
			data_in_0_9_in_data = data_store_0_8;
		end else if (eq_206_out) begin 
			data_in_0_9_in_data = data_store_3_38;
		end else begin
			data_in_0_9_in_data = 0;
		end
	end
	// controller for data_in_1_11.data_in_1_11_in_data
	always @(*) begin
		if (eq_210_out) begin 
			data_in_1_11_in_data = data_store_0_0;
		end else if (eq_211_out) begin 
			data_in_1_11_in_data = data_store_1_10;
		end else begin
			data_in_1_11_in_data = 0;
		end
	end
	// controller for data_in_1_13.data_in_1_13_in_data
	always @(*) begin
		if (eq_210_out) begin 
			data_in_1_13_in_data = data_store_0_2;
		end else if (eq_211_out) begin 
			data_in_1_13_in_data = data_store_1_12;
		end else begin
			data_in_1_13_in_data = 0;
		end
	end
	// controller for data_in_1_15.data_in_1_15_in_data
	always @(*) begin
		if (eq_210_out) begin 
			data_in_1_15_in_data = data_store_0_4;
		end else if (eq_211_out) begin 
			data_in_1_15_in_data = data_store_1_14;
		end else begin
			data_in_1_15_in_data = 0;
		end
	end
	// controller for data_in_1_17.data_in_1_17_in_data
	always @(*) begin
		if (eq_210_out) begin 
			data_in_1_17_in_data = data_store_0_6;
		end else if (eq_211_out) begin 
			data_in_1_17_in_data = data_store_1_16;
		end else begin
			data_in_1_17_in_data = 0;
		end
	end
	// controller for data_in_1_19.data_in_1_19_in_data
	always @(*) begin
		if (eq_210_out) begin 
			data_in_1_19_in_data = data_store_0_8;
		end else if (eq_211_out) begin 
			data_in_1_19_in_data = data_store_1_18;
		end else begin
			data_in_1_19_in_data = 0;
		end
	end
	// controller for data_in_2_21.data_in_2_21_in_data
	always @(*) begin
		if (eq_212_out) begin 
			data_in_2_21_in_data = data_store_1_10;
		end else if (eq_213_out) begin 
			data_in_2_21_in_data = data_store_2_20;
		end else begin
			data_in_2_21_in_data = 0;
		end
	end
	// controller for data_in_2_23.data_in_2_23_in_data
	always @(*) begin
		if (eq_212_out) begin 
			data_in_2_23_in_data = data_store_1_12;
		end else if (eq_213_out) begin 
			data_in_2_23_in_data = data_store_2_22;
		end else begin
			data_in_2_23_in_data = 0;
		end
	end
	// controller for data_in_2_25.data_in_2_25_in_data
	always @(*) begin
		if (eq_212_out) begin 
			data_in_2_25_in_data = data_store_1_14;
		end else if (eq_213_out) begin 
			data_in_2_25_in_data = data_store_2_24;
		end else begin
			data_in_2_25_in_data = 0;
		end
	end
	// controller for data_in_2_27.data_in_2_27_in_data
	always @(*) begin
		if (eq_212_out) begin 
			data_in_2_27_in_data = data_store_1_16;
		end else if (eq_213_out) begin 
			data_in_2_27_in_data = data_store_2_26;
		end else begin
			data_in_2_27_in_data = 0;
		end
	end
	// controller for data_in_2_29.data_in_2_29_in_data
	always @(*) begin
		if (eq_212_out) begin 
			data_in_2_29_in_data = data_store_1_18;
		end else if (eq_213_out) begin 
			data_in_2_29_in_data = data_store_2_28;
		end else begin
			data_in_2_29_in_data = 0;
		end
	end
	// controller for data_in_3_31.data_in_3_31_in_data
	always @(*) begin
		if (eq_216_out) begin 
			data_in_3_31_in_data = data_store_2_20;
		end else if (eq_217_out) begin 
			data_in_3_31_in_data = data_store_3_30;
		end else begin
			data_in_3_31_in_data = 0;
		end
	end
	// controller for data_in_3_33.data_in_3_33_in_data
	always @(*) begin
		if (eq_216_out) begin 
			data_in_3_33_in_data = data_store_2_22;
		end else if (eq_217_out) begin 
			data_in_3_33_in_data = data_store_3_32;
		end else begin
			data_in_3_33_in_data = 0;
		end
	end
	// controller for data_in_3_35.data_in_3_35_in_data
	always @(*) begin
		if (eq_216_out) begin 
			data_in_3_35_in_data = data_store_2_24;
		end else if (eq_217_out) begin 
			data_in_3_35_in_data = data_store_3_34;
		end else begin
			data_in_3_35_in_data = 0;
		end
	end
	// controller for data_in_3_37.data_in_3_37_in_data
	always @(*) begin
		if (eq_216_out) begin 
			data_in_3_37_in_data = data_store_2_26;
		end else if (eq_217_out) begin 
			data_in_3_37_in_data = data_store_3_36;
		end else begin
			data_in_3_37_in_data = 0;
		end
	end
	// controller for data_in_3_39.data_in_3_39_in_data
	always @(*) begin
		if (eq_216_out) begin 
			data_in_3_39_in_data = data_store_2_28;
		end else if (eq_217_out) begin 
			data_in_3_39_in_data = data_store_3_38;
		end else begin
			data_in_3_39_in_data = 0;
		end
	end
	// controller for eq_100.eq_100_in0
	// controller for eq_100.eq_100_in1
	// Insensitive connections
	assign eq_100_in0 = 32'd2;
	assign eq_100_in1 = state_3_entry_BB_reg;
	// controller for eq_102.eq_102_in0
	// controller for eq_102.eq_102_in1
	// Insensitive connections
	assign eq_102_in0 = 32'd8;
	assign eq_102_in1 = state_3_entry_BB_reg;
	// controller for eq_103.eq_103_in0
	// controller for eq_103.eq_103_in1
	// Insensitive connections
	assign eq_103_in0 = 32'd2;
	assign eq_103_in1 = state_4_entry_BB_reg;
	// controller for eq_104.eq_104_in0
	// controller for eq_104.eq_104_in1
	// Insensitive connections
	assign eq_104_in0 = 32'd2;
	assign eq_104_in1 = state_5_entry_BB_reg;
	// controller for eq_105.eq_105_in0
	// controller for eq_105.eq_105_in1
	// Insensitive connections
	assign eq_105_in0 = 32'd0;
	assign eq_105_in1 = state_0_entry_BB_reg;
	// controller for eq_106.eq_106_in0
	// controller for eq_106.eq_106_in1
	// Insensitive connections
	assign eq_106_in0 = 32'd1;
	assign eq_106_in1 = state_0_entry_BB_reg;
	// controller for eq_109.eq_109_in0
	// controller for eq_109.eq_109_in1
	// Insensitive connections
	assign eq_109_in0 = 32'd3;
	assign eq_109_in1 = state_0_entry_BB_reg;
	// controller for eq_112.eq_112_in0
	// controller for eq_112.eq_112_in1
	// Insensitive connections
	assign eq_112_in0 = 32'd4;
	assign eq_112_in1 = state_0_entry_BB_reg;
	// controller for eq_115.eq_115_in0
	// controller for eq_115.eq_115_in1
	// Insensitive connections
	assign eq_115_in0 = 32'd5;
	assign eq_115_in1 = state_0_entry_BB_reg;
	// controller for eq_118.eq_118_in0
	// controller for eq_118.eq_118_in1
	// Insensitive connections
	assign eq_118_in0 = 32'd6;
	assign eq_118_in1 = state_1_entry_BB_reg;
	// controller for eq_119.eq_119_in0
	// controller for eq_119.eq_119_in1
	// Insensitive connections
	assign eq_119_in0 = 32'd6;
	assign eq_119_in1 = state_2_entry_BB_reg;
	// controller for eq_120.eq_120_in0
	// controller for eq_120.eq_120_in1
	// Insensitive connections
	assign eq_120_in0 = 32'd7;
	assign eq_120_in1 = state_2_entry_BB_reg;
	// controller for eq_123.eq_123_in0
	// controller for eq_123.eq_123_in1
	// Insensitive connections
	assign eq_123_in0 = 32'd8;
	assign eq_123_in1 = state_2_entry_BB_reg;
	// controller for eq_126.eq_126_in0
	// controller for eq_126.eq_126_in1
	// Insensitive connections
	assign eq_126_in0 = 32'd2;
	assign eq_126_in1 = state_3_entry_BB_reg;
	// controller for eq_129.eq_129_in0
	// controller for eq_129.eq_129_in1
	// Insensitive connections
	assign eq_129_in0 = 32'd8;
	assign eq_129_in1 = state_3_entry_BB_reg;
	// controller for eq_130.eq_130_in0
	// controller for eq_130.eq_130_in1
	// Insensitive connections
	assign eq_130_in0 = 32'd2;
	assign eq_130_in1 = state_4_entry_BB_reg;
	// controller for eq_131.eq_131_in0
	// controller for eq_131.eq_131_in1
	// Insensitive connections
	assign eq_131_in0 = 32'd2;
	assign eq_131_in1 = state_5_entry_BB_reg;
	// controller for eq_137.eq_137_in0
	// controller for eq_137.eq_137_in1
	// Insensitive connections
	assign eq_137_in0 = 32'd0;
	assign eq_137_in1 = state_0_entry_BB_reg;
	// controller for eq_138.eq_138_in0
	// controller for eq_138.eq_138_in1
	// Insensitive connections
	assign eq_138_in0 = 32'd1;
	assign eq_138_in1 = state_0_entry_BB_reg;
	// controller for eq_139.eq_139_in0
	// controller for eq_139.eq_139_in1
	// Insensitive connections
	assign eq_139_in0 = 32'd3;
	assign eq_139_in1 = state_0_entry_BB_reg;
	// controller for eq_140.eq_140_in0
	// controller for eq_140.eq_140_in1
	// Insensitive connections
	assign eq_140_in0 = 32'd5;
	assign eq_140_in1 = state_0_entry_BB_reg;
	// controller for eq_143.eq_143_in0
	// controller for eq_143.eq_143_in1
	// Insensitive connections
	assign eq_143_in0 = 32'd0;
	assign eq_143_in1 = state_0_entry_BB_reg;
	// controller for eq_144.eq_144_in0
	// controller for eq_144.eq_144_in1
	// Insensitive connections
	assign eq_144_in0 = 32'd1;
	assign eq_144_in1 = state_0_entry_BB_reg;
	// controller for eq_145.eq_145_in0
	// controller for eq_145.eq_145_in1
	// Insensitive connections
	assign eq_145_in0 = 32'd3;
	assign eq_145_in1 = state_0_entry_BB_reg;
	// controller for eq_146.eq_146_in0
	// controller for eq_146.eq_146_in1
	// Insensitive connections
	assign eq_146_in0 = 32'd5;
	assign eq_146_in1 = state_0_entry_BB_reg;
	// controller for eq_155.eq_155_in0
	// controller for eq_155.eq_155_in1
	// Insensitive connections
	assign eq_155_in0 = 32'd6;
	assign eq_155_in1 = state_2_entry_BB_reg;
	// controller for eq_156.eq_156_in0
	// controller for eq_156.eq_156_in1
	// Insensitive connections
	assign eq_156_in0 = 32'd7;
	assign eq_156_in1 = state_2_entry_BB_reg;
	// controller for eq_205.eq_205_in0
	// controller for eq_205.eq_205_in1
	// Insensitive connections
	assign eq_205_in0 = 32'd0;
	assign eq_205_in1 = state_0_last_state;
	// controller for eq_206.eq_206_in0
	// controller for eq_206.eq_206_in1
	// Insensitive connections
	assign eq_206_in0 = 32'd3;
	assign eq_206_in1 = state_0_last_state;
	// controller for eq_210.eq_210_in0
	// controller for eq_210.eq_210_in1
	// Insensitive connections
	assign eq_210_in0 = 32'd0;
	assign eq_210_in1 = state_1_last_state;
	// controller for eq_211.eq_211_in0
	// controller for eq_211.eq_211_in1
	// Insensitive connections
	assign eq_211_in0 = 32'd1;
	assign eq_211_in1 = state_1_last_state;
	// controller for eq_212.eq_212_in0
	// controller for eq_212.eq_212_in1
	// Insensitive connections
	assign eq_212_in0 = 32'd1;
	assign eq_212_in1 = state_2_last_state;
	// controller for eq_213.eq_213_in0
	// controller for eq_213.eq_213_in1
	// Insensitive connections
	assign eq_213_in0 = 32'd2;
	assign eq_213_in1 = state_2_last_state;
	// controller for eq_216.eq_216_in0
	// controller for eq_216.eq_216_in1
	// Insensitive connections
	assign eq_216_in0 = 32'd2;
	assign eq_216_in1 = state_3_last_state;
	// controller for eq_217.eq_217_in0
	// controller for eq_217.eq_217_in1
	// Insensitive connections
	assign eq_217_in0 = 32'd3;
	assign eq_217_in1 = state_3_last_state;
	// controller for eq_218.eq_218_in0
	// controller for eq_218.eq_218_in1
	// Insensitive connections
	assign eq_218_in0 = 32'd3;
	assign eq_218_in1 = state_4_last_state;
	// controller for eq_219.eq_219_in0
	// controller for eq_219.eq_219_in1
	// Insensitive connections
	assign eq_219_in0 = 32'd4;
	assign eq_219_in1 = state_4_last_state;
	// controller for eq_220.eq_220_in0
	// controller for eq_220.eq_220_in1
	// Insensitive connections
	assign eq_220_in0 = 32'd4;
	assign eq_220_in1 = state_5_last_state;
	// controller for eq_221.eq_221_in0
	// controller for eq_221.eq_221_in1
	// Insensitive connections
	assign eq_221_in0 = 32'd5;
	assign eq_221_in1 = state_5_last_state;
	// controller for eq_85.eq_85_in0
	// controller for eq_85.eq_85_in1
	// Insensitive connections
	assign eq_85_in0 = 32'd0;
	assign eq_85_in1 = state_0_entry_BB_reg;
	// controller for eq_86.eq_86_in0
	// controller for eq_86.eq_86_in1
	// Insensitive connections
	assign eq_86_in0 = 32'd1;
	assign eq_86_in1 = state_0_entry_BB_reg;
	// controller for eq_88.eq_88_in0
	// controller for eq_88.eq_88_in1
	// Insensitive connections
	assign eq_88_in0 = 32'd3;
	assign eq_88_in1 = state_0_entry_BB_reg;
	// controller for eq_90.eq_90_in0
	// controller for eq_90.eq_90_in1
	// Insensitive connections
	assign eq_90_in0 = 32'd4;
	assign eq_90_in1 = state_0_entry_BB_reg;
	// controller for eq_92.eq_92_in0
	// controller for eq_92.eq_92_in1
	// Insensitive connections
	assign eq_92_in0 = 32'd5;
	assign eq_92_in1 = state_0_entry_BB_reg;
	// controller for eq_94.eq_94_in0
	// controller for eq_94.eq_94_in1
	// Insensitive connections
	assign eq_94_in0 = 32'd6;
	assign eq_94_in1 = state_1_entry_BB_reg;
	// controller for eq_95.eq_95_in0
	// controller for eq_95.eq_95_in1
	// Insensitive connections
	assign eq_95_in0 = 32'd6;
	assign eq_95_in1 = state_2_entry_BB_reg;
	// controller for eq_96.eq_96_in0
	// controller for eq_96.eq_96_in1
	// Insensitive connections
	assign eq_96_in0 = 32'd7;
	assign eq_96_in1 = state_2_entry_BB_reg;
	// controller for eq_98.eq_98_in0
	// controller for eq_98.eq_98_in1
	// Insensitive connections
	assign eq_98_in0 = 32'd8;
	assign eq_98_in1 = state_2_entry_BB_reg;
	// controller for icmp_13.cmp_in0_icmp_13
	// controller for icmp_13.cmp_in1_icmp_13
	// Insensitive connections
	assign cmp_in0_icmp_13 = sgt_out_sext_12;
	assign cmp_in1_icmp_13 = 32'd0;
	// controller for icmp_15.cmp_in0_icmp_15
	// controller for icmp_15.cmp_in1_icmp_15
	// Insensitive connections
	assign cmp_in0_icmp_15 = sgt_out_sext_8;
	assign cmp_in1_icmp_15 = 32'd0;
	// controller for icmp_31.cmp_in0_icmp_31
	// controller for icmp_31.cmp_in1_icmp_31
	// Insensitive connections
	assign cmp_in0_icmp_31 = sgt_out_sext_30;
	assign cmp_in1_icmp_31 = 32'd0;
	// controller for icmp_33.cmp_in0_icmp_33
	// controller for icmp_33.cmp_in1_icmp_33
	// Insensitive connections
	assign cmp_in0_icmp_33 = data_in_3_35_out_data;
	assign cmp_in1_icmp_33 = data_in_3_31_out_data;
	// controller for notOp_107.notOp_107_in0
	// Insensitive connections
	assign notOp_107_in0 = eq_106_out;
	// controller for notOp_110.notOp_110_in0
	// Insensitive connections
	assign notOp_110_in0 = eq_109_out;
	// controller for notOp_113.notOp_113_in0
	// Insensitive connections
	assign notOp_113_in0 = eq_112_out;
	// controller for notOp_116.notOp_116_in0
	// Insensitive connections
	assign notOp_116_in0 = eq_115_out;
	// controller for notOp_121.notOp_121_in0
	// Insensitive connections
	assign notOp_121_in0 = eq_120_out;
	// controller for notOp_124.notOp_124_in0
	// Insensitive connections
	assign notOp_124_in0 = eq_123_out;
	// controller for notOp_127.notOp_127_in0
	// Insensitive connections
	assign notOp_127_in0 = eq_126_out;
	// controller for notOp_185.notOp_185_in0
	// Insensitive connections
	assign notOp_185_in0 = andOp_49_out;
	// controller for notOp_187.notOp_187_in0
	// Insensitive connections
	assign notOp_187_in0 = andOp_58_out;
	// controller for notOp_189.notOp_189_in0
	// Insensitive connections
	assign notOp_189_in0 = andOp_76_out;
	// controller for notOp_191.notOp_191_in0
	// Insensitive connections
	assign notOp_191_in0 = andOp_60_out;
	// controller for notOp_193.notOp_193_in0
	// Insensitive connections
	assign notOp_193_in0 = andOp_180_out;
	// controller for notOp_195.notOp_195_in0
	// Insensitive connections
	assign notOp_195_in0 = andOp_70_out;
	// controller for notOp_197.notOp_197_in0
	// Insensitive connections
	assign notOp_197_in0 = andOp_181_out;
	// controller for notOp_199.notOp_199_in0
	// Insensitive connections
	assign notOp_199_in0 = andOp_182_out;
	// controller for notOp_201.notOp_201_in0
	// Insensitive connections
	assign notOp_201_in0 = andOp_183_out;
	// controller for notOp_203.notOp_203_in0
	// Insensitive connections
	assign notOp_203_in0 = andOp_184_out;
	// controller for notOp_42.notOp_42_in0
	// Insensitive connections
	assign notOp_42_in0 = andOp_41_out;
	// controller for notOp_45.notOp_45_in0
	// Insensitive connections
	assign notOp_45_in0 = andOp_44_out;
	// controller for notOp_48.notOp_48_in0
	// Insensitive connections
	assign notOp_48_in0 = andOp_47_out;
	// controller for notOp_50.notOp_50_in0
	// Insensitive connections
	assign notOp_50_in0 = cmp_out_icmp_13;
	// controller for notOp_54.notOp_54_in0
	// Insensitive connections
	assign notOp_54_in0 = andOp_53_out;
	// controller for notOp_57.notOp_57_in0
	// Insensitive connections
	assign notOp_57_in0 = andOp_56_out;
	// controller for notOp_59.notOp_59_in0
	// Insensitive connections
	assign notOp_59_in0 = cmp_out_icmp_15;
	// controller for notOp_63.notOp_63_in0
	// Insensitive connections
	assign notOp_63_in0 = andOp_62_out;
	// controller for notOp_66.notOp_66_in0
	// Insensitive connections
	assign notOp_66_in0 = andOp_65_out;
	// controller for notOp_69.notOp_69_in0
	// Insensitive connections
	assign notOp_69_in0 = andOp_68_out;
	// controller for notOp_71.notOp_71_in0
	// Insensitive connections
	assign notOp_71_in0 = cmp_out_icmp_31;
	// controller for notOp_75.notOp_75_in0
	// Insensitive connections
	assign notOp_75_in0 = andOp_74_out;
	// controller for notOp_77.notOp_77_in0
	// Insensitive connections
	assign notOp_77_in0 = cmp_out_icmp_33;
	// controller for notOp_81.notOp_81_in0
	// Insensitive connections
	assign notOp_81_in0 = andOp_80_out;
	// controller for notOp_83.notOp_83_in0
	// Insensitive connections
	assign notOp_83_in0 = cmp_out_icmp_33;
	// controller for orOp_101.orOp_101_in0
	// controller for orOp_101.orOp_101_in1
	// Insensitive connections
	assign orOp_101_in0 = eq_100_out;
	assign orOp_101_in1 = andOp_78_out;
	// controller for orOp_87.orOp_87_in0
	// controller for orOp_87.orOp_87_in1
	// Insensitive connections
	assign orOp_87_in0 = eq_86_out;
	assign orOp_87_in1 = andOp_53_out;
	// controller for orOp_89.orOp_89_in0
	// controller for orOp_89.orOp_89_in1
	// Insensitive connections
	assign orOp_89_in0 = eq_88_out;
	assign orOp_89_in1 = andOp_41_out;
	// controller for orOp_91.orOp_91_in0
	// controller for orOp_91.orOp_91_in1
	// Insensitive connections
	assign orOp_91_in0 = eq_90_out;
	assign orOp_91_in1 = andOp_51_out;
	// controller for orOp_93.orOp_93_in0
	// controller for orOp_93.orOp_93_in1
	// Insensitive connections
	assign orOp_93_in0 = eq_92_out;
	assign orOp_93_in1 = andOp_44_out;
	// controller for orOp_97.orOp_97_in0
	// controller for orOp_97.orOp_97_in1
	// Insensitive connections
	assign orOp_97_in0 = eq_96_out;
	assign orOp_97_in1 = andOp_62_out;
	// controller for orOp_99.orOp_99_in0
	// controller for orOp_99.orOp_99_in1
	// Insensitive connections
	assign orOp_99_in0 = eq_98_out;
	assign orOp_99_in1 = andOp_72_out;
	// controller for phi_5.phi_in_phi_5
	// controller for phi_5.phi_last_block_phi_5
	// controller for phi_5.phi_s_phi_5
	// Insensitive connections
	assign phi_in_phi_5 = concat_163_out;
	assign phi_last_block_phi_5 = bb_1_predecessor_in_state_0_out_data;
	assign phi_s_phi_5 = concat_164_out;
	// controller for ret_40.valid_reg
	always @(*) begin
		if (andOp_179_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// controller for sext_12.sgt_in0_sext_12
	// Insensitive connections
	assign sgt_in0_sext_12 = arg_3_s_axi_awready;
	// controller for sext_21.sgt_in0_sext_21
	// Insensitive connections
	assign sgt_in0_sext_21 = data_in_2_27_out_data;
	// controller for sext_30.sgt_in0_sext_30
	// Insensitive connections
	assign sgt_in0_sext_30 = arg_3_s_axi_wready;
	// controller for sext_8.sgt_in0_sext_8
	// Insensitive connections
	assign sgt_in0_sext_8 = arg_0_read_ready;
	// controller for tmp_output_136.tmp_output_136_in_data
	always @(*) begin
		if (eq_137_out) begin 
			tmp_output_136_in_data = arg_1_rdata;
		end else if (eq_139_out) begin 
			tmp_output_136_in_data = data_in_0_1_out_data;
		end else begin
			tmp_output_136_in_data = 0;
		end
	end
	// controller for tmp_output_142.tmp_output_142_in_data
	always @(*) begin
		if (eq_143_out) begin 
			tmp_output_142_in_data = arg_2_rdata;
		end else if (eq_145_out) begin 
			tmp_output_142_in_data = data_in_0_3_out_data;
		end else begin
			tmp_output_142_in_data = 0;
		end
	end
	// controller for tmp_output_154.tmp_output_154_in_data
	always @(*) begin
		if (eq_155_out) begin 
			tmp_output_154_in_data = arg_0_out_data;
		end else if (eq_156_out) begin 
			tmp_output_154_in_data = data_in_2_29_out_data;
		end else begin
			tmp_output_154_in_data = 0;
		end
	end
	// controller for trunc_23.trunc_in_trunc_23
	// Insensitive connections
	assign trunc_in_trunc_23 = add_out_add_22;
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			data_store_0_0 <= 0;
		end else begin
			if (andOp_207_out) begin
				data_store_0_0 <= arg_1_rdata;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_2 <= 0;
		end else begin
			if (andOp_208_out) begin
				data_store_0_2 <= arg_2_rdata;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_4 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_4 <= data_in_0_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_6 <= 0;
		end else begin
			if (andOp_209_out) begin
				data_store_0_6 <= phi_out_phi_5;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_8 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_8 <= data_in_0_9_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_10 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_10 <= data_in_1_11_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_12 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_12 <= data_in_1_13_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_14 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_14 <= data_in_1_15_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_16 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_16 <= data_in_1_17_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_18 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_18 <= data_in_1_19_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_20 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_20 <= data_in_2_21_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_22 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_22 <= data_in_2_23_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_24 <= 0;
		end else begin
			if (andOp_214_out) begin
				data_store_2_24 <= trunc_out_trunc_23;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_26 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_26 <= data_in_2_27_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_28 <= 0;
		end else begin
			if (andOp_215_out) begin
				data_store_2_28 <= arg_0_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_30 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_30 <= data_in_3_31_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_32 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_32 <= data_in_3_33_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_34 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_34 <= data_in_3_35_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_36 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_36 <= data_in_3_37_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_38 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_38 <= data_in_3_39_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_180_out) begin
				global_state <= 32'd2;
			end
			if (andOp_181_out) begin
				global_state <= 32'd3;
			end
			if (andOp_182_out) begin
				global_state <= 32'd4;
			end
			if (andOp_183_out) begin
				global_state <= 32'd5;
			end
			if (andOp_184_out) begin
				global_state <= 32'd5;
			end
			if (andOp_49_out) begin
				global_state <= 32'd0;
			end
			if (andOp_58_out) begin
				global_state <= 32'd0;
			end
			if (andOp_60_out) begin
				global_state <= 32'd1;
			end
			if (andOp_70_out) begin
				global_state <= 32'd2;
			end
			if (andOp_76_out) begin
				global_state <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
			if (andOp_49_out) begin
				state_0_entry_BB_reg <= 32'd3;
			end
			if (andOp_58_out) begin
				state_0_entry_BB_reg <= 32'd5;
			end
			if (andOp_76_out) begin
				state_0_entry_BB_reg <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (andOp_190_out) begin
				state_0_is_active <= 1'd0;
			end
			if (andOp_49_out) begin
				state_0_is_active <= 1'd1;
			end
			if (andOp_58_out) begin
				state_0_is_active <= 1'd1;
			end
			if (andOp_76_out) begin
				state_0_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
			if (andOp_49_out) begin
				state_0_last_BB_reg <= 32'd3;
			end
			if (andOp_58_out) begin
				state_0_last_BB_reg <= 32'd5;
			end
			if (andOp_76_out) begin
				state_0_last_BB_reg <= 32'd8;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
			if (andOp_49_out) begin
				state_0_last_state <= 32'd0;
			end
			if (andOp_58_out) begin
				state_0_last_state <= 32'd0;
			end
			if (andOp_76_out) begin
				state_0_last_state <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_60_out) begin
				state_1_entry_BB_reg <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_192_out) begin
				state_1_is_active <= 1'd0;
			end
			if (andOp_60_out) begin
				state_1_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_60_out) begin
				state_1_last_BB_reg <= 32'd5;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_60_out) begin
				state_1_last_state <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_180_out) begin
				state_2_entry_BB_reg <= 32'd6;
			end
			if (andOp_70_out) begin
				state_2_entry_BB_reg <= 32'd7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_180_out) begin
				state_2_is_active <= 1'd1;
			end
			if (andOp_196_out) begin
				state_2_is_active <= 1'd0;
			end
			if (andOp_70_out) begin
				state_2_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_180_out) begin
				state_2_last_BB_reg <= bb_6_predecessor_in_state_1_out_data;
			end
			if (andOp_70_out) begin
				state_2_last_BB_reg <= 32'd7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_180_out) begin
				state_2_last_state <= 32'd1;
			end
			if (andOp_70_out) begin
				state_2_last_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_181_out) begin
				state_3_entry_BB_reg <= 32'd8;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_181_out) begin
				state_3_is_active <= 1'd1;
			end
			if (andOp_198_out) begin
				state_3_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_181_out) begin
				state_3_last_BB_reg <= bb_8_predecessor_in_state_2_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_state <= 0;
		end else begin
			if (andOp_181_out) begin
				state_3_last_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_182_out) begin
				state_4_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_182_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_200_out) begin
				state_4_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_182_out) begin
				state_4_last_BB_reg <= bb_2_predecessor_in_state_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_state <= 0;
		end else begin
			if (andOp_182_out) begin
				state_4_last_state <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_entry_BB_reg <= 0;
		end else begin
			if (andOp_183_out) begin
				state_5_entry_BB_reg <= 32'd2;
			end
			if (andOp_184_out) begin
				state_5_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_is_active <= 0;
		end else begin
			if (andOp_183_out) begin
				state_5_is_active <= 1'd1;
			end
			if (andOp_184_out) begin
				state_5_is_active <= 1'd1;
			end
			if (andOp_204_out) begin
				state_5_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_last_BB_reg <= 0;
		end else begin
			if (andOp_183_out) begin
				state_5_last_BB_reg <= bb_2_predecessor_in_state_4_out_data;
			end
			if (andOp_184_out) begin
				state_5_last_BB_reg <= bb_2_predecessor_in_state_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_last_state <= 0;
		end else begin
			if (andOp_183_out) begin
				state_5_last_state <= 32'd4;
			end
			if (andOp_184_out) begin
				state_5_last_state <= 32'd5;
			end
		end
	end

endmodule

