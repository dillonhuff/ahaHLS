module axi_rb(input [0:0] clk, input [0:0] rst, output [0:0] valid, output [31:0] arg_0_in_data, input [31:0] arg_0_out_data, input [0:0] arg_0_read_ready, output [0:0] arg_0_read_valid, input [0:0] arg_0_write_ready, output [0:0] arg_0_write_valid, output [7:0] arg_1_raddr, input [7:0] arg_1_rdata, output [7:0] arg_1_waddr, output [7:0] arg_1_wdata, output [0:0] arg_1_wen, output [15:0] arg_2_raddr, input [15:0] arg_2_rdata, output [15:0] arg_2_waddr, output [15:0] arg_2_wdata, output [0:0] arg_2_wen, output [15:0] arg_3_s_axi_araddr, output [1:0] arg_3_s_axi_arburst, output [7:0] arg_3_s_axi_arlen, input [0:0] arg_3_s_axi_arready, output [2:0] arg_3_s_axi_arsize, output [0:0] arg_3_s_axi_arvalid, output [15:0] arg_3_s_axi_awaddr, output [1:0] arg_3_s_axi_awburst, output [7:0] arg_3_s_axi_awlen, input [0:0] arg_3_s_axi_awready, output [2:0] arg_3_s_axi_awsize, output [0:0] arg_3_s_axi_awvalid, output [0:0] arg_3_s_axi_bready, input [0:0] arg_3_s_axi_bvalid, input [31:0] arg_3_s_axi_rdata, output [0:0] arg_3_s_axi_rready, input [0:0] arg_3_s_axi_rvalid, output [31:0] arg_3_s_axi_wdata, input [0:0] arg_3_s_axi_wready, output [3:0] arg_3_s_axi_wstrb, output [0:0] arg_3_s_axi_wvalid);

	reg [0:0] valid_reg;
	reg [31:0] arg_0_in_data_reg;
	reg [0:0] arg_0_read_valid_reg;
	reg [0:0] arg_0_write_valid_reg;
	reg [7:0] arg_1_raddr_reg;
	reg [7:0] arg_1_waddr_reg;
	reg [7:0] arg_1_wdata_reg;
	reg [0:0] arg_1_wen_reg;
	reg [15:0] arg_2_raddr_reg;
	reg [15:0] arg_2_waddr_reg;
	reg [15:0] arg_2_wdata_reg;
	reg [0:0] arg_2_wen_reg;
	reg [15:0] arg_3_s_axi_araddr_reg;
	reg [1:0] arg_3_s_axi_arburst_reg;
	reg [7:0] arg_3_s_axi_arlen_reg;
	reg [2:0] arg_3_s_axi_arsize_reg;
	reg [0:0] arg_3_s_axi_arvalid_reg;
	reg [15:0] arg_3_s_axi_awaddr_reg;
	reg [1:0] arg_3_s_axi_awburst_reg;
	reg [7:0] arg_3_s_axi_awlen_reg;
	reg [2:0] arg_3_s_axi_awsize_reg;
	reg [0:0] arg_3_s_axi_awvalid_reg;
	reg [0:0] arg_3_s_axi_bready_reg;
	reg [0:0] arg_3_s_axi_rready_reg;
	reg [31:0] arg_3_s_axi_wdata_reg;
	reg [3:0] arg_3_s_axi_wstrb_reg;
	reg [0:0] arg_3_s_axi_wvalid_reg;

	assign valid = valid_reg;
	assign arg_0_in_data = arg_0_in_data_reg;
	assign arg_0_read_valid = arg_0_read_valid_reg;
	assign arg_0_write_valid = arg_0_write_valid_reg;
	assign arg_1_raddr = arg_1_raddr_reg;
	assign arg_1_waddr = arg_1_waddr_reg;
	assign arg_1_wdata = arg_1_wdata_reg;
	assign arg_1_wen = arg_1_wen_reg;
	assign arg_2_raddr = arg_2_raddr_reg;
	assign arg_2_waddr = arg_2_waddr_reg;
	assign arg_2_wdata = arg_2_wdata_reg;
	assign arg_2_wen = arg_2_wen_reg;
	assign arg_3_s_axi_araddr = arg_3_s_axi_araddr_reg;
	assign arg_3_s_axi_arburst = arg_3_s_axi_arburst_reg;
	assign arg_3_s_axi_arlen = arg_3_s_axi_arlen_reg;
	assign arg_3_s_axi_arsize = arg_3_s_axi_arsize_reg;
	assign arg_3_s_axi_arvalid = arg_3_s_axi_arvalid_reg;
	assign arg_3_s_axi_awaddr = arg_3_s_axi_awaddr_reg;
	assign arg_3_s_axi_awburst = arg_3_s_axi_awburst_reg;
	assign arg_3_s_axi_awlen = arg_3_s_axi_awlen_reg;
	assign arg_3_s_axi_awsize = arg_3_s_axi_awsize_reg;
	assign arg_3_s_axi_awvalid = arg_3_s_axi_awvalid_reg;
	assign arg_3_s_axi_bready = arg_3_s_axi_bready_reg;
	assign arg_3_s_axi_rready = arg_3_s_axi_rready_reg;
	assign arg_3_s_axi_wdata = arg_3_s_axi_wdata_reg;
	assign arg_3_s_axi_wstrb = arg_3_s_axi_wstrb_reg;
	assign arg_3_s_axi_wvalid = arg_3_s_axi_wvalid_reg;

	// Start debug wires and ports

	initial begin
	end





	// End debug wires and ports

	// Start Functional Units
	br_dummy br_unit();

	wire [31:0] sext_sext10_in;
	wire [63:0] sext_sext10_out;
	sext sext_sext10(.in(sext_sext10_in), .out(sext_sext10_out));

	wire [31:0] icmp_icmp11_in0;
	wire [31:0] icmp_icmp11_in1;
	wire [0:0] icmp_icmp11_out;
	eq #(.WIDTH(32)) icmp_icmp11(.in0(icmp_icmp11_in0), .in1(icmp_icmp11_in1), .out(icmp_icmp11_out));

	wire [31:0] sext_sext14_in;
	wire [63:0] sext_sext14_out;
	sext sext_sext14(.in(sext_sext14_in), .out(sext_sext14_out));

	wire [31:0] icmp_icmp16_in0;
	wire [31:0] icmp_icmp16_in1;
	wire [0:0] icmp_icmp16_out;
	eq #(.WIDTH(32)) icmp_icmp16(.in0(icmp_icmp16_in0), .in1(icmp_icmp16_in1), .out(icmp_icmp16_out));

	wire [31:0] sext_sext25_in;
	wire [63:0] sext_sext25_out;
	sext sext_sext25(.in(sext_sext25_in), .out(sext_sext25_out));

	wire [31:0] icmp_icmp26_in0;
	wire [31:0] icmp_icmp26_in1;
	wire [0:0] icmp_icmp26_out;
	eq #(.WIDTH(32)) icmp_icmp26(.in0(icmp_icmp26_in0), .in1(icmp_icmp26_in1), .out(icmp_icmp26_out));

	wire [31:0] sext_sext28_in;
	wire [63:0] sext_sext28_out;
	sext sext_sext28(.in(sext_sext28_in), .out(sext_sext28_out));

	wire [31:0] add_add29_in0;
	wire [31:0] add_add29_in1;
	wire [31:0] add_add29_out;
	add #(.WIDTH(32)) add_add29(.in0(add_add29_in0), .in1(add_add29_in1), .out(add_add29_out));

	wire [7:0] icmp_icmp32_in0;
	wire [7:0] icmp_icmp32_in1;
	wire [0:0] icmp_icmp32_out;
	slt #(.WIDTH(8)) icmp_icmp32(.in0(icmp_icmp32_in0), .in1(icmp_icmp32_in1), .out(icmp_icmp32_out));

	wire [31:0] trunc_trunc30_in;
	wire [7:0] trunc_trunc30_out;
	trunc #(.IN_WIDTH(32), .OUT_WIDTH(8)) trunc_trunc30(.in(trunc_trunc30_in), .out(trunc_trunc30_out));

	wire [15:0] phi_phi18_in;
	wire [31:0] phi_phi18_last_block;
	wire [63:0] phi_phi18_s;
	wire [31:0] phi_phi18_out;
	phi #(.NB_PAIR(2), .WIDTH(8)) phi_phi18(.in(phi_phi18_in), .last_block(phi_phi18_last_block), .out(phi_phi18_out), .s(phi_phi18_s));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] bb_1_active_in_state_0_in_data;
	wire [0:0] bb_1_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_0(.in_data(bb_1_active_in_state_0_in_data), .out_data(bb_1_active_in_state_0_out_data));

	reg [31:0] bb_1_predecessor_in_state_0_in_data;
	wire [31:0] bb_1_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_0(.in_data(bb_1_predecessor_in_state_0_in_data), .out_data(bb_1_predecessor_in_state_0_out_data));

	reg [0:0] br_1_happened_in_state_0_in_data;
	wire [0:0] br_1_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened_in_state_0(.in_data(br_1_happened_in_state_0_in_data), .out_data(br_1_happened_in_state_0_out_data));

	reg [0:0] bb_5_active_in_state_0_in_data;
	wire [0:0] bb_5_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_5_active_in_state_0(.in_data(bb_5_active_in_state_0_in_data), .out_data(bb_5_active_in_state_0_out_data));

	reg [31:0] bb_5_predecessor_in_state_0_in_data;
	wire [31:0] bb_5_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_5_predecessor_in_state_0(.in_data(bb_5_predecessor_in_state_0_in_data), .out_data(bb_5_predecessor_in_state_0_out_data));

	reg [0:0] br_5_happened_in_state_0_in_data;
	wire [0:0] br_5_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_5_happened_in_state_0(.in_data(br_5_happened_in_state_0_in_data), .out_data(br_5_happened_in_state_0_out_data));

	reg [0:0] bb_4_active_in_state_0_in_data;
	wire [0:0] bb_4_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_0(.in_data(bb_4_active_in_state_0_in_data), .out_data(bb_4_active_in_state_0_out_data));

	reg [31:0] bb_4_predecessor_in_state_0_in_data;
	wire [31:0] bb_4_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_0(.in_data(bb_4_predecessor_in_state_0_in_data), .out_data(bb_4_predecessor_in_state_0_out_data));

	reg [0:0] br_4_happened_in_state_0_in_data;
	wire [0:0] br_4_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_0(.in_data(br_4_happened_in_state_0_in_data), .out_data(br_4_happened_in_state_0_out_data));

	reg [0:0] bb_3_active_in_state_0_in_data;
	wire [0:0] bb_3_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_0(.in_data(bb_3_active_in_state_0_in_data), .out_data(bb_3_active_in_state_0_out_data));

	reg [31:0] bb_3_predecessor_in_state_0_in_data;
	wire [31:0] bb_3_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_0(.in_data(bb_3_predecessor_in_state_0_in_data), .out_data(bb_3_predecessor_in_state_0_out_data));

	reg [0:0] br_3_happened_in_state_0_in_data;
	wire [0:0] br_3_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_0(.in_data(br_3_happened_in_state_0_in_data), .out_data(br_3_happened_in_state_0_out_data));

	reg [0:0] bb_6_active_in_state_1_in_data;
	wire [0:0] bb_6_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_6_active_in_state_1(.in_data(bb_6_active_in_state_1_in_data), .out_data(bb_6_active_in_state_1_out_data));

	reg [31:0] bb_6_predecessor_in_state_1_in_data;
	wire [31:0] bb_6_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_6_predecessor_in_state_1(.in_data(bb_6_predecessor_in_state_1_in_data), .out_data(bb_6_predecessor_in_state_1_out_data));

	reg [0:0] br_6_happened_in_state_1_in_data;
	wire [0:0] br_6_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_6_happened_in_state_1(.in_data(br_6_happened_in_state_1_in_data), .out_data(br_6_happened_in_state_1_out_data));

	reg [0:0] bb_7_active_in_state_1_in_data;
	wire [0:0] bb_7_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_7_active_in_state_1(.in_data(bb_7_active_in_state_1_in_data), .out_data(bb_7_active_in_state_1_out_data));

	reg [31:0] bb_7_predecessor_in_state_1_in_data;
	wire [31:0] bb_7_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_7_predecessor_in_state_1(.in_data(bb_7_predecessor_in_state_1_in_data), .out_data(bb_7_predecessor_in_state_1_out_data));

	reg [0:0] br_7_happened_in_state_1_in_data;
	wire [0:0] br_7_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_7_happened_in_state_1(.in_data(br_7_happened_in_state_1_in_data), .out_data(br_7_happened_in_state_1_out_data));

	reg [0:0] bb_8_active_in_state_1_in_data;
	wire [0:0] bb_8_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active_in_state_1(.in_data(bb_8_active_in_state_1_in_data), .out_data(bb_8_active_in_state_1_out_data));

	reg [31:0] bb_8_predecessor_in_state_1_in_data;
	wire [31:0] bb_8_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor_in_state_1(.in_data(bb_8_predecessor_in_state_1_in_data), .out_data(bb_8_predecessor_in_state_1_out_data));

	reg [0:0] br_8_happened_in_state_1_in_data;
	wire [0:0] br_8_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_8_happened_in_state_1(.in_data(br_8_happened_in_state_1_in_data), .out_data(br_8_happened_in_state_1_out_data));

	reg [0:0] bb_2_active_in_state_2_in_data;
	wire [0:0] bb_2_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_2(.in_data(bb_2_active_in_state_2_in_data), .out_data(bb_2_active_in_state_2_out_data));

	reg [31:0] bb_2_predecessor_in_state_2_in_data;
	wire [31:0] bb_2_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_2(.in_data(bb_2_predecessor_in_state_2_in_data), .out_data(bb_2_predecessor_in_state_2_out_data));

	reg [0:0] bb_8_active_in_state_2_in_data;
	wire [0:0] bb_8_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active_in_state_2(.in_data(bb_8_active_in_state_2_in_data), .out_data(bb_8_active_in_state_2_out_data));

	reg [31:0] bb_8_predecessor_in_state_2_in_data;
	wire [31:0] bb_8_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor_in_state_2(.in_data(bb_8_predecessor_in_state_2_in_data), .out_data(bb_8_predecessor_in_state_2_out_data));

	reg [0:0] br_8_happened_in_state_2_in_data;
	wire [0:0] br_8_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_8_happened_in_state_2(.in_data(br_8_happened_in_state_2_in_data), .out_data(br_8_happened_in_state_2_out_data));

	reg [7:0] data_in_0_1_in_data;
	wire [7:0] data_in_0_1_out_data;
	hls_wire #(.WIDTH(8)) data_in_0_1(.in_data(data_in_0_1_in_data), .out_data(data_in_0_1_out_data));

	reg [15:0] data_in_0_3_in_data;
	wire [15:0] data_in_0_3_out_data;
	hls_wire #(.WIDTH(16)) data_in_0_3(.in_data(data_in_0_3_in_data), .out_data(data_in_0_3_out_data));

	reg [31:0] data_in_0_5_in_data;
	wire [31:0] data_in_0_5_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_5(.in_data(data_in_0_5_in_data), .out_data(data_in_0_5_out_data));

	reg [7:0] data_in_0_7_in_data;
	wire [7:0] data_in_0_7_out_data;
	hls_wire #(.WIDTH(8)) data_in_0_7(.in_data(data_in_0_7_in_data), .out_data(data_in_0_7_out_data));

	reg [7:0] data_in_0_9_in_data;
	wire [7:0] data_in_0_9_out_data;
	hls_wire #(.WIDTH(8)) data_in_0_9(.in_data(data_in_0_9_in_data), .out_data(data_in_0_9_out_data));

	reg [7:0] data_in_1_11_in_data;
	wire [7:0] data_in_1_11_out_data;
	hls_wire #(.WIDTH(8)) data_in_1_11(.in_data(data_in_1_11_in_data), .out_data(data_in_1_11_out_data));

	reg [15:0] data_in_1_13_in_data;
	wire [15:0] data_in_1_13_out_data;
	hls_wire #(.WIDTH(16)) data_in_1_13(.in_data(data_in_1_13_in_data), .out_data(data_in_1_13_out_data));

	reg [31:0] data_in_1_15_in_data;
	wire [31:0] data_in_1_15_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_15(.in_data(data_in_1_15_in_data), .out_data(data_in_1_15_out_data));

	reg [7:0] data_in_1_17_in_data;
	wire [7:0] data_in_1_17_out_data;
	hls_wire #(.WIDTH(8)) data_in_1_17(.in_data(data_in_1_17_in_data), .out_data(data_in_1_17_out_data));

	reg [7:0] data_in_1_19_in_data;
	wire [7:0] data_in_1_19_out_data;
	hls_wire #(.WIDTH(8)) data_in_1_19(.in_data(data_in_1_19_in_data), .out_data(data_in_1_19_out_data));

	reg [7:0] data_in_2_21_in_data;
	wire [7:0] data_in_2_21_out_data;
	hls_wire #(.WIDTH(8)) data_in_2_21(.in_data(data_in_2_21_in_data), .out_data(data_in_2_21_out_data));

	reg [15:0] data_in_2_23_in_data;
	wire [15:0] data_in_2_23_out_data;
	hls_wire #(.WIDTH(16)) data_in_2_23(.in_data(data_in_2_23_in_data), .out_data(data_in_2_23_out_data));

	reg [31:0] data_in_2_25_in_data;
	wire [31:0] data_in_2_25_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_25(.in_data(data_in_2_25_in_data), .out_data(data_in_2_25_out_data));

	reg [7:0] data_in_2_27_in_data;
	wire [7:0] data_in_2_27_out_data;
	hls_wire #(.WIDTH(8)) data_in_2_27(.in_data(data_in_2_27_in_data), .out_data(data_in_2_27_out_data));

	reg [7:0] data_in_2_29_in_data;
	wire [7:0] data_in_2_29_out_data;
	hls_wire #(.WIDTH(8)) data_in_2_29(.in_data(data_in_2_29_in_data), .out_data(data_in_2_29_out_data));

	wire [0:0] andOp_30_in0;
	wire [0:0] andOp_30_in1;
	wire [0:0] andOp_30_out;
	andOp #(.WIDTH(1)) andOp_30(.in0(andOp_30_in0), .in1(andOp_30_in1), .out(andOp_30_out));

	wire [0:0] notOp_31_in0;
	wire [0:0] notOp_31_out;
	notOp #(.WIDTH(1)) notOp_31(.in(notOp_31_in0), .out(notOp_31_out));

	wire [0:0] andOp_32_in0;
	wire [0:0] andOp_32_in1;
	wire [0:0] andOp_32_out;
	andOp #(.WIDTH(1)) andOp_32(.in0(andOp_32_in0), .in1(andOp_32_in1), .out(andOp_32_out));

	wire [0:0] notOp_33_in0;
	wire [0:0] notOp_33_out;
	notOp #(.WIDTH(1)) notOp_33(.in(notOp_33_in0), .out(notOp_33_out));

	wire [0:0] andOp_34_in0;
	wire [0:0] andOp_34_in1;
	wire [0:0] andOp_34_out;
	andOp #(.WIDTH(1)) andOp_34(.in0(andOp_34_in0), .in1(andOp_34_in1), .out(andOp_34_out));

	wire [0:0] notOp_35_in0;
	wire [0:0] notOp_35_out;
	notOp #(.WIDTH(1)) notOp_35(.in(notOp_35_in0), .out(notOp_35_out));

	wire [0:0] andOp_36_in0;
	wire [0:0] andOp_36_in1;
	wire [0:0] andOp_36_out;
	andOp #(.WIDTH(1)) andOp_36(.in0(andOp_36_in0), .in1(andOp_36_in1), .out(andOp_36_out));

	wire [0:0] notOp_37_in0;
	wire [0:0] notOp_37_out;
	notOp #(.WIDTH(1)) notOp_37(.in(notOp_37_in0), .out(notOp_37_out));

	wire [0:0] andOp_38_in0;
	wire [0:0] andOp_38_in1;
	wire [0:0] andOp_38_out;
	andOp #(.WIDTH(1)) andOp_38(.in0(andOp_38_in0), .in1(andOp_38_in1), .out(andOp_38_out));

	wire [0:0] andOp_39_in0;
	wire [0:0] andOp_39_in1;
	wire [0:0] andOp_39_out;
	andOp #(.WIDTH(1)) andOp_39(.in0(andOp_39_in0), .in1(andOp_39_in1), .out(andOp_39_out));

	wire [0:0] notOp_40_in0;
	wire [0:0] notOp_40_out;
	notOp #(.WIDTH(1)) notOp_40(.in(notOp_40_in0), .out(notOp_40_out));

	wire [0:0] andOp_41_in0;
	wire [0:0] andOp_41_in1;
	wire [0:0] andOp_41_out;
	andOp #(.WIDTH(1)) andOp_41(.in0(andOp_41_in0), .in1(andOp_41_in1), .out(andOp_41_out));

	wire [0:0] notOp_42_in0;
	wire [0:0] notOp_42_out;
	notOp #(.WIDTH(1)) notOp_42(.in(notOp_42_in0), .out(notOp_42_out));

	wire [0:0] andOp_43_in0;
	wire [0:0] andOp_43_in1;
	wire [0:0] andOp_43_out;
	andOp #(.WIDTH(1)) andOp_43(.in0(andOp_43_in0), .in1(andOp_43_in1), .out(andOp_43_out));

	wire [0:0] notOp_44_in0;
	wire [0:0] notOp_44_out;
	notOp #(.WIDTH(1)) notOp_44(.in(notOp_44_in0), .out(notOp_44_out));

	wire [0:0] andOp_45_in0;
	wire [0:0] andOp_45_in1;
	wire [0:0] andOp_45_out;
	andOp #(.WIDTH(1)) andOp_45(.in0(andOp_45_in0), .in1(andOp_45_in1), .out(andOp_45_out));

	wire [0:0] andOp_46_in0;
	wire [0:0] andOp_46_in1;
	wire [0:0] andOp_46_out;
	andOp #(.WIDTH(1)) andOp_46(.in0(andOp_46_in0), .in1(andOp_46_in1), .out(andOp_46_out));

	wire [0:0] notOp_47_in0;
	wire [0:0] notOp_47_out;
	notOp #(.WIDTH(1)) notOp_47(.in(notOp_47_in0), .out(notOp_47_out));

	wire [0:0] andOp_48_in0;
	wire [0:0] andOp_48_in1;
	wire [0:0] andOp_48_out;
	andOp #(.WIDTH(1)) andOp_48(.in0(andOp_48_in0), .in1(andOp_48_in1), .out(andOp_48_out));

	wire [0:0] notOp_49_in0;
	wire [0:0] notOp_49_out;
	notOp #(.WIDTH(1)) notOp_49(.in(notOp_49_in0), .out(notOp_49_out));

	wire [0:0] andOp_50_in0;
	wire [0:0] andOp_50_in1;
	wire [0:0] andOp_50_out;
	andOp #(.WIDTH(1)) andOp_50(.in0(andOp_50_in0), .in1(andOp_50_in1), .out(andOp_50_out));

	wire [0:0] notOp_51_in0;
	wire [0:0] notOp_51_out;
	notOp #(.WIDTH(1)) notOp_51(.in(notOp_51_in0), .out(notOp_51_out));

	wire [0:0] andOp_52_in0;
	wire [0:0] andOp_52_in1;
	wire [0:0] andOp_52_out;
	andOp #(.WIDTH(1)) andOp_52(.in0(andOp_52_in0), .in1(andOp_52_in1), .out(andOp_52_out));

	wire [0:0] andOp_53_in0;
	wire [0:0] andOp_53_in1;
	wire [0:0] andOp_53_out;
	andOp #(.WIDTH(1)) andOp_53(.in0(andOp_53_in0), .in1(andOp_53_in1), .out(andOp_53_out));

	wire [0:0] notOp_54_in0;
	wire [0:0] notOp_54_out;
	notOp #(.WIDTH(1)) notOp_54(.in(notOp_54_in0), .out(notOp_54_out));

	wire [0:0] andOp_55_in0;
	wire [0:0] andOp_55_in1;
	wire [0:0] andOp_55_out;
	andOp #(.WIDTH(1)) andOp_55(.in0(andOp_55_in0), .in1(andOp_55_in1), .out(andOp_55_out));

	wire [0:0] notOp_56_in0;
	wire [0:0] notOp_56_out;
	notOp #(.WIDTH(1)) notOp_56(.in(notOp_56_in0), .out(notOp_56_out));

	wire [0:0] andOp_57_in0;
	wire [0:0] andOp_57_in1;
	wire [0:0] andOp_57_out;
	andOp #(.WIDTH(1)) andOp_57(.in0(andOp_57_in0), .in1(andOp_57_in1), .out(andOp_57_out));

	wire [0:0] andOp_58_in0;
	wire [0:0] andOp_58_in1;
	wire [0:0] andOp_58_out;
	andOp #(.WIDTH(1)) andOp_58(.in0(andOp_58_in0), .in1(andOp_58_in1), .out(andOp_58_out));

	wire [0:0] notOp_59_in0;
	wire [0:0] notOp_59_out;
	notOp #(.WIDTH(1)) notOp_59(.in(notOp_59_in0), .out(notOp_59_out));

	wire [0:0] andOp_60_in0;
	wire [0:0] andOp_60_in1;
	wire [0:0] andOp_60_out;
	andOp #(.WIDTH(1)) andOp_60(.in0(andOp_60_in0), .in1(andOp_60_in1), .out(andOp_60_out));

	wire [0:0] notOp_61_in0;
	wire [0:0] notOp_61_out;
	notOp #(.WIDTH(1)) notOp_61(.in(notOp_61_in0), .out(notOp_61_out));

	wire [0:0] andOp_62_in0;
	wire [0:0] andOp_62_in1;
	wire [0:0] andOp_62_out;
	andOp #(.WIDTH(1)) andOp_62(.in0(andOp_62_in0), .in1(andOp_62_in1), .out(andOp_62_out));

	wire [31:0] eq_63_in0;
	wire [31:0] eq_63_in1;
	wire [0:0] eq_63_out;
	eq #(.WIDTH(32)) eq_63(.in0(eq_63_in0), .in1(eq_63_in1), .out(eq_63_out));

	wire [31:0] eq_64_in0;
	wire [31:0] eq_64_in1;
	wire [0:0] eq_64_out;
	eq #(.WIDTH(32)) eq_64(.in0(eq_64_in0), .in1(eq_64_in1), .out(eq_64_out));

	wire [0:0] orOp_65_in0;
	wire [0:0] orOp_65_in1;
	wire [0:0] orOp_65_out;
	orOp #(.WIDTH(1)) orOp_65(.in0(orOp_65_in0), .in1(orOp_65_in1), .out(orOp_65_out));

	wire [31:0] eq_66_in0;
	wire [31:0] eq_66_in1;
	wire [0:0] eq_66_out;
	eq #(.WIDTH(32)) eq_66(.in0(eq_66_in0), .in1(eq_66_in1), .out(eq_66_out));

	wire [0:0] orOp_67_in0;
	wire [0:0] orOp_67_in1;
	wire [0:0] orOp_67_out;
	orOp #(.WIDTH(1)) orOp_67(.in0(orOp_67_in0), .in1(orOp_67_in1), .out(orOp_67_out));

	wire [31:0] eq_68_in0;
	wire [31:0] eq_68_in1;
	wire [0:0] eq_68_out;
	eq #(.WIDTH(32)) eq_68(.in0(eq_68_in0), .in1(eq_68_in1), .out(eq_68_out));

	wire [0:0] orOp_69_in0;
	wire [0:0] orOp_69_in1;
	wire [0:0] orOp_69_out;
	orOp #(.WIDTH(1)) orOp_69(.in0(orOp_69_in0), .in1(orOp_69_in1), .out(orOp_69_out));

	wire [31:0] eq_70_in0;
	wire [31:0] eq_70_in1;
	wire [0:0] eq_70_out;
	eq #(.WIDTH(32)) eq_70(.in0(eq_70_in0), .in1(eq_70_in1), .out(eq_70_out));

	wire [0:0] orOp_71_in0;
	wire [0:0] orOp_71_in1;
	wire [0:0] orOp_71_out;
	orOp #(.WIDTH(1)) orOp_71(.in0(orOp_71_in0), .in1(orOp_71_in1), .out(orOp_71_out));

	wire [31:0] eq_72_in0;
	wire [31:0] eq_72_in1;
	wire [0:0] eq_72_out;
	eq #(.WIDTH(32)) eq_72(.in0(eq_72_in0), .in1(eq_72_in1), .out(eq_72_out));

	wire [31:0] eq_73_in0;
	wire [31:0] eq_73_in1;
	wire [0:0] eq_73_out;
	eq #(.WIDTH(32)) eq_73(.in0(eq_73_in0), .in1(eq_73_in1), .out(eq_73_out));

	wire [0:0] orOp_74_in0;
	wire [0:0] orOp_74_in1;
	wire [0:0] orOp_74_out;
	orOp #(.WIDTH(1)) orOp_74(.in0(orOp_74_in0), .in1(orOp_74_in1), .out(orOp_74_out));

	wire [31:0] eq_75_in0;
	wire [31:0] eq_75_in1;
	wire [0:0] eq_75_out;
	eq #(.WIDTH(32)) eq_75(.in0(eq_75_in0), .in1(eq_75_in1), .out(eq_75_out));

	wire [0:0] orOp_76_in0;
	wire [0:0] orOp_76_in1;
	wire [0:0] orOp_76_out;
	orOp #(.WIDTH(1)) orOp_76(.in0(orOp_76_in0), .in1(orOp_76_in1), .out(orOp_76_out));

	wire [31:0] eq_77_in0;
	wire [31:0] eq_77_in1;
	wire [0:0] eq_77_out;
	eq #(.WIDTH(32)) eq_77(.in0(eq_77_in0), .in1(eq_77_in1), .out(eq_77_out));

	wire [0:0] orOp_78_in0;
	wire [0:0] orOp_78_in1;
	wire [0:0] orOp_78_out;
	orOp #(.WIDTH(1)) orOp_78(.in0(orOp_78_in0), .in1(orOp_78_in1), .out(orOp_78_out));

	wire [31:0] eq_79_in0;
	wire [31:0] eq_79_in1;
	wire [0:0] eq_79_out;
	eq #(.WIDTH(32)) eq_79(.in0(eq_79_in0), .in1(eq_79_in1), .out(eq_79_out));

	wire [31:0] eq_80_in0;
	wire [31:0] eq_80_in1;
	wire [0:0] eq_80_out;
	eq #(.WIDTH(32)) eq_80(.in0(eq_80_in0), .in1(eq_80_in1), .out(eq_80_out));

	wire [31:0] eq_81_in0;
	wire [31:0] eq_81_in1;
	wire [0:0] eq_81_out;
	eq #(.WIDTH(32)) eq_81(.in0(eq_81_in0), .in1(eq_81_in1), .out(eq_81_out));

	wire [0:0] notOp_82_in0;
	wire [0:0] notOp_82_out;
	notOp #(.WIDTH(1)) notOp_82(.in(notOp_82_in0), .out(notOp_82_out));

	wire [0:0] andOp_83_in0;
	wire [0:0] andOp_83_in1;
	wire [0:0] andOp_83_out;
	andOp #(.WIDTH(1)) andOp_83(.in0(andOp_83_in0), .in1(andOp_83_in1), .out(andOp_83_out));

	wire [31:0] eq_84_in0;
	wire [31:0] eq_84_in1;
	wire [0:0] eq_84_out;
	eq #(.WIDTH(32)) eq_84(.in0(eq_84_in0), .in1(eq_84_in1), .out(eq_84_out));

	wire [0:0] notOp_85_in0;
	wire [0:0] notOp_85_out;
	notOp #(.WIDTH(1)) notOp_85(.in(notOp_85_in0), .out(notOp_85_out));

	wire [0:0] andOp_86_in0;
	wire [0:0] andOp_86_in1;
	wire [0:0] andOp_86_out;
	andOp #(.WIDTH(1)) andOp_86(.in0(andOp_86_in0), .in1(andOp_86_in1), .out(andOp_86_out));

	wire [31:0] eq_87_in0;
	wire [31:0] eq_87_in1;
	wire [0:0] eq_87_out;
	eq #(.WIDTH(32)) eq_87(.in0(eq_87_in0), .in1(eq_87_in1), .out(eq_87_out));

	wire [0:0] notOp_88_in0;
	wire [0:0] notOp_88_out;
	notOp #(.WIDTH(1)) notOp_88(.in(notOp_88_in0), .out(notOp_88_out));

	wire [0:0] andOp_89_in0;
	wire [0:0] andOp_89_in1;
	wire [0:0] andOp_89_out;
	andOp #(.WIDTH(1)) andOp_89(.in0(andOp_89_in0), .in1(andOp_89_in1), .out(andOp_89_out));

	wire [31:0] eq_90_in0;
	wire [31:0] eq_90_in1;
	wire [0:0] eq_90_out;
	eq #(.WIDTH(32)) eq_90(.in0(eq_90_in0), .in1(eq_90_in1), .out(eq_90_out));

	wire [0:0] notOp_91_in0;
	wire [0:0] notOp_91_out;
	notOp #(.WIDTH(1)) notOp_91(.in(notOp_91_in0), .out(notOp_91_out));

	wire [0:0] andOp_92_in0;
	wire [0:0] andOp_92_in1;
	wire [0:0] andOp_92_out;
	andOp #(.WIDTH(1)) andOp_92(.in0(andOp_92_in0), .in1(andOp_92_in1), .out(andOp_92_out));

	wire [31:0] eq_93_in0;
	wire [31:0] eq_93_in1;
	wire [0:0] eq_93_out;
	eq #(.WIDTH(32)) eq_93(.in0(eq_93_in0), .in1(eq_93_in1), .out(eq_93_out));

	wire [31:0] eq_94_in0;
	wire [31:0] eq_94_in1;
	wire [0:0] eq_94_out;
	eq #(.WIDTH(32)) eq_94(.in0(eq_94_in0), .in1(eq_94_in1), .out(eq_94_out));

	wire [0:0] notOp_95_in0;
	wire [0:0] notOp_95_out;
	notOp #(.WIDTH(1)) notOp_95(.in(notOp_95_in0), .out(notOp_95_out));

	wire [0:0] andOp_96_in0;
	wire [0:0] andOp_96_in1;
	wire [0:0] andOp_96_out;
	andOp #(.WIDTH(1)) andOp_96(.in0(andOp_96_in0), .in1(andOp_96_in1), .out(andOp_96_out));

	wire [31:0] eq_97_in0;
	wire [31:0] eq_97_in1;
	wire [0:0] eq_97_out;
	eq #(.WIDTH(32)) eq_97(.in0(eq_97_in0), .in1(eq_97_in1), .out(eq_97_out));

	wire [0:0] notOp_98_in0;
	wire [0:0] notOp_98_out;
	notOp #(.WIDTH(1)) notOp_98(.in(notOp_98_in0), .out(notOp_98_out));

	wire [0:0] andOp_99_in0;
	wire [0:0] andOp_99_in1;
	wire [0:0] andOp_99_out;
	andOp #(.WIDTH(1)) andOp_99(.in0(andOp_99_in0), .in1(andOp_99_in1), .out(andOp_99_out));

	wire [31:0] eq_100_in0;
	wire [31:0] eq_100_in1;
	wire [0:0] eq_100_out;
	eq #(.WIDTH(32)) eq_100(.in0(eq_100_in0), .in1(eq_100_in1), .out(eq_100_out));

	wire [0:0] notOp_101_in0;
	wire [0:0] notOp_101_out;
	notOp #(.WIDTH(1)) notOp_101(.in(notOp_101_in0), .out(notOp_101_out));

	wire [0:0] andOp_102_in0;
	wire [0:0] andOp_102_in1;
	wire [0:0] andOp_102_out;
	andOp #(.WIDTH(1)) andOp_102(.in0(andOp_102_in0), .in1(andOp_102_in1), .out(andOp_102_out));

	wire [31:0] eq_103_in0;
	wire [31:0] eq_103_in1;
	wire [0:0] eq_103_out;
	eq #(.WIDTH(32)) eq_103(.in0(eq_103_in0), .in1(eq_103_in1), .out(eq_103_out));

	wire [0:0] andOp_104_in0;
	wire [0:0] andOp_104_in1;
	wire [0:0] andOp_104_out;
	andOp #(.WIDTH(1)) andOp_104(.in0(andOp_104_in0), .in1(andOp_104_in1), .out(andOp_104_out));

	wire [0:0] andOp_105_in0;
	wire [0:0] andOp_105_in1;
	wire [0:0] andOp_105_out;
	andOp #(.WIDTH(1)) andOp_105(.in0(andOp_105_in0), .in1(andOp_105_in1), .out(andOp_105_out));

	wire [0:0] andOp_106_in0;
	wire [0:0] andOp_106_in1;
	wire [0:0] andOp_106_out;
	andOp #(.WIDTH(1)) andOp_106(.in0(andOp_106_in0), .in1(andOp_106_in1), .out(andOp_106_out));

	wire [0:0] andOp_107_in0;
	wire [0:0] andOp_107_in1;
	wire [0:0] andOp_107_out;
	andOp #(.WIDTH(1)) andOp_107(.in0(andOp_107_in0), .in1(andOp_107_in1), .out(andOp_107_out));

	wire [0:0] andOp_108_in0;
	wire [0:0] andOp_108_in1;
	wire [0:0] andOp_108_out;
	andOp #(.WIDTH(1)) andOp_108(.in0(andOp_108_in0), .in1(andOp_108_in1), .out(andOp_108_out));

	wire [0:0] andOp_109_in0;
	wire [0:0] andOp_109_in1;
	wire [0:0] andOp_109_out;
	andOp #(.WIDTH(1)) andOp_109(.in0(andOp_109_in0), .in1(andOp_109_in1), .out(andOp_109_out));

	wire [0:0] andOp_110_in0;
	wire [0:0] andOp_110_in1;
	wire [0:0] andOp_110_out;
	andOp #(.WIDTH(1)) andOp_110(.in0(andOp_110_in0), .in1(andOp_110_in1), .out(andOp_110_out));

	reg [7:0] tmp_output_111_in_data;
	wire [7:0] tmp_output_111_out_data;
	hls_wire #(.WIDTH(8)) tmp_output_111(.in_data(tmp_output_111_in_data), .out_data(tmp_output_111_out_data));

	wire [31:0] eq_112_in0;
	wire [31:0] eq_112_in1;
	wire [0:0] eq_112_out;
	eq #(.WIDTH(32)) eq_112(.in0(eq_112_in0), .in1(eq_112_in1), .out(eq_112_out));

	wire [31:0] eq_113_in0;
	wire [31:0] eq_113_in1;
	wire [0:0] eq_113_out;
	eq #(.WIDTH(32)) eq_113(.in0(eq_113_in0), .in1(eq_113_in1), .out(eq_113_out));

	wire [31:0] eq_114_in0;
	wire [31:0] eq_114_in1;
	wire [0:0] eq_114_out;
	eq #(.WIDTH(32)) eq_114(.in0(eq_114_in0), .in1(eq_114_in1), .out(eq_114_out));

	wire [31:0] eq_115_in0;
	wire [31:0] eq_115_in1;
	wire [0:0] eq_115_out;
	eq #(.WIDTH(32)) eq_115(.in0(eq_115_in0), .in1(eq_115_in1), .out(eq_115_out));

	wire [0:0] andOp_116_in0;
	wire [0:0] andOp_116_in1;
	wire [0:0] andOp_116_out;
	andOp #(.WIDTH(1)) andOp_116(.in0(andOp_116_in0), .in1(andOp_116_in1), .out(andOp_116_out));

	reg [15:0] tmp_output_117_in_data;
	wire [15:0] tmp_output_117_out_data;
	hls_wire #(.WIDTH(16)) tmp_output_117(.in_data(tmp_output_117_in_data), .out_data(tmp_output_117_out_data));

	wire [31:0] eq_118_in0;
	wire [31:0] eq_118_in1;
	wire [0:0] eq_118_out;
	eq #(.WIDTH(32)) eq_118(.in0(eq_118_in0), .in1(eq_118_in1), .out(eq_118_out));

	wire [31:0] eq_119_in0;
	wire [31:0] eq_119_in1;
	wire [0:0] eq_119_out;
	eq #(.WIDTH(32)) eq_119(.in0(eq_119_in0), .in1(eq_119_in1), .out(eq_119_out));

	wire [31:0] eq_120_in0;
	wire [31:0] eq_120_in1;
	wire [0:0] eq_120_out;
	eq #(.WIDTH(32)) eq_120(.in0(eq_120_in0), .in1(eq_120_in1), .out(eq_120_out));

	wire [31:0] eq_121_in0;
	wire [31:0] eq_121_in1;
	wire [0:0] eq_121_out;
	eq #(.WIDTH(32)) eq_121(.in0(eq_121_in0), .in1(eq_121_in1), .out(eq_121_out));

	wire [0:0] andOp_122_in0;
	wire [0:0] andOp_122_in1;
	wire [0:0] andOp_122_out;
	andOp #(.WIDTH(1)) andOp_122(.in0(andOp_122_in0), .in1(andOp_122_in1), .out(andOp_122_out));

	wire [0:0] andOp_123_in0;
	wire [0:0] andOp_123_in1;
	wire [0:0] andOp_123_out;
	andOp #(.WIDTH(1)) andOp_123(.in0(andOp_123_in0), .in1(andOp_123_in1), .out(andOp_123_out));

	wire [0:0] andOp_124_in0;
	wire [0:0] andOp_124_in1;
	wire [0:0] andOp_124_out;
	andOp #(.WIDTH(1)) andOp_124(.in0(andOp_124_in0), .in1(andOp_124_in1), .out(andOp_124_out));

	wire [0:0] andOp_125_in0;
	wire [0:0] andOp_125_in1;
	wire [0:0] andOp_125_out;
	andOp #(.WIDTH(1)) andOp_125(.in0(andOp_125_in0), .in1(andOp_125_in1), .out(andOp_125_out));

	wire [0:0] andOp_126_in0;
	wire [0:0] andOp_126_in1;
	wire [0:0] andOp_126_out;
	andOp #(.WIDTH(1)) andOp_126(.in0(andOp_126_in0), .in1(andOp_126_in1), .out(andOp_126_out));

	wire [0:0] andOp_127_in0;
	wire [0:0] andOp_127_in1;
	wire [0:0] andOp_127_out;
	andOp #(.WIDTH(1)) andOp_127(.in0(andOp_127_in0), .in1(andOp_127_in1), .out(andOp_127_out));

	wire [0:0] andOp_128_in0;
	wire [0:0] andOp_128_in1;
	wire [0:0] andOp_128_out;
	andOp #(.WIDTH(1)) andOp_128(.in0(andOp_128_in0), .in1(andOp_128_in1), .out(andOp_128_out));

	wire [0:0] andOp_129_in0;
	wire [0:0] andOp_129_in1;
	wire [0:0] andOp_129_out;
	andOp #(.WIDTH(1)) andOp_129(.in0(andOp_129_in0), .in1(andOp_129_in1), .out(andOp_129_out));

	wire [7:0] concat_130_in0;
	wire [7:0] concat_130_in1;
	wire [15:0] concat_130_out;
	concat #(.IN0_WIDTH(8), .IN1_WIDTH(8)) concat_130(.in0(concat_130_in0), .in1(concat_130_in1), .out(concat_130_out));

	wire [31:0] concat_131_in0;
	wire [31:0] concat_131_in1;
	wire [63:0] concat_131_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_131(.in0(concat_131_in0), .in1(concat_131_in1), .out(concat_131_out));

	wire [0:0] andOp_132_in0;
	wire [0:0] andOp_132_in1;
	wire [0:0] andOp_132_out;
	andOp #(.WIDTH(1)) andOp_132(.in0(andOp_132_in0), .in1(andOp_132_in1), .out(andOp_132_out));

	wire [0:0] andOp_133_in0;
	wire [0:0] andOp_133_in1;
	wire [0:0] andOp_133_out;
	andOp #(.WIDTH(1)) andOp_133(.in0(andOp_133_in0), .in1(andOp_133_in1), .out(andOp_133_out));

	wire [0:0] andOp_134_in0;
	wire [0:0] andOp_134_in1;
	wire [0:0] andOp_134_out;
	andOp #(.WIDTH(1)) andOp_134(.in0(andOp_134_in0), .in1(andOp_134_in1), .out(andOp_134_out));

	reg [31:0] tmp_output_135_in_data;
	wire [31:0] tmp_output_135_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_135(.in_data(tmp_output_135_in_data), .out_data(tmp_output_135_out_data));

	wire [31:0] eq_136_in0;
	wire [31:0] eq_136_in1;
	wire [0:0] eq_136_out;
	eq #(.WIDTH(32)) eq_136(.in0(eq_136_in0), .in1(eq_136_in1), .out(eq_136_out));

	wire [31:0] eq_137_in0;
	wire [31:0] eq_137_in1;
	wire [0:0] eq_137_out;
	eq #(.WIDTH(32)) eq_137(.in0(eq_137_in0), .in1(eq_137_in1), .out(eq_137_out));

	wire [0:0] andOp_138_in0;
	wire [0:0] andOp_138_in1;
	wire [0:0] andOp_138_out;
	andOp #(.WIDTH(1)) andOp_138(.in0(andOp_138_in0), .in1(andOp_138_in1), .out(andOp_138_out));

	wire [0:0] andOp_139_in0;
	wire [0:0] andOp_139_in1;
	wire [0:0] andOp_139_out;
	andOp #(.WIDTH(1)) andOp_139(.in0(andOp_139_in0), .in1(andOp_139_in1), .out(andOp_139_out));

	wire [0:0] andOp_140_in0;
	wire [0:0] andOp_140_in1;
	wire [0:0] andOp_140_out;
	andOp #(.WIDTH(1)) andOp_140(.in0(andOp_140_in0), .in1(andOp_140_in1), .out(andOp_140_out));

	wire [0:0] andOp_141_in0;
	wire [0:0] andOp_141_in1;
	wire [0:0] andOp_141_out;
	andOp #(.WIDTH(1)) andOp_141(.in0(andOp_141_in0), .in1(andOp_141_in1), .out(andOp_141_out));

	wire [0:0] andOp_142_in0;
	wire [0:0] andOp_142_in1;
	wire [0:0] andOp_142_out;
	andOp #(.WIDTH(1)) andOp_142(.in0(andOp_142_in0), .in1(andOp_142_in1), .out(andOp_142_out));

	wire [0:0] andOp_143_in0;
	wire [0:0] andOp_143_in1;
	wire [0:0] andOp_143_out;
	andOp #(.WIDTH(1)) andOp_143(.in0(andOp_143_in0), .in1(andOp_143_in1), .out(andOp_143_out));

	wire [0:0] andOp_144_in0;
	wire [0:0] andOp_144_in1;
	wire [0:0] andOp_144_out;
	andOp #(.WIDTH(1)) andOp_144(.in0(andOp_144_in0), .in1(andOp_144_in1), .out(andOp_144_out));

	wire [0:0] andOp_145_in0;
	wire [0:0] andOp_145_in1;
	wire [0:0] andOp_145_out;
	andOp #(.WIDTH(1)) andOp_145(.in0(andOp_145_in0), .in1(andOp_145_in1), .out(andOp_145_out));

	wire [0:0] andOp_146_in0;
	wire [0:0] andOp_146_in1;
	wire [0:0] andOp_146_out;
	andOp #(.WIDTH(1)) andOp_146(.in0(andOp_146_in0), .in1(andOp_146_in1), .out(andOp_146_out));

	wire [0:0] notOp_147_in0;
	wire [0:0] notOp_147_out;
	notOp #(.WIDTH(1)) notOp_147(.in(notOp_147_in0), .out(notOp_147_out));

	wire [0:0] andOp_148_in0;
	wire [0:0] andOp_148_in1;
	wire [0:0] andOp_148_out;
	andOp #(.WIDTH(1)) andOp_148(.in0(andOp_148_in0), .in1(andOp_148_in1), .out(andOp_148_out));

	wire [0:0] notOp_149_in0;
	wire [0:0] notOp_149_out;
	notOp #(.WIDTH(1)) notOp_149(.in(notOp_149_in0), .out(notOp_149_out));

	wire [0:0] andOp_150_in0;
	wire [0:0] andOp_150_in1;
	wire [0:0] andOp_150_out;
	andOp #(.WIDTH(1)) andOp_150(.in0(andOp_150_in0), .in1(andOp_150_in1), .out(andOp_150_out));

	wire [0:0] notOp_151_in0;
	wire [0:0] notOp_151_out;
	notOp #(.WIDTH(1)) notOp_151(.in(notOp_151_in0), .out(notOp_151_out));

	wire [0:0] andOp_152_in0;
	wire [0:0] andOp_152_in1;
	wire [0:0] andOp_152_out;
	andOp #(.WIDTH(1)) andOp_152(.in0(andOp_152_in0), .in1(andOp_152_in1), .out(andOp_152_out));

	wire [0:0] notOp_153_in0;
	wire [0:0] notOp_153_out;
	notOp #(.WIDTH(1)) notOp_153(.in(notOp_153_in0), .out(notOp_153_out));

	wire [0:0] andOp_154_in0;
	wire [0:0] andOp_154_in1;
	wire [0:0] andOp_154_out;
	andOp #(.WIDTH(1)) andOp_154(.in0(andOp_154_in0), .in1(andOp_154_in1), .out(andOp_154_out));

	wire [0:0] notOp_155_in0;
	wire [0:0] notOp_155_out;
	notOp #(.WIDTH(1)) notOp_155(.in(notOp_155_in0), .out(notOp_155_out));

	wire [0:0] andOp_156_in0;
	wire [0:0] andOp_156_in1;
	wire [0:0] andOp_156_out;
	andOp #(.WIDTH(1)) andOp_156(.in0(andOp_156_in0), .in1(andOp_156_in1), .out(andOp_156_out));

	wire [0:0] notOp_157_in0;
	wire [0:0] notOp_157_out;
	notOp #(.WIDTH(1)) notOp_157(.in(notOp_157_in0), .out(notOp_157_out));

	wire [0:0] andOp_158_in0;
	wire [0:0] andOp_158_in1;
	wire [0:0] andOp_158_out;
	andOp #(.WIDTH(1)) andOp_158(.in0(andOp_158_in0), .in1(andOp_158_in1), .out(andOp_158_out));

	wire [0:0] notOp_159_in0;
	wire [0:0] notOp_159_out;
	notOp #(.WIDTH(1)) notOp_159(.in(notOp_159_in0), .out(notOp_159_out));

	wire [0:0] andOp_160_in0;
	wire [0:0] andOp_160_in1;
	wire [0:0] andOp_160_out;
	andOp #(.WIDTH(1)) andOp_160(.in0(andOp_160_in0), .in1(andOp_160_in1), .out(andOp_160_out));

	wire [31:0] eq_161_in0;
	wire [31:0] eq_161_in1;
	wire [0:0] eq_161_out;
	eq #(.WIDTH(32)) eq_161(.in0(eq_161_in0), .in1(eq_161_in1), .out(eq_161_out));

	wire [31:0] eq_162_in0;
	wire [31:0] eq_162_in1;
	wire [0:0] eq_162_out;
	eq #(.WIDTH(32)) eq_162(.in0(eq_162_in0), .in1(eq_162_in1), .out(eq_162_out));

	wire [0:0] andOp_163_in0;
	wire [0:0] andOp_163_in1;
	wire [0:0] andOp_163_out;
	andOp #(.WIDTH(1)) andOp_163(.in0(andOp_163_in0), .in1(andOp_163_in1), .out(andOp_163_out));

	wire [0:0] andOp_164_in0;
	wire [0:0] andOp_164_in1;
	wire [0:0] andOp_164_out;
	andOp #(.WIDTH(1)) andOp_164(.in0(andOp_164_in0), .in1(andOp_164_in1), .out(andOp_164_out));

	wire [0:0] andOp_165_in0;
	wire [0:0] andOp_165_in1;
	wire [0:0] andOp_165_out;
	andOp #(.WIDTH(1)) andOp_165(.in0(andOp_165_in0), .in1(andOp_165_in1), .out(andOp_165_out));

	wire [31:0] eq_166_in0;
	wire [31:0] eq_166_in1;
	wire [0:0] eq_166_out;
	eq #(.WIDTH(32)) eq_166(.in0(eq_166_in0), .in1(eq_166_in1), .out(eq_166_out));

	wire [31:0] eq_167_in0;
	wire [31:0] eq_167_in1;
	wire [0:0] eq_167_out;
	eq #(.WIDTH(32)) eq_167(.in0(eq_167_in0), .in1(eq_167_in1), .out(eq_167_out));

	wire [0:0] andOp_168_in0;
	wire [0:0] andOp_168_in1;
	wire [0:0] andOp_168_out;
	andOp #(.WIDTH(1)) andOp_168(.in0(andOp_168_in0), .in1(andOp_168_in1), .out(andOp_168_out));

	wire [0:0] andOp_169_in0;
	wire [0:0] andOp_169_in1;
	wire [0:0] andOp_169_out;
	andOp #(.WIDTH(1)) andOp_169(.in0(andOp_169_in0), .in1(andOp_169_in1), .out(andOp_169_out));

	wire [31:0] eq_170_in0;
	wire [31:0] eq_170_in1;
	wire [0:0] eq_170_out;
	eq #(.WIDTH(32)) eq_170(.in0(eq_170_in0), .in1(eq_170_in1), .out(eq_170_out));

	wire [31:0] eq_171_in0;
	wire [31:0] eq_171_in1;
	wire [0:0] eq_171_out;
	eq #(.WIDTH(32)) eq_171(.in0(eq_171_in0), .in1(eq_171_in1), .out(eq_171_out));

	// End Functional Units

	reg [7:0] data_store_0_0;
	reg [15:0] data_store_0_2;
	reg [31:0] data_store_0_4;
	reg [7:0] data_store_0_6;
	reg [7:0] data_store_0_8;
	reg [7:0] data_store_1_10;
	reg [15:0] data_store_1_12;
	reg [31:0] data_store_1_14;
	reg [7:0] data_store_1_16;
	reg [7:0] data_store_1_18;
	reg [7:0] data_store_2_20;
	reg [15:0] data_store_2_22;
	reg [31:0] data_store_2_24;
	reg [7:0] data_store_2_26;
	reg [7:0] data_store_2_28;
	reg [31:0] global_state;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;

	// controller for add_add29.add_add29_in0
	// controller for add_add29.add_add29_in1
	// Insensitive connections
	assign add_add29_in0 = sext_sext28_out;
	assign add_add29_in1 = 32'd1;
	// controller for andOp_102.andOp_102_in0
	// controller for andOp_102.andOp_102_in1
	// Insensitive connections
	assign andOp_102_in0 = notOp_101_out;
	assign andOp_102_in1 = andOp_57_out;
	// controller for andOp_104.andOp_104_in0
	// controller for andOp_104.andOp_104_in1
	// Insensitive connections
	assign andOp_104_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_104_in1 = state_0_is_active;
	// controller for andOp_105.andOp_105_in0
	// controller for andOp_105.andOp_105_in1
	// Insensitive connections
	assign andOp_105_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_105_in1 = state_0_is_active;
	// controller for andOp_106.andOp_106_in0
	// controller for andOp_106.andOp_106_in1
	// Insensitive connections
	assign andOp_106_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_106_in1 = state_0_is_active;
	// controller for andOp_107.andOp_107_in0
	// controller for andOp_107.andOp_107_in1
	// Insensitive connections
	assign andOp_107_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_107_in1 = state_0_is_active;
	// controller for andOp_108.andOp_108_in0
	// controller for andOp_108.andOp_108_in1
	// Insensitive connections
	assign andOp_108_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_108_in1 = state_0_is_active;
	// controller for andOp_109.andOp_109_in0
	// controller for andOp_109.andOp_109_in1
	// Insensitive connections
	assign andOp_109_in0 = bb_5_active_in_state_0_out_data;
	assign andOp_109_in1 = state_0_is_active;
	// controller for andOp_110.andOp_110_in0
	// controller for andOp_110.andOp_110_in1
	// Insensitive connections
	assign andOp_110_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_110_in1 = state_0_is_active;
	// controller for andOp_116.andOp_116_in0
	// controller for andOp_116.andOp_116_in1
	// Insensitive connections
	assign andOp_116_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_116_in1 = state_0_is_active;
	// controller for andOp_122.andOp_122_in0
	// controller for andOp_122.andOp_122_in1
	// Insensitive connections
	assign andOp_122_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_122_in1 = state_0_is_active;
	// controller for andOp_123.andOp_123_in0
	// controller for andOp_123.andOp_123_in1
	// Insensitive connections
	assign andOp_123_in0 = bb_6_active_in_state_1_out_data;
	assign andOp_123_in1 = state_1_is_active;
	// controller for andOp_124.andOp_124_in0
	// controller for andOp_124.andOp_124_in1
	// Insensitive connections
	assign andOp_124_in0 = bb_6_active_in_state_1_out_data;
	assign andOp_124_in1 = state_1_is_active;
	// controller for andOp_125.andOp_125_in0
	// controller for andOp_125.andOp_125_in1
	// Insensitive connections
	assign andOp_125_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_125_in1 = state_0_is_active;
	// controller for andOp_126.andOp_126_in0
	// controller for andOp_126.andOp_126_in1
	// Insensitive connections
	assign andOp_126_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_126_in1 = state_0_is_active;
	// controller for andOp_127.andOp_127_in0
	// controller for andOp_127.andOp_127_in1
	// Insensitive connections
	assign andOp_127_in0 = bb_5_active_in_state_0_out_data;
	assign andOp_127_in1 = state_0_is_active;
	// controller for andOp_128.andOp_128_in0
	// controller for andOp_128.andOp_128_in1
	// Insensitive connections
	assign andOp_128_in0 = bb_5_active_in_state_0_out_data;
	assign andOp_128_in1 = state_0_is_active;
	// controller for andOp_129.andOp_129_in0
	// controller for andOp_129.andOp_129_in1
	// Insensitive connections
	assign andOp_129_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_129_in1 = state_0_is_active;
	// controller for andOp_132.andOp_132_in0
	// controller for andOp_132.andOp_132_in1
	// Insensitive connections
	assign andOp_132_in0 = bb_7_active_in_state_1_out_data;
	assign andOp_132_in1 = state_1_is_active;
	// controller for andOp_133.andOp_133_in0
	// controller for andOp_133.andOp_133_in1
	// Insensitive connections
	assign andOp_133_in0 = bb_7_active_in_state_1_out_data;
	assign andOp_133_in1 = state_1_is_active;
	// controller for andOp_134.andOp_134_in0
	// controller for andOp_134.andOp_134_in1
	// Insensitive connections
	assign andOp_134_in0 = bb_7_active_in_state_1_out_data;
	assign andOp_134_in1 = state_1_is_active;
	// controller for andOp_138.andOp_138_in0
	// controller for andOp_138.andOp_138_in1
	// Insensitive connections
	assign andOp_138_in0 = bb_7_active_in_state_1_out_data;
	assign andOp_138_in1 = state_1_is_active;
	// controller for andOp_139.andOp_139_in0
	// controller for andOp_139.andOp_139_in1
	// Insensitive connections
	assign andOp_139_in0 = bb_7_active_in_state_1_out_data;
	assign andOp_139_in1 = state_1_is_active;
	// controller for andOp_140.andOp_140_in0
	// controller for andOp_140.andOp_140_in1
	// Insensitive connections
	assign andOp_140_in0 = bb_8_active_in_state_1_out_data;
	assign andOp_140_in1 = state_1_is_active;
	// controller for andOp_141.andOp_141_in0
	// controller for andOp_141.andOp_141_in1
	// Insensitive connections
	assign andOp_141_in0 = bb_8_active_in_state_1_out_data;
	assign andOp_141_in1 = state_1_is_active;
	// controller for andOp_142.andOp_142_in0
	// controller for andOp_142.andOp_142_in1
	// Insensitive connections
	assign andOp_142_in0 = bb_8_active_in_state_1_out_data;
	assign andOp_142_in1 = state_1_is_active;
	// controller for andOp_143.andOp_143_in0
	// controller for andOp_143.andOp_143_in1
	// Insensitive connections
	assign andOp_143_in0 = bb_2_active_in_state_2_out_data;
	assign andOp_143_in1 = state_2_is_active;
	// controller for andOp_144.andOp_144_in0
	// controller for andOp_144.andOp_144_in1
	// Insensitive connections
	assign andOp_144_in0 = bb_8_active_in_state_2_out_data;
	assign andOp_144_in1 = state_2_is_active;
	// controller for andOp_145.andOp_145_in0
	// controller for andOp_145.andOp_145_in1
	// Insensitive connections
	assign andOp_145_in0 = bb_8_active_in_state_1_out_data;
	assign andOp_145_in1 = state_1_is_active;
	// controller for andOp_146.andOp_146_in0
	// controller for andOp_146.andOp_146_in1
	// Insensitive connections
	assign andOp_146_in0 = bb_2_active_in_state_2_out_data;
	assign andOp_146_in1 = state_2_is_active;
	// controller for andOp_148.andOp_148_in0
	// controller for andOp_148.andOp_148_in1
	// Insensitive connections
	assign andOp_148_in0 = notOp_147_out;
	assign andOp_148_in1 = 1'd1;
	// controller for andOp_150.andOp_150_in0
	// controller for andOp_150.andOp_150_in1
	// Insensitive connections
	assign andOp_150_in0 = notOp_149_out;
	assign andOp_150_in1 = andOp_148_out;
	// controller for andOp_152.andOp_152_in0
	// controller for andOp_152.andOp_152_in1
	// Insensitive connections
	assign andOp_152_in0 = notOp_151_out;
	assign andOp_152_in1 = andOp_150_out;
	// controller for andOp_154.andOp_154_in0
	// controller for andOp_154.andOp_154_in1
	// Insensitive connections
	assign andOp_154_in0 = notOp_153_out;
	assign andOp_154_in1 = 1'd1;
	// controller for andOp_156.andOp_156_in0
	// controller for andOp_156.andOp_156_in1
	// Insensitive connections
	assign andOp_156_in0 = notOp_155_out;
	assign andOp_156_in1 = andOp_154_out;
	// controller for andOp_158.andOp_158_in0
	// controller for andOp_158.andOp_158_in1
	// Insensitive connections
	assign andOp_158_in0 = notOp_157_out;
	assign andOp_158_in1 = 1'd1;
	// controller for andOp_160.andOp_160_in0
	// controller for andOp_160.andOp_160_in1
	// Insensitive connections
	assign andOp_160_in0 = notOp_159_out;
	assign andOp_160_in1 = andOp_158_out;
	// controller for andOp_163.andOp_163_in0
	// controller for andOp_163.andOp_163_in1
	// Insensitive connections
	assign andOp_163_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_163_in1 = state_0_is_active;
	// controller for andOp_164.andOp_164_in0
	// controller for andOp_164.andOp_164_in1
	// Insensitive connections
	assign andOp_164_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_164_in1 = state_0_is_active;
	// controller for andOp_165.andOp_165_in0
	// controller for andOp_165.andOp_165_in1
	// Insensitive connections
	assign andOp_165_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_165_in1 = state_0_is_active;
	// controller for andOp_168.andOp_168_in0
	// controller for andOp_168.andOp_168_in1
	// Insensitive connections
	assign andOp_168_in0 = bb_6_active_in_state_1_out_data;
	assign andOp_168_in1 = state_1_is_active;
	// controller for andOp_169.andOp_169_in0
	// controller for andOp_169.andOp_169_in1
	// Insensitive connections
	assign andOp_169_in0 = bb_8_active_in_state_1_out_data;
	assign andOp_169_in1 = state_1_is_active;
	// controller for andOp_30.andOp_30_in0
	// controller for andOp_30.andOp_30_in1
	// Insensitive connections
	assign andOp_30_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_30_in1 = state_0_is_active;
	// controller for andOp_32.andOp_32_in0
	// controller for andOp_32.andOp_32_in1
	// Insensitive connections
	assign andOp_32_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_32_in1 = state_0_is_active;
	// controller for andOp_34.andOp_34_in0
	// controller for andOp_34.andOp_34_in1
	// Insensitive connections
	assign andOp_34_in0 = bb_5_active_in_state_0_out_data;
	assign andOp_34_in1 = state_0_is_active;
	// controller for andOp_36.andOp_36_in0
	// controller for andOp_36.andOp_36_in1
	// Insensitive connections
	assign andOp_36_in0 = andOp_34_out;
	assign andOp_36_in1 = icmp_icmp16_out;
	// controller for andOp_38.andOp_38_in0
	// controller for andOp_38.andOp_38_in1
	// Insensitive connections
	assign andOp_38_in0 = andOp_34_out;
	assign andOp_38_in1 = notOp_37_out;
	// controller for andOp_39.andOp_39_in0
	// controller for andOp_39.andOp_39_in1
	// Insensitive connections
	assign andOp_39_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_39_in1 = state_0_is_active;
	// controller for andOp_41.andOp_41_in0
	// controller for andOp_41.andOp_41_in1
	// Insensitive connections
	assign andOp_41_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_41_in1 = state_0_is_active;
	// controller for andOp_43.andOp_43_in0
	// controller for andOp_43.andOp_43_in1
	// Insensitive connections
	assign andOp_43_in0 = andOp_41_out;
	assign andOp_43_in1 = icmp_icmp11_out;
	// controller for andOp_45.andOp_45_in0
	// controller for andOp_45.andOp_45_in1
	// Insensitive connections
	assign andOp_45_in0 = andOp_41_out;
	assign andOp_45_in1 = notOp_44_out;
	// controller for andOp_46.andOp_46_in0
	// controller for andOp_46.andOp_46_in1
	// Insensitive connections
	assign andOp_46_in0 = bb_6_active_in_state_1_out_data;
	assign andOp_46_in1 = state_1_is_active;
	// controller for andOp_48.andOp_48_in0
	// controller for andOp_48.andOp_48_in1
	// Insensitive connections
	assign andOp_48_in0 = bb_7_active_in_state_1_out_data;
	assign andOp_48_in1 = state_1_is_active;
	// controller for andOp_50.andOp_50_in0
	// controller for andOp_50.andOp_50_in1
	// Insensitive connections
	assign andOp_50_in0 = andOp_48_out;
	assign andOp_50_in1 = icmp_icmp26_out;
	// controller for andOp_52.andOp_52_in0
	// controller for andOp_52.andOp_52_in1
	// Insensitive connections
	assign andOp_52_in0 = andOp_48_out;
	assign andOp_52_in1 = notOp_51_out;
	// controller for andOp_53.andOp_53_in0
	// controller for andOp_53.andOp_53_in1
	// Insensitive connections
	assign andOp_53_in0 = bb_8_active_in_state_2_out_data;
	assign andOp_53_in1 = state_2_is_active;
	// controller for andOp_55.andOp_55_in0
	// controller for andOp_55.andOp_55_in1
	// Insensitive connections
	assign andOp_55_in0 = andOp_53_out;
	assign andOp_55_in1 = icmp_icmp32_out;
	// controller for andOp_57.andOp_57_in0
	// controller for andOp_57.andOp_57_in1
	// Insensitive connections
	assign andOp_57_in0 = andOp_53_out;
	assign andOp_57_in1 = notOp_56_out;
	// controller for andOp_58.andOp_58_in0
	// controller for andOp_58.andOp_58_in1
	// Insensitive connections
	assign andOp_58_in0 = bb_8_active_in_state_2_out_data;
	assign andOp_58_in1 = state_2_is_active;
	// controller for andOp_60.andOp_60_in0
	// controller for andOp_60.andOp_60_in1
	// Insensitive connections
	assign andOp_60_in0 = andOp_58_out;
	assign andOp_60_in1 = icmp_icmp32_out;
	// controller for andOp_62.andOp_62_in0
	// controller for andOp_62.andOp_62_in1
	// Insensitive connections
	assign andOp_62_in0 = andOp_58_out;
	assign andOp_62_in1 = notOp_61_out;
	// controller for andOp_83.andOp_83_in0
	// controller for andOp_83.andOp_83_in1
	// Insensitive connections
	assign andOp_83_in0 = notOp_82_out;
	assign andOp_83_in1 = andOp_39_out;
	// controller for andOp_86.andOp_86_in0
	// controller for andOp_86.andOp_86_in1
	// Insensitive connections
	assign andOp_86_in0 = notOp_85_out;
	assign andOp_86_in1 = andOp_32_out;
	// controller for andOp_89.andOp_89_in0
	// controller for andOp_89.andOp_89_in1
	// Insensitive connections
	assign andOp_89_in0 = notOp_88_out;
	assign andOp_89_in1 = andOp_45_out;
	// controller for andOp_92.andOp_92_in0
	// controller for andOp_92.andOp_92_in1
	// Insensitive connections
	assign andOp_92_in0 = notOp_91_out;
	assign andOp_92_in1 = andOp_30_out;
	// controller for andOp_96.andOp_96_in0
	// controller for andOp_96.andOp_96_in1
	// Insensitive connections
	assign andOp_96_in0 = notOp_95_out;
	assign andOp_96_in1 = andOp_46_out;
	// controller for andOp_99.andOp_99_in0
	// controller for andOp_99.andOp_99_in1
	// Insensitive connections
	assign andOp_99_in0 = notOp_98_out;
	assign andOp_99_in1 = andOp_52_out;
	// controller for arg_0.arg_0_in_data_reg
	always @(*) begin
		if (andOp_134_out) begin 
			arg_0_in_data_reg = tmp_output_135_out_data;
		end else begin
			arg_0_in_data_reg = 0;
		end
	end
	// controller for arg_0.arg_0_write_valid_reg
	always @(*) begin
		if (andOp_133_out) begin 
			arg_0_write_valid_reg = 32'd1;
		end else begin
			arg_0_write_valid_reg = 0;
		end
	end
	// controller for arg_1.arg_1_raddr_reg
	always @(*) begin
		if (andOp_104_out) begin 
			arg_1_raddr_reg = arg_1_rdata;
		end else begin
			arg_1_raddr_reg = 0;
		end
	end
	// controller for arg_2.arg_2_raddr_reg
	always @(*) begin
		if (andOp_105_out) begin 
			arg_2_raddr_reg = arg_2_rdata;
		end else begin
			arg_2_raddr_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_araddr_reg
	always @(*) begin
		if (andOp_116_out) begin 
			arg_3_s_axi_araddr_reg = tmp_output_117_out_data;
		end else begin
			arg_3_s_axi_araddr_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_arburst_reg
	always @(*) begin
		if (andOp_108_out) begin 
			arg_3_s_axi_arburst_reg = 2'd1;
		end else begin
			arg_3_s_axi_arburst_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_arlen_reg
	always @(*) begin
		if (andOp_110_out) begin 
			arg_3_s_axi_arlen_reg = tmp_output_111_out_data;
		end else begin
			arg_3_s_axi_arlen_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_arsize_reg
	always @(*) begin
		if (andOp_107_out) begin 
			arg_3_s_axi_arsize_reg = -(3'd3);
		end else begin
			arg_3_s_axi_arsize_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_arvalid_reg
	always @(*) begin
		if (andOp_106_out) begin 
			arg_3_s_axi_arvalid_reg = 32'd1;
		end else begin
			arg_3_s_axi_arvalid_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_rready_reg
	always @(*) begin
		if (andOp_123_out) begin 
			arg_3_s_axi_rready_reg = 32'd1;
		end else begin
			arg_3_s_axi_rready_reg = 0;
		end
	end
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_63_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_80_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_0.bb_1_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_0_in_data = orOp_65_out;
		end else begin
			bb_1_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_0.bb_1_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_83_out) begin 
			bb_1_predecessor_in_state_0_in_data = 32'd4;
		end else if (eq_81_out) begin 
			bb_1_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_2.bb_2_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_2_in_data = orOp_78_out;
		end else begin
			bb_2_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_2.bb_2_predecessor_in_state_2_in_data
	always @(*) begin
		if (andOp_102_out) begin 
			bb_2_predecessor_in_state_2_in_data = 32'd8;
		end else if (eq_100_out) begin 
			bb_2_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_0.bb_3_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_0_in_data = orOp_71_out;
		end else begin
			bb_3_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_0.bb_3_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_92_out) begin 
			bb_3_predecessor_in_state_0_in_data = 32'd0;
		end else if (eq_90_out) begin 
			bb_3_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_0.bb_4_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_0_in_data = orOp_69_out;
		end else begin
			bb_4_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_0.bb_4_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_89_out) begin 
			bb_4_predecessor_in_state_0_in_data = 32'd3;
		end else if (eq_87_out) begin 
			bb_4_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_5_active_in_state_0.bb_5_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_5_active_in_state_0_in_data = orOp_67_out;
		end else begin
			bb_5_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_5_predecessor_in_state_0.bb_5_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_86_out) begin 
			bb_5_predecessor_in_state_0_in_data = 32'd1;
		end else if (eq_84_out) begin 
			bb_5_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_5_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_6_active_in_state_1.bb_6_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_6_active_in_state_1_in_data = eq_72_out;
		end else begin
			bb_6_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_6_predecessor_in_state_1.bb_6_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_93_out) begin 
			bb_6_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_6_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_7_active_in_state_1.bb_7_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_7_active_in_state_1_in_data = orOp_74_out;
		end else begin
			bb_7_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_7_predecessor_in_state_1.bb_7_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_96_out) begin 
			bb_7_predecessor_in_state_1_in_data = 32'd6;
		end else if (eq_94_out) begin 
			bb_7_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_7_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_8_active_in_state_1.bb_8_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_state_1_in_data = orOp_76_out;
		end else begin
			bb_8_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_8_active_in_state_2.bb_8_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_state_2_in_data = eq_79_out;
		end else begin
			bb_8_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_8_predecessor_in_state_1.bb_8_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_99_out) begin 
			bb_8_predecessor_in_state_1_in_data = 32'd7;
		end else if (eq_97_out) begin 
			bb_8_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_8_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_8_predecessor_in_state_2.bb_8_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_103_out) begin 
			bb_8_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_8_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_30_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_31_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_1_happened_in_state_0.br_1_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_32_out) begin 
			br_1_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_33_out) begin 
			br_1_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_1_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_0.br_3_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_41_out) begin 
			br_3_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_42_out) begin 
			br_3_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_0.br_4_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_39_out) begin 
			br_4_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_40_out) begin 
			br_4_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_5_happened_in_state_0.br_5_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_34_out) begin 
			br_5_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_35_out) begin 
			br_5_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_5_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_6_happened_in_state_1.br_6_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_46_out) begin 
			br_6_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_47_out) begin 
			br_6_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_6_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_7_happened_in_state_1.br_7_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_48_out) begin 
			br_7_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_49_out) begin 
			br_7_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_7_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_8_happened_in_state_1.br_8_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_53_out) begin 
			br_8_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_54_out) begin 
			br_8_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_8_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_8_happened_in_state_2.br_8_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_58_out) begin 
			br_8_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_59_out) begin 
			br_8_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_8_happened_in_state_2_in_data = 0;
		end
	end
	// controller for concat_130.concat_130_in0
	// controller for concat_130.concat_130_in1
	// Insensitive connections
	assign concat_130_in0 = 8'd0;
	assign concat_130_in1 = data_in_0_7_out_data;
	// controller for concat_131.concat_131_in0
	// controller for concat_131.concat_131_in1
	// Insensitive connections
	assign concat_131_in0 = 32'd4;
	assign concat_131_in1 = 32'd8;
	// controller for data_in_0_1.data_in_0_1_in_data
	always @(*) begin
		if (eq_161_out) begin 
			data_in_0_1_in_data = data_store_0_0;
		end else if (eq_162_out) begin 
			data_in_0_1_in_data = data_store_2_20;
		end else begin
			data_in_0_1_in_data = 0;
		end
	end
	// controller for data_in_0_3.data_in_0_3_in_data
	always @(*) begin
		if (eq_161_out) begin 
			data_in_0_3_in_data = data_store_0_2;
		end else if (eq_162_out) begin 
			data_in_0_3_in_data = data_store_2_22;
		end else begin
			data_in_0_3_in_data = 0;
		end
	end
	// controller for data_in_0_5.data_in_0_5_in_data
	always @(*) begin
		if (eq_161_out) begin 
			data_in_0_5_in_data = data_store_0_4;
		end else if (eq_162_out) begin 
			data_in_0_5_in_data = data_store_2_24;
		end else begin
			data_in_0_5_in_data = 0;
		end
	end
	// controller for data_in_0_7.data_in_0_7_in_data
	always @(*) begin
		if (eq_161_out) begin 
			data_in_0_7_in_data = data_store_0_6;
		end else if (eq_162_out) begin 
			data_in_0_7_in_data = data_store_2_26;
		end else begin
			data_in_0_7_in_data = 0;
		end
	end
	// controller for data_in_0_9.data_in_0_9_in_data
	always @(*) begin
		if (eq_161_out) begin 
			data_in_0_9_in_data = data_store_0_8;
		end else if (eq_162_out) begin 
			data_in_0_9_in_data = data_store_2_28;
		end else begin
			data_in_0_9_in_data = 0;
		end
	end
	// controller for data_in_1_11.data_in_1_11_in_data
	always @(*) begin
		if (eq_166_out) begin 
			data_in_1_11_in_data = data_store_0_0;
		end else if (eq_167_out) begin 
			data_in_1_11_in_data = data_store_1_10;
		end else begin
			data_in_1_11_in_data = 0;
		end
	end
	// controller for data_in_1_13.data_in_1_13_in_data
	always @(*) begin
		if (eq_166_out) begin 
			data_in_1_13_in_data = data_store_0_2;
		end else if (eq_167_out) begin 
			data_in_1_13_in_data = data_store_1_12;
		end else begin
			data_in_1_13_in_data = 0;
		end
	end
	// controller for data_in_1_15.data_in_1_15_in_data
	always @(*) begin
		if (eq_166_out) begin 
			data_in_1_15_in_data = data_store_0_4;
		end else if (eq_167_out) begin 
			data_in_1_15_in_data = data_store_1_14;
		end else begin
			data_in_1_15_in_data = 0;
		end
	end
	// controller for data_in_1_17.data_in_1_17_in_data
	always @(*) begin
		if (eq_166_out) begin 
			data_in_1_17_in_data = data_store_0_6;
		end else if (eq_167_out) begin 
			data_in_1_17_in_data = data_store_1_16;
		end else begin
			data_in_1_17_in_data = 0;
		end
	end
	// controller for data_in_1_19.data_in_1_19_in_data
	always @(*) begin
		if (eq_166_out) begin 
			data_in_1_19_in_data = data_store_0_8;
		end else if (eq_167_out) begin 
			data_in_1_19_in_data = data_store_1_18;
		end else begin
			data_in_1_19_in_data = 0;
		end
	end
	// controller for data_in_2_21.data_in_2_21_in_data
	always @(*) begin
		if (eq_170_out) begin 
			data_in_2_21_in_data = data_store_1_10;
		end else if (eq_171_out) begin 
			data_in_2_21_in_data = data_store_2_20;
		end else begin
			data_in_2_21_in_data = 0;
		end
	end
	// controller for data_in_2_23.data_in_2_23_in_data
	always @(*) begin
		if (eq_170_out) begin 
			data_in_2_23_in_data = data_store_1_12;
		end else if (eq_171_out) begin 
			data_in_2_23_in_data = data_store_2_22;
		end else begin
			data_in_2_23_in_data = 0;
		end
	end
	// controller for data_in_2_25.data_in_2_25_in_data
	always @(*) begin
		if (eq_170_out) begin 
			data_in_2_25_in_data = data_store_1_14;
		end else if (eq_171_out) begin 
			data_in_2_25_in_data = data_store_2_24;
		end else begin
			data_in_2_25_in_data = 0;
		end
	end
	// controller for data_in_2_27.data_in_2_27_in_data
	always @(*) begin
		if (eq_170_out) begin 
			data_in_2_27_in_data = data_store_1_16;
		end else if (eq_171_out) begin 
			data_in_2_27_in_data = data_store_2_26;
		end else begin
			data_in_2_27_in_data = 0;
		end
	end
	// controller for data_in_2_29.data_in_2_29_in_data
	always @(*) begin
		if (eq_170_out) begin 
			data_in_2_29_in_data = data_store_1_18;
		end else if (eq_171_out) begin 
			data_in_2_29_in_data = data_store_2_28;
		end else begin
			data_in_2_29_in_data = 0;
		end
	end
	// controller for eq_100.eq_100_in0
	// controller for eq_100.eq_100_in1
	// Insensitive connections
	assign eq_100_in0 = 32'd2;
	assign eq_100_in1 = state_2_entry_BB_reg;
	// controller for eq_103.eq_103_in0
	// controller for eq_103.eq_103_in1
	// Insensitive connections
	assign eq_103_in0 = 32'd8;
	assign eq_103_in1 = state_2_entry_BB_reg;
	// controller for eq_112.eq_112_in0
	// controller for eq_112.eq_112_in1
	// Insensitive connections
	assign eq_112_in0 = 32'd0;
	assign eq_112_in1 = state_0_entry_BB_reg;
	// controller for eq_113.eq_113_in0
	// controller for eq_113.eq_113_in1
	// Insensitive connections
	assign eq_113_in0 = 32'd1;
	assign eq_113_in1 = state_0_entry_BB_reg;
	// controller for eq_114.eq_114_in0
	// controller for eq_114.eq_114_in1
	// Insensitive connections
	assign eq_114_in0 = 32'd5;
	assign eq_114_in1 = state_0_entry_BB_reg;
	// controller for eq_115.eq_115_in0
	// controller for eq_115.eq_115_in1
	// Insensitive connections
	assign eq_115_in0 = 32'd3;
	assign eq_115_in1 = state_0_entry_BB_reg;
	// controller for eq_118.eq_118_in0
	// controller for eq_118.eq_118_in1
	// Insensitive connections
	assign eq_118_in0 = 32'd0;
	assign eq_118_in1 = state_0_entry_BB_reg;
	// controller for eq_119.eq_119_in0
	// controller for eq_119.eq_119_in1
	// Insensitive connections
	assign eq_119_in0 = 32'd1;
	assign eq_119_in1 = state_0_entry_BB_reg;
	// controller for eq_120.eq_120_in0
	// controller for eq_120.eq_120_in1
	// Insensitive connections
	assign eq_120_in0 = 32'd5;
	assign eq_120_in1 = state_0_entry_BB_reg;
	// controller for eq_121.eq_121_in0
	// controller for eq_121.eq_121_in1
	// Insensitive connections
	assign eq_121_in0 = 32'd3;
	assign eq_121_in1 = state_0_entry_BB_reg;
	// controller for eq_136.eq_136_in0
	// controller for eq_136.eq_136_in1
	// Insensitive connections
	assign eq_136_in0 = 32'd6;
	assign eq_136_in1 = state_1_entry_BB_reg;
	// controller for eq_137.eq_137_in0
	// controller for eq_137.eq_137_in1
	// Insensitive connections
	assign eq_137_in0 = 32'd7;
	assign eq_137_in1 = state_1_entry_BB_reg;
	// controller for eq_161.eq_161_in0
	// controller for eq_161.eq_161_in1
	// Insensitive connections
	assign eq_161_in0 = 32'd0;
	assign eq_161_in1 = state_0_last_state;
	// controller for eq_162.eq_162_in0
	// controller for eq_162.eq_162_in1
	// Insensitive connections
	assign eq_162_in0 = 32'd2;
	assign eq_162_in1 = state_0_last_state;
	// controller for eq_166.eq_166_in0
	// controller for eq_166.eq_166_in1
	// Insensitive connections
	assign eq_166_in0 = 32'd0;
	assign eq_166_in1 = state_1_last_state;
	// controller for eq_167.eq_167_in0
	// controller for eq_167.eq_167_in1
	// Insensitive connections
	assign eq_167_in0 = 32'd1;
	assign eq_167_in1 = state_1_last_state;
	// controller for eq_170.eq_170_in0
	// controller for eq_170.eq_170_in1
	// Insensitive connections
	assign eq_170_in0 = 32'd1;
	assign eq_170_in1 = state_2_last_state;
	// controller for eq_171.eq_171_in0
	// controller for eq_171.eq_171_in1
	// Insensitive connections
	assign eq_171_in0 = 32'd2;
	assign eq_171_in1 = state_2_last_state;
	// controller for eq_63.eq_63_in0
	// controller for eq_63.eq_63_in1
	// Insensitive connections
	assign eq_63_in0 = 32'd0;
	assign eq_63_in1 = state_0_entry_BB_reg;
	// controller for eq_64.eq_64_in0
	// controller for eq_64.eq_64_in1
	// Insensitive connections
	assign eq_64_in0 = 32'd1;
	assign eq_64_in1 = state_0_entry_BB_reg;
	// controller for eq_66.eq_66_in0
	// controller for eq_66.eq_66_in1
	// Insensitive connections
	assign eq_66_in0 = 32'd5;
	assign eq_66_in1 = state_0_entry_BB_reg;
	// controller for eq_68.eq_68_in0
	// controller for eq_68.eq_68_in1
	// Insensitive connections
	assign eq_68_in0 = 32'd4;
	assign eq_68_in1 = state_0_entry_BB_reg;
	// controller for eq_70.eq_70_in0
	// controller for eq_70.eq_70_in1
	// Insensitive connections
	assign eq_70_in0 = 32'd3;
	assign eq_70_in1 = state_0_entry_BB_reg;
	// controller for eq_72.eq_72_in0
	// controller for eq_72.eq_72_in1
	// Insensitive connections
	assign eq_72_in0 = 32'd6;
	assign eq_72_in1 = state_1_entry_BB_reg;
	// controller for eq_73.eq_73_in0
	// controller for eq_73.eq_73_in1
	// Insensitive connections
	assign eq_73_in0 = 32'd7;
	assign eq_73_in1 = state_1_entry_BB_reg;
	// controller for eq_75.eq_75_in0
	// controller for eq_75.eq_75_in1
	// Insensitive connections
	assign eq_75_in0 = 32'd8;
	assign eq_75_in1 = state_1_entry_BB_reg;
	// controller for eq_77.eq_77_in0
	// controller for eq_77.eq_77_in1
	// Insensitive connections
	assign eq_77_in0 = 32'd2;
	assign eq_77_in1 = state_2_entry_BB_reg;
	// controller for eq_79.eq_79_in0
	// controller for eq_79.eq_79_in1
	// Insensitive connections
	assign eq_79_in0 = 32'd8;
	assign eq_79_in1 = state_2_entry_BB_reg;
	// controller for eq_80.eq_80_in0
	// controller for eq_80.eq_80_in1
	// Insensitive connections
	assign eq_80_in0 = 32'd0;
	assign eq_80_in1 = state_0_entry_BB_reg;
	// controller for eq_81.eq_81_in0
	// controller for eq_81.eq_81_in1
	// Insensitive connections
	assign eq_81_in0 = 32'd1;
	assign eq_81_in1 = state_0_entry_BB_reg;
	// controller for eq_84.eq_84_in0
	// controller for eq_84.eq_84_in1
	// Insensitive connections
	assign eq_84_in0 = 32'd5;
	assign eq_84_in1 = state_0_entry_BB_reg;
	// controller for eq_87.eq_87_in0
	// controller for eq_87.eq_87_in1
	// Insensitive connections
	assign eq_87_in0 = 32'd4;
	assign eq_87_in1 = state_0_entry_BB_reg;
	// controller for eq_90.eq_90_in0
	// controller for eq_90.eq_90_in1
	// Insensitive connections
	assign eq_90_in0 = 32'd3;
	assign eq_90_in1 = state_0_entry_BB_reg;
	// controller for eq_93.eq_93_in0
	// controller for eq_93.eq_93_in1
	// Insensitive connections
	assign eq_93_in0 = 32'd6;
	assign eq_93_in1 = state_1_entry_BB_reg;
	// controller for eq_94.eq_94_in0
	// controller for eq_94.eq_94_in1
	// Insensitive connections
	assign eq_94_in0 = 32'd7;
	assign eq_94_in1 = state_1_entry_BB_reg;
	// controller for eq_97.eq_97_in0
	// controller for eq_97.eq_97_in1
	// Insensitive connections
	assign eq_97_in0 = 32'd8;
	assign eq_97_in1 = state_1_entry_BB_reg;
	// controller for icmp_icmp11.icmp_icmp11_in0
	// controller for icmp_icmp11.icmp_icmp11_in1
	// Insensitive connections
	assign icmp_icmp11_in0 = sext_sext10_out;
	assign icmp_icmp11_in1 = 32'd0;
	// controller for icmp_icmp16.icmp_icmp16_in0
	// controller for icmp_icmp16.icmp_icmp16_in1
	// Insensitive connections
	assign icmp_icmp16_in0 = sext_sext14_out;
	assign icmp_icmp16_in1 = 32'd0;
	// controller for icmp_icmp26.icmp_icmp26_in0
	// controller for icmp_icmp26.icmp_icmp26_in1
	// Insensitive connections
	assign icmp_icmp26_in0 = sext_sext25_out;
	assign icmp_icmp26_in1 = 32'd0;
	// controller for icmp_icmp32.icmp_icmp32_in0
	// controller for icmp_icmp32.icmp_icmp32_in1
	// Insensitive connections
	assign icmp_icmp32_in0 = data_in_2_27_out_data;
	assign icmp_icmp32_in1 = data_in_2_21_out_data;
	// controller for notOp_101.notOp_101_in0
	// Insensitive connections
	assign notOp_101_in0 = eq_100_out;
	// controller for notOp_147.notOp_147_in0
	// Insensitive connections
	assign notOp_147_in0 = andOp_36_out;
	// controller for notOp_149.notOp_149_in0
	// Insensitive connections
	assign notOp_149_in0 = andOp_43_out;
	// controller for notOp_151.notOp_151_in0
	// Insensitive connections
	assign notOp_151_in0 = andOp_55_out;
	// controller for notOp_153.notOp_153_in0
	// Insensitive connections
	assign notOp_153_in0 = andOp_38_out;
	// controller for notOp_155.notOp_155_in0
	// Insensitive connections
	assign notOp_155_in0 = andOp_50_out;
	// controller for notOp_157.notOp_157_in0
	// Insensitive connections
	assign notOp_157_in0 = andOp_145_out;
	// controller for notOp_159.notOp_159_in0
	// Insensitive connections
	assign notOp_159_in0 = andOp_146_out;
	// controller for notOp_31.notOp_31_in0
	// Insensitive connections
	assign notOp_31_in0 = andOp_30_out;
	// controller for notOp_33.notOp_33_in0
	// Insensitive connections
	assign notOp_33_in0 = andOp_32_out;
	// controller for notOp_35.notOp_35_in0
	// Insensitive connections
	assign notOp_35_in0 = andOp_34_out;
	// controller for notOp_37.notOp_37_in0
	// Insensitive connections
	assign notOp_37_in0 = icmp_icmp16_out;
	// controller for notOp_40.notOp_40_in0
	// Insensitive connections
	assign notOp_40_in0 = andOp_39_out;
	// controller for notOp_42.notOp_42_in0
	// Insensitive connections
	assign notOp_42_in0 = andOp_41_out;
	// controller for notOp_44.notOp_44_in0
	// Insensitive connections
	assign notOp_44_in0 = icmp_icmp11_out;
	// controller for notOp_47.notOp_47_in0
	// Insensitive connections
	assign notOp_47_in0 = andOp_46_out;
	// controller for notOp_49.notOp_49_in0
	// Insensitive connections
	assign notOp_49_in0 = andOp_48_out;
	// controller for notOp_51.notOp_51_in0
	// Insensitive connections
	assign notOp_51_in0 = icmp_icmp26_out;
	// controller for notOp_54.notOp_54_in0
	// Insensitive connections
	assign notOp_54_in0 = andOp_53_out;
	// controller for notOp_56.notOp_56_in0
	// Insensitive connections
	assign notOp_56_in0 = icmp_icmp32_out;
	// controller for notOp_59.notOp_59_in0
	// Insensitive connections
	assign notOp_59_in0 = andOp_58_out;
	// controller for notOp_61.notOp_61_in0
	// Insensitive connections
	assign notOp_61_in0 = icmp_icmp32_out;
	// controller for notOp_82.notOp_82_in0
	// Insensitive connections
	assign notOp_82_in0 = eq_81_out;
	// controller for notOp_85.notOp_85_in0
	// Insensitive connections
	assign notOp_85_in0 = eq_84_out;
	// controller for notOp_88.notOp_88_in0
	// Insensitive connections
	assign notOp_88_in0 = eq_87_out;
	// controller for notOp_91.notOp_91_in0
	// Insensitive connections
	assign notOp_91_in0 = eq_90_out;
	// controller for notOp_95.notOp_95_in0
	// Insensitive connections
	assign notOp_95_in0 = eq_94_out;
	// controller for notOp_98.notOp_98_in0
	// Insensitive connections
	assign notOp_98_in0 = eq_97_out;
	// controller for orOp_65.orOp_65_in0
	// controller for orOp_65.orOp_65_in1
	// Insensitive connections
	assign orOp_65_in0 = eq_64_out;
	assign orOp_65_in1 = andOp_39_out;
	// controller for orOp_67.orOp_67_in0
	// controller for orOp_67.orOp_67_in1
	// Insensitive connections
	assign orOp_67_in0 = eq_66_out;
	assign orOp_67_in1 = andOp_32_out;
	// controller for orOp_69.orOp_69_in0
	// controller for orOp_69.orOp_69_in1
	// Insensitive connections
	assign orOp_69_in0 = eq_68_out;
	assign orOp_69_in1 = andOp_45_out;
	// controller for orOp_71.orOp_71_in0
	// controller for orOp_71.orOp_71_in1
	// Insensitive connections
	assign orOp_71_in0 = eq_70_out;
	assign orOp_71_in1 = andOp_30_out;
	// controller for orOp_74.orOp_74_in0
	// controller for orOp_74.orOp_74_in1
	// Insensitive connections
	assign orOp_74_in0 = eq_73_out;
	assign orOp_74_in1 = andOp_46_out;
	// controller for orOp_76.orOp_76_in0
	// controller for orOp_76.orOp_76_in1
	// Insensitive connections
	assign orOp_76_in0 = eq_75_out;
	assign orOp_76_in1 = andOp_52_out;
	// controller for orOp_78.orOp_78_in0
	// controller for orOp_78.orOp_78_in1
	// Insensitive connections
	assign orOp_78_in0 = eq_77_out;
	assign orOp_78_in1 = andOp_57_out;
	// controller for phi_phi18.phi_phi18_in
	// controller for phi_phi18.phi_phi18_last_block
	// controller for phi_phi18.phi_phi18_s
	// Insensitive connections
	assign phi_phi18_in = concat_130_out;
	assign phi_phi18_last_block = bb_1_predecessor_in_state_0_out_data;
	assign phi_phi18_s = concat_131_out;
	// controller for ret31.valid_reg
	always @(*) begin
		if (andOp_143_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// controller for sext_sext10.sext_sext10_in
	// Insensitive connections
	assign sext_sext10_in = arg_3_s_axi_arready;
	// controller for sext_sext14.sext_sext14_in
	// Insensitive connections
	assign sext_sext14_in = arg_3_s_axi_rvalid;
	// controller for sext_sext25.sext_sext25_in
	// Insensitive connections
	assign sext_sext25_in = arg_0_write_ready;
	// controller for sext_sext28.sext_sext28_in
	// Insensitive connections
	assign sext_sext28_in = data_in_1_19_out_data;
	// controller for tmp_output_111.tmp_output_111_in_data
	always @(*) begin
		if (eq_112_out) begin 
			tmp_output_111_in_data = arg_1_rdata;
		end else if (eq_115_out) begin 
			tmp_output_111_in_data = data_in_0_1_out_data;
		end else begin
			tmp_output_111_in_data = 0;
		end
	end
	// controller for tmp_output_117.tmp_output_117_in_data
	always @(*) begin
		if (eq_118_out) begin 
			tmp_output_117_in_data = arg_2_rdata;
		end else if (eq_121_out) begin 
			tmp_output_117_in_data = data_in_0_3_out_data;
		end else begin
			tmp_output_117_in_data = 0;
		end
	end
	// controller for tmp_output_135.tmp_output_135_in_data
	always @(*) begin
		if (eq_136_out) begin 
			tmp_output_135_in_data = arg_3_s_axi_rdata;
		end else if (eq_137_out) begin 
			tmp_output_135_in_data = data_in_1_15_out_data;
		end else begin
			tmp_output_135_in_data = 0;
		end
	end
	// controller for trunc_trunc30.trunc_trunc30_in
	// Insensitive connections
	assign trunc_trunc30_in = add_add29_out;
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			data_store_0_0 <= 0;
		end else begin
			if (andOp_163_out) begin
				data_store_0_0 <= arg_1_rdata;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_2 <= 0;
		end else begin
			if (andOp_164_out) begin
				data_store_0_2 <= arg_2_rdata;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_4 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_4 <= data_in_0_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_6 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_6 <= data_in_0_7_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_8 <= 0;
		end else begin
			if (andOp_165_out) begin
				data_store_0_8 <= phi_phi18_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_10 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_10 <= data_in_1_11_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_12 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_12 <= data_in_1_13_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_14 <= 0;
		end else begin
			if (andOp_168_out) begin
				data_store_1_14 <= arg_3_s_axi_rdata;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_16 <= 0;
		end else begin
			if (andOp_169_out) begin
				data_store_1_16 <= trunc_trunc30_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_18 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_18 <= data_in_1_19_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_20 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_20 <= data_in_2_21_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_22 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_22 <= data_in_2_23_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_24 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_24 <= data_in_2_25_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_26 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_26 <= data_in_2_27_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_28 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_28 <= data_in_2_29_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_145_out) begin
				global_state <= 32'd2;
			end
			if (andOp_146_out) begin
				global_state <= 32'd2;
			end
			if (andOp_36_out) begin
				global_state <= 32'd0;
			end
			if (andOp_38_out) begin
				global_state <= 32'd1;
			end
			if (andOp_43_out) begin
				global_state <= 32'd0;
			end
			if (andOp_50_out) begin
				global_state <= 32'd1;
			end
			if (andOp_55_out) begin
				global_state <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
			if (andOp_36_out) begin
				state_0_entry_BB_reg <= 32'd5;
			end
			if (andOp_43_out) begin
				state_0_entry_BB_reg <= 32'd3;
			end
			if (andOp_55_out) begin
				state_0_entry_BB_reg <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (andOp_152_out) begin
				state_0_is_active <= 1'd0;
			end
			if (andOp_36_out) begin
				state_0_is_active <= 1'd1;
			end
			if (andOp_43_out) begin
				state_0_is_active <= 1'd1;
			end
			if (andOp_55_out) begin
				state_0_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
			if (andOp_36_out) begin
				state_0_last_BB_reg <= 32'd5;
			end
			if (andOp_43_out) begin
				state_0_last_BB_reg <= 32'd3;
			end
			if (andOp_55_out) begin
				state_0_last_BB_reg <= 32'd8;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
			if (andOp_36_out) begin
				state_0_last_state <= 32'd0;
			end
			if (andOp_43_out) begin
				state_0_last_state <= 32'd0;
			end
			if (andOp_55_out) begin
				state_0_last_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_38_out) begin
				state_1_entry_BB_reg <= 32'd6;
			end
			if (andOp_50_out) begin
				state_1_entry_BB_reg <= 32'd7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_156_out) begin
				state_1_is_active <= 1'd0;
			end
			if (andOp_38_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_50_out) begin
				state_1_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_38_out) begin
				state_1_last_BB_reg <= 32'd5;
			end
			if (andOp_50_out) begin
				state_1_last_BB_reg <= 32'd7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_38_out) begin
				state_1_last_state <= 32'd0;
			end
			if (andOp_50_out) begin
				state_1_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_145_out) begin
				state_2_entry_BB_reg <= 32'd8;
			end
			if (andOp_146_out) begin
				state_2_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_145_out) begin
				state_2_is_active <= 1'd1;
			end
			if (andOp_146_out) begin
				state_2_is_active <= 1'd1;
			end
			if (andOp_160_out) begin
				state_2_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_145_out) begin
				state_2_last_BB_reg <= bb_8_predecessor_in_state_1_out_data;
			end
			if (andOp_146_out) begin
				state_2_last_BB_reg <= bb_2_predecessor_in_state_2_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_145_out) begin
				state_2_last_state <= 32'd1;
			end
			if (andOp_146_out) begin
				state_2_last_state <= 32'd2;
			end
		end
	end

endmodule

