module matrix_add(input [0:0] clk, input [0:0] rst, output [0:0] valid, output [8:0] a_debug_addr, input [31:0] a_debug_data, output [8:0] a_debug_write_addr, output [31:0] a_debug_write_data, output [0:0] a_debug_write_en, output [8:0] a_raddr_0, input [31:0] a_rdata_0, output [0:0] a_rst, output [8:0] a_waddr_0, output [31:0] a_wdata_0, output [0:0] a_wen_0, output [8:0] b_debug_addr, input [31:0] b_debug_data, output [8:0] b_debug_write_addr, output [31:0] b_debug_write_data, output [0:0] b_debug_write_en, output [8:0] b_raddr_0, input [31:0] b_rdata_0, output [0:0] b_rst, output [8:0] b_waddr_0, output [31:0] b_wdata_0, output [0:0] b_wen_0, output [8:0] c_debug_addr, input [31:0] c_debug_data, output [8:0] c_debug_write_addr, output [31:0] c_debug_write_data, output [0:0] c_debug_write_en, output [8:0] c_raddr_0, input [31:0] c_rdata_0, output [0:0] c_rst, output [8:0] c_waddr_0, output [31:0] c_wdata_0, output [0:0] c_wen_0);

	reg [0:0] valid_reg;
	reg [8:0] a_debug_addr_reg;
	reg [8:0] a_debug_write_addr_reg;
	reg [31:0] a_debug_write_data_reg;
	reg [0:0] a_debug_write_en_reg;
	reg [8:0] a_raddr_0_reg;
	reg [0:0] a_rst_reg;
	reg [8:0] a_waddr_0_reg;
	reg [31:0] a_wdata_0_reg;
	reg [0:0] a_wen_0_reg;
	reg [8:0] b_debug_addr_reg;
	reg [8:0] b_debug_write_addr_reg;
	reg [31:0] b_debug_write_data_reg;
	reg [0:0] b_debug_write_en_reg;
	reg [8:0] b_raddr_0_reg;
	reg [0:0] b_rst_reg;
	reg [8:0] b_waddr_0_reg;
	reg [31:0] b_wdata_0_reg;
	reg [0:0] b_wen_0_reg;
	reg [8:0] c_debug_addr_reg;
	reg [8:0] c_debug_write_addr_reg;
	reg [31:0] c_debug_write_data_reg;
	reg [0:0] c_debug_write_en_reg;
	reg [8:0] c_raddr_0_reg;
	reg [0:0] c_rst_reg;
	reg [8:0] c_waddr_0_reg;
	reg [31:0] c_wdata_0_reg;
	reg [0:0] c_wen_0_reg;

	assign valid = valid_reg;
	assign a_debug_addr = a_debug_addr_reg;
	assign a_debug_write_addr = a_debug_write_addr_reg;
	assign a_debug_write_data = a_debug_write_data_reg;
	assign a_debug_write_en = a_debug_write_en_reg;
	assign a_raddr_0 = a_raddr_0_reg;
	assign a_rst = a_rst_reg;
	assign a_waddr_0 = a_waddr_0_reg;
	assign a_wdata_0 = a_wdata_0_reg;
	assign a_wen_0 = a_wen_0_reg;
	assign b_debug_addr = b_debug_addr_reg;
	assign b_debug_write_addr = b_debug_write_addr_reg;
	assign b_debug_write_data = b_debug_write_data_reg;
	assign b_debug_write_en = b_debug_write_en_reg;
	assign b_raddr_0 = b_raddr_0_reg;
	assign b_rst = b_rst_reg;
	assign b_waddr_0 = b_waddr_0_reg;
	assign b_wdata_0 = b_wdata_0_reg;
	assign b_wen_0 = b_wen_0_reg;
	assign c_debug_addr = c_debug_addr_reg;
	assign c_debug_write_addr = c_debug_write_addr_reg;
	assign c_debug_write_data = c_debug_write_data_reg;
	assign c_debug_write_en = c_debug_write_en_reg;
	assign c_raddr_0 = c_raddr_0_reg;
	assign c_rst = c_rst_reg;
	assign c_waddr_0 = c_waddr_0_reg;
	assign c_wdata_0 = c_wdata_0_reg;
	assign c_wen_0 = c_wen_0_reg;

	// Start debug wires and ports

	initial begin
	end






	// End debug wires and ports

	// Start Functional Units
	br_dummy br_unit();

	wire [31:0] add_add17_in0;
	wire [31:0] add_add17_in1;
	wire [31:0] add_add17_out;
	add #(.WIDTH(32)) add_add17(.in0(add_add17_in0), .in1(add_add17_in1), .out(add_add17_out));

	wire [31:0] icmp_icmp18_in0;
	wire [31:0] icmp_icmp18_in1;
	wire [0:0] icmp_icmp18_out;
	eq #(.WIDTH(32)) icmp_icmp18(.in0(icmp_icmp18_in0), .in1(icmp_icmp18_in1), .out(icmp_icmp18_out));

	wire [63:0] phi_phi2_in;
	wire [31:0] phi_phi2_last_block;
	wire [63:0] phi_phi2_s;
	wire [31:0] phi_phi2_out;
	phi #(.DEBUG_ID(1), .NB_PAIR(2), .WIDTH(32)) phi_phi2(.in(phi_phi2_in), .last_block(phi_phi2_last_block), .out(phi_phi2_out), .s(phi_phi2_s));

	wire [31:0] add_add3_in0;
	wire [31:0] add_add3_in1;
	wire [31:0] add_add3_out;
	add #(.WIDTH(32)) add_add3(.in0(add_add3_in0), .in1(add_add3_in1), .out(add_add3_out));

	wire [31:0] add_add15_in0;
	wire [31:0] add_add15_in1;
	wire [31:0] add_add15_out;
	add #(.WIDTH(32)) add_add15(.in0(add_add15_in0), .in1(add_add15_in1), .out(add_add15_out));

	wire [31:0] add_add4_in0;
	wire [31:0] add_add4_in1;
	wire [31:0] add_add4_out;
	add #(.WIDTH(32)) add_add4(.in0(add_add4_in0), .in1(add_add4_in1), .out(add_add4_out));

	wire [31:0] icmp_icmp5_in0;
	wire [31:0] icmp_icmp5_in1;
	wire [0:0] icmp_icmp5_out;
	eq #(.WIDTH(32)) icmp_icmp5(.in0(icmp_icmp5_in0), .in1(icmp_icmp5_in1), .out(icmp_icmp5_out));

	wire [63:0] phi_phi7_in;
	wire [31:0] phi_phi7_last_block;
	wire [63:0] phi_phi7_s;
	wire [31:0] phi_phi7_out;
	phi #(.DEBUG_ID(2), .NB_PAIR(2), .WIDTH(32)) phi_phi7(.in(phi_phi7_in), .last_block(phi_phi7_last_block), .out(phi_phi7_out), .s(phi_phi7_s));

	wire [31:0] shl_shl8_in0;
	wire [31:0] shl_shl8_in1;
	wire [31:0] shl_shl8_out;
	shlOp #(.WIDTH(32)) shl_shl8(.in0(shl_shl8_in0), .in1(shl_shl8_in1), .out(shl_shl8_out));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] bb_4_active_in_state_1_in_data;
	wire [0:0] bb_4_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_1(.in_data(bb_4_active_in_state_1_in_data), .out_data(bb_4_active_in_state_1_out_data));

	reg [31:0] bb_4_predecessor_in_state_1_in_data;
	wire [31:0] bb_4_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_1(.in_data(bb_4_predecessor_in_state_1_in_data), .out_data(bb_4_predecessor_in_state_1_out_data));

	reg [0:0] br_4_happened_in_state_1_in_data;
	wire [0:0] br_4_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_1(.in_data(br_4_happened_in_state_1_in_data), .out_data(br_4_happened_in_state_1_out_data));

	reg [0:0] bb_1_active_in_state_1_in_data;
	wire [0:0] bb_1_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_1(.in_data(bb_1_active_in_state_1_in_data), .out_data(bb_1_active_in_state_1_out_data));

	reg [31:0] bb_1_predecessor_in_state_1_in_data;
	wire [31:0] bb_1_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_1(.in_data(bb_1_predecessor_in_state_1_in_data), .out_data(bb_1_predecessor_in_state_1_out_data));

	reg [0:0] br_1_happened_in_state_1_in_data;
	wire [0:0] br_1_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened_in_state_1(.in_data(br_1_happened_in_state_1_in_data), .out_data(br_1_happened_in_state_1_out_data));

	reg [0:0] bb_4_active_in_state_2_in_data;
	wire [0:0] bb_4_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_2(.in_data(bb_4_active_in_state_2_in_data), .out_data(bb_4_active_in_state_2_out_data));

	reg [31:0] bb_4_predecessor_in_state_2_in_data;
	wire [31:0] bb_4_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_2(.in_data(bb_4_predecessor_in_state_2_in_data), .out_data(bb_4_predecessor_in_state_2_out_data));

	reg [0:0] br_4_happened_in_state_2_in_data;
	wire [0:0] br_4_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_2(.in_data(br_4_happened_in_state_2_in_data), .out_data(br_4_happened_in_state_2_out_data));

	reg [0:0] bb_4_active_in_state_3_in_data;
	wire [0:0] bb_4_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_3(.in_data(bb_4_active_in_state_3_in_data), .out_data(bb_4_active_in_state_3_out_data));

	reg [31:0] bb_4_predecessor_in_state_3_in_data;
	wire [31:0] bb_4_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_3(.in_data(bb_4_predecessor_in_state_3_in_data), .out_data(bb_4_predecessor_in_state_3_out_data));

	reg [0:0] br_4_happened_in_state_3_in_data;
	wire [0:0] br_4_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_3(.in_data(br_4_happened_in_state_3_in_data), .out_data(br_4_happened_in_state_3_out_data));

	reg [0:0] bb_4_active_in_state_4_in_data;
	wire [0:0] bb_4_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_4(.in_data(bb_4_active_in_state_4_in_data), .out_data(bb_4_active_in_state_4_out_data));

	reg [31:0] bb_4_predecessor_in_state_4_in_data;
	wire [31:0] bb_4_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_4(.in_data(bb_4_predecessor_in_state_4_in_data), .out_data(bb_4_predecessor_in_state_4_out_data));

	reg [0:0] br_4_happened_in_state_4_in_data;
	wire [0:0] br_4_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_4(.in_data(br_4_happened_in_state_4_in_data), .out_data(br_4_happened_in_state_4_out_data));

	reg [0:0] bb_4_active_in_state_5_in_data;
	wire [0:0] bb_4_active_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_5(.in_data(bb_4_active_in_state_5_in_data), .out_data(bb_4_active_in_state_5_out_data));

	reg [31:0] bb_4_predecessor_in_state_5_in_data;
	wire [31:0] bb_4_predecessor_in_state_5_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_5(.in_data(bb_4_predecessor_in_state_5_in_data), .out_data(bb_4_predecessor_in_state_5_out_data));

	reg [0:0] br_4_happened_in_state_5_in_data;
	wire [0:0] br_4_happened_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_5(.in_data(br_4_happened_in_state_5_in_data), .out_data(br_4_happened_in_state_5_out_data));

	reg [0:0] bb_4_active_in_state_6_in_data;
	wire [0:0] bb_4_active_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_6(.in_data(bb_4_active_in_state_6_in_data), .out_data(bb_4_active_in_state_6_out_data));

	reg [31:0] bb_4_predecessor_in_state_6_in_data;
	wire [31:0] bb_4_predecessor_in_state_6_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_6(.in_data(bb_4_predecessor_in_state_6_in_data), .out_data(bb_4_predecessor_in_state_6_out_data));

	reg [0:0] br_4_happened_in_state_6_in_data;
	wire [0:0] br_4_happened_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_6(.in_data(br_4_happened_in_state_6_in_data), .out_data(br_4_happened_in_state_6_out_data));

	reg [0:0] bb_3_active_in_state_6_in_data;
	wire [0:0] bb_3_active_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_6(.in_data(bb_3_active_in_state_6_in_data), .out_data(bb_3_active_in_state_6_out_data));

	reg [31:0] bb_3_predecessor_in_state_6_in_data;
	wire [31:0] bb_3_predecessor_in_state_6_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_6(.in_data(bb_3_predecessor_in_state_6_in_data), .out_data(bb_3_predecessor_in_state_6_out_data));

	reg [0:0] br_3_happened_in_state_6_in_data;
	wire [0:0] br_3_happened_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_6(.in_data(br_3_happened_in_state_6_in_data), .out_data(br_3_happened_in_state_6_out_data));

	reg [0:0] bb_2_active_in_state_7_in_data;
	wire [0:0] bb_2_active_in_state_7_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_7(.in_data(bb_2_active_in_state_7_in_data), .out_data(bb_2_active_in_state_7_out_data));

	reg [31:0] bb_2_predecessor_in_state_7_in_data;
	wire [31:0] bb_2_predecessor_in_state_7_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_7(.in_data(bb_2_predecessor_in_state_7_in_data), .out_data(bb_2_predecessor_in_state_7_out_data));

	reg [31:0] data_in_0_1_in_data;
	wire [31:0] data_in_0_1_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_1(.in_data(data_in_0_1_in_data), .out_data(data_in_0_1_out_data));

	reg [31:0] data_in_0_3_in_data;
	wire [31:0] data_in_0_3_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_3(.in_data(data_in_0_3_in_data), .out_data(data_in_0_3_out_data));

	reg [31:0] data_in_0_5_in_data;
	wire [31:0] data_in_0_5_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_5(.in_data(data_in_0_5_in_data), .out_data(data_in_0_5_out_data));

	reg [31:0] data_in_0_7_in_data;
	wire [31:0] data_in_0_7_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_7(.in_data(data_in_0_7_in_data), .out_data(data_in_0_7_out_data));

	reg [31:0] data_in_1_9_in_data;
	wire [31:0] data_in_1_9_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_9(.in_data(data_in_1_9_in_data), .out_data(data_in_1_9_out_data));

	reg [31:0] data_in_1_12_in_data;
	wire [31:0] data_in_1_12_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_12(.in_data(data_in_1_12_in_data), .out_data(data_in_1_12_out_data));

	reg [31:0] data_in_1_14_in_data;
	wire [31:0] data_in_1_14_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_14(.in_data(data_in_1_14_in_data), .out_data(data_in_1_14_out_data));

	reg [31:0] data_in_1_16_in_data;
	wire [31:0] data_in_1_16_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_16(.in_data(data_in_1_16_in_data), .out_data(data_in_1_16_out_data));

	reg [31:0] data_in_2_18_in_data;
	wire [31:0] data_in_2_18_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_18(.in_data(data_in_2_18_in_data), .out_data(data_in_2_18_out_data));

	reg [31:0] data_in_2_20_in_data;
	wire [31:0] data_in_2_20_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_20(.in_data(data_in_2_20_in_data), .out_data(data_in_2_20_out_data));

	reg [31:0] data_in_2_22_in_data;
	wire [31:0] data_in_2_22_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_22(.in_data(data_in_2_22_in_data), .out_data(data_in_2_22_out_data));

	reg [31:0] data_in_2_24_in_data;
	wire [31:0] data_in_2_24_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_24(.in_data(data_in_2_24_in_data), .out_data(data_in_2_24_out_data));

	reg [31:0] data_in_2_26_in_data;
	wire [31:0] data_in_2_26_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_26(.in_data(data_in_2_26_in_data), .out_data(data_in_2_26_out_data));

	reg [31:0] data_in_3_29_in_data;
	wire [31:0] data_in_3_29_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_29(.in_data(data_in_3_29_in_data), .out_data(data_in_3_29_out_data));

	reg [31:0] data_in_3_30_in_data;
	wire [31:0] data_in_3_30_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_30(.in_data(data_in_3_30_in_data), .out_data(data_in_3_30_out_data));

	reg [31:0] data_in_3_32_in_data;
	wire [31:0] data_in_3_32_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_32(.in_data(data_in_3_32_in_data), .out_data(data_in_3_32_out_data));

	reg [31:0] data_in_3_34_in_data;
	wire [31:0] data_in_3_34_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_34(.in_data(data_in_3_34_in_data), .out_data(data_in_3_34_out_data));

	reg [31:0] data_in_3_36_in_data;
	wire [31:0] data_in_3_36_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_36(.in_data(data_in_3_36_in_data), .out_data(data_in_3_36_out_data));

	reg [31:0] data_in_3_37_in_data;
	wire [31:0] data_in_3_37_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_37(.in_data(data_in_3_37_in_data), .out_data(data_in_3_37_out_data));

	reg [31:0] data_in_4_39_in_data;
	wire [31:0] data_in_4_39_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_39(.in_data(data_in_4_39_in_data), .out_data(data_in_4_39_out_data));

	reg [31:0] data_in_4_41_in_data;
	wire [31:0] data_in_4_41_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_41(.in_data(data_in_4_41_in_data), .out_data(data_in_4_41_out_data));

	reg [31:0] data_in_4_43_in_data;
	wire [31:0] data_in_4_43_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_43(.in_data(data_in_4_43_in_data), .out_data(data_in_4_43_out_data));

	reg [31:0] data_in_4_45_in_data;
	wire [31:0] data_in_4_45_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_45(.in_data(data_in_4_45_in_data), .out_data(data_in_4_45_out_data));

	reg [31:0] data_in_5_47_in_data;
	wire [31:0] data_in_5_47_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_47(.in_data(data_in_5_47_in_data), .out_data(data_in_5_47_out_data));

	reg [31:0] data_in_5_49_in_data;
	wire [31:0] data_in_5_49_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_49(.in_data(data_in_5_49_in_data), .out_data(data_in_5_49_out_data));

	reg [31:0] data_in_5_51_in_data;
	wire [31:0] data_in_5_51_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_51(.in_data(data_in_5_51_in_data), .out_data(data_in_5_51_out_data));

	reg [31:0] data_in_5_53_in_data;
	wire [31:0] data_in_5_53_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_53(.in_data(data_in_5_53_in_data), .out_data(data_in_5_53_out_data));

	reg [31:0] data_in_6_55_in_data;
	wire [31:0] data_in_6_55_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_55(.in_data(data_in_6_55_in_data), .out_data(data_in_6_55_out_data));

	reg [31:0] data_in_6_57_in_data;
	wire [31:0] data_in_6_57_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_57(.in_data(data_in_6_57_in_data), .out_data(data_in_6_57_out_data));

	reg [31:0] data_in_6_59_in_data;
	wire [31:0] data_in_6_59_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_59(.in_data(data_in_6_59_in_data), .out_data(data_in_6_59_out_data));

	reg [31:0] data_in_6_61_in_data;
	wire [31:0] data_in_6_61_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_61(.in_data(data_in_6_61_in_data), .out_data(data_in_6_61_out_data));

	wire [0:0] andOp_62_in0;
	wire [0:0] andOp_62_in1;
	wire [0:0] andOp_62_out;
	andOp #(.WIDTH(1)) andOp_62(.in0(andOp_62_in0), .in1(andOp_62_in1), .out(andOp_62_out));

	wire [0:0] notOp_63_in0;
	wire [0:0] notOp_63_out;
	notOp #(.WIDTH(1)) notOp_63(.in(notOp_63_in0), .out(notOp_63_out));

	wire [0:0] andOp_64_in0;
	wire [0:0] andOp_64_in1;
	wire [0:0] andOp_64_out;
	andOp #(.WIDTH(1)) andOp_64(.in0(andOp_64_in0), .in1(andOp_64_in1), .out(andOp_64_out));

	wire [0:0] notOp_65_in0;
	wire [0:0] notOp_65_out;
	notOp #(.WIDTH(1)) notOp_65(.in(notOp_65_in0), .out(notOp_65_out));

	wire [0:0] andOp_66_in0;
	wire [0:0] andOp_66_in1;
	wire [0:0] andOp_66_out;
	andOp #(.WIDTH(1)) andOp_66(.in0(andOp_66_in0), .in1(andOp_66_in1), .out(andOp_66_out));

	wire [0:0] notOp_67_in0;
	wire [0:0] notOp_67_out;
	notOp #(.WIDTH(1)) notOp_67(.in(notOp_67_in0), .out(notOp_67_out));

	wire [0:0] andOp_68_in0;
	wire [0:0] andOp_68_in1;
	wire [0:0] andOp_68_out;
	andOp #(.WIDTH(1)) andOp_68(.in0(andOp_68_in0), .in1(andOp_68_in1), .out(andOp_68_out));

	wire [0:0] andOp_69_in0;
	wire [0:0] andOp_69_in1;
	wire [0:0] andOp_69_out;
	andOp #(.WIDTH(1)) andOp_69(.in0(andOp_69_in0), .in1(andOp_69_in1), .out(andOp_69_out));

	wire [0:0] notOp_70_in0;
	wire [0:0] notOp_70_out;
	notOp #(.WIDTH(1)) notOp_70(.in(notOp_70_in0), .out(notOp_70_out));

	wire [0:0] andOp_71_in0;
	wire [0:0] andOp_71_in1;
	wire [0:0] andOp_71_out;
	andOp #(.WIDTH(1)) andOp_71(.in0(andOp_71_in0), .in1(andOp_71_in1), .out(andOp_71_out));

	wire [0:0] notOp_72_in0;
	wire [0:0] notOp_72_out;
	notOp #(.WIDTH(1)) notOp_72(.in(notOp_72_in0), .out(notOp_72_out));

	wire [0:0] andOp_73_in0;
	wire [0:0] andOp_73_in1;
	wire [0:0] andOp_73_out;
	andOp #(.WIDTH(1)) andOp_73(.in0(andOp_73_in0), .in1(andOp_73_in1), .out(andOp_73_out));

	wire [0:0] notOp_74_in0;
	wire [0:0] notOp_74_out;
	notOp #(.WIDTH(1)) notOp_74(.in(notOp_74_in0), .out(notOp_74_out));

	wire [0:0] andOp_75_in0;
	wire [0:0] andOp_75_in1;
	wire [0:0] andOp_75_out;
	andOp #(.WIDTH(1)) andOp_75(.in0(andOp_75_in0), .in1(andOp_75_in1), .out(andOp_75_out));

	wire [0:0] andOp_76_in0;
	wire [0:0] andOp_76_in1;
	wire [0:0] andOp_76_out;
	andOp #(.WIDTH(1)) andOp_76(.in0(andOp_76_in0), .in1(andOp_76_in1), .out(andOp_76_out));

	wire [0:0] notOp_77_in0;
	wire [0:0] notOp_77_out;
	notOp #(.WIDTH(1)) notOp_77(.in(notOp_77_in0), .out(notOp_77_out));

	wire [0:0] andOp_78_in0;
	wire [0:0] andOp_78_in1;
	wire [0:0] andOp_78_out;
	andOp #(.WIDTH(1)) andOp_78(.in0(andOp_78_in0), .in1(andOp_78_in1), .out(andOp_78_out));

	wire [0:0] notOp_79_in0;
	wire [0:0] notOp_79_out;
	notOp #(.WIDTH(1)) notOp_79(.in(notOp_79_in0), .out(notOp_79_out));

	wire [0:0] andOp_80_in0;
	wire [0:0] andOp_80_in1;
	wire [0:0] andOp_80_out;
	andOp #(.WIDTH(1)) andOp_80(.in0(andOp_80_in0), .in1(andOp_80_in1), .out(andOp_80_out));

	wire [0:0] andOp_81_in0;
	wire [0:0] andOp_81_in1;
	wire [0:0] andOp_81_out;
	andOp #(.WIDTH(1)) andOp_81(.in0(andOp_81_in0), .in1(andOp_81_in1), .out(andOp_81_out));

	wire [0:0] notOp_82_in0;
	wire [0:0] notOp_82_out;
	notOp #(.WIDTH(1)) notOp_82(.in(notOp_82_in0), .out(notOp_82_out));

	wire [0:0] andOp_83_in0;
	wire [0:0] andOp_83_in1;
	wire [0:0] andOp_83_out;
	andOp #(.WIDTH(1)) andOp_83(.in0(andOp_83_in0), .in1(andOp_83_in1), .out(andOp_83_out));

	wire [0:0] notOp_84_in0;
	wire [0:0] notOp_84_out;
	notOp #(.WIDTH(1)) notOp_84(.in(notOp_84_in0), .out(notOp_84_out));

	wire [0:0] andOp_85_in0;
	wire [0:0] andOp_85_in1;
	wire [0:0] andOp_85_out;
	andOp #(.WIDTH(1)) andOp_85(.in0(andOp_85_in0), .in1(andOp_85_in1), .out(andOp_85_out));

	wire [0:0] andOp_86_in0;
	wire [0:0] andOp_86_in1;
	wire [0:0] andOp_86_out;
	andOp #(.WIDTH(1)) andOp_86(.in0(andOp_86_in0), .in1(andOp_86_in1), .out(andOp_86_out));

	wire [0:0] notOp_87_in0;
	wire [0:0] notOp_87_out;
	notOp #(.WIDTH(1)) notOp_87(.in(notOp_87_in0), .out(notOp_87_out));

	wire [0:0] andOp_88_in0;
	wire [0:0] andOp_88_in1;
	wire [0:0] andOp_88_out;
	andOp #(.WIDTH(1)) andOp_88(.in0(andOp_88_in0), .in1(andOp_88_in1), .out(andOp_88_out));

	wire [0:0] notOp_89_in0;
	wire [0:0] notOp_89_out;
	notOp #(.WIDTH(1)) notOp_89(.in(notOp_89_in0), .out(notOp_89_out));

	wire [0:0] andOp_90_in0;
	wire [0:0] andOp_90_in1;
	wire [0:0] andOp_90_out;
	andOp #(.WIDTH(1)) andOp_90(.in0(andOp_90_in0), .in1(andOp_90_in1), .out(andOp_90_out));

	wire [0:0] andOp_91_in0;
	wire [0:0] andOp_91_in1;
	wire [0:0] andOp_91_out;
	andOp #(.WIDTH(1)) andOp_91(.in0(andOp_91_in0), .in1(andOp_91_in1), .out(andOp_91_out));

	wire [0:0] notOp_92_in0;
	wire [0:0] notOp_92_out;
	notOp #(.WIDTH(1)) notOp_92(.in(notOp_92_in0), .out(notOp_92_out));

	wire [0:0] andOp_93_in0;
	wire [0:0] andOp_93_in1;
	wire [0:0] andOp_93_out;
	andOp #(.WIDTH(1)) andOp_93(.in0(andOp_93_in0), .in1(andOp_93_in1), .out(andOp_93_out));

	wire [0:0] notOp_94_in0;
	wire [0:0] notOp_94_out;
	notOp #(.WIDTH(1)) notOp_94(.in(notOp_94_in0), .out(notOp_94_out));

	wire [0:0] andOp_95_in0;
	wire [0:0] andOp_95_in1;
	wire [0:0] andOp_95_out;
	andOp #(.WIDTH(1)) andOp_95(.in0(andOp_95_in0), .in1(andOp_95_in1), .out(andOp_95_out));

	wire [0:0] andOp_96_in0;
	wire [0:0] andOp_96_in1;
	wire [0:0] andOp_96_out;
	andOp #(.WIDTH(1)) andOp_96(.in0(andOp_96_in0), .in1(andOp_96_in1), .out(andOp_96_out));

	wire [0:0] notOp_97_in0;
	wire [0:0] notOp_97_out;
	notOp #(.WIDTH(1)) notOp_97(.in(notOp_97_in0), .out(notOp_97_out));

	wire [0:0] andOp_98_in0;
	wire [0:0] andOp_98_in1;
	wire [0:0] andOp_98_out;
	andOp #(.WIDTH(1)) andOp_98(.in0(andOp_98_in0), .in1(andOp_98_in1), .out(andOp_98_out));

	wire [0:0] notOp_99_in0;
	wire [0:0] notOp_99_out;
	notOp #(.WIDTH(1)) notOp_99(.in(notOp_99_in0), .out(notOp_99_out));

	wire [0:0] andOp_100_in0;
	wire [0:0] andOp_100_in1;
	wire [0:0] andOp_100_out;
	andOp #(.WIDTH(1)) andOp_100(.in0(andOp_100_in0), .in1(andOp_100_in1), .out(andOp_100_out));

	wire [31:0] eq_101_in0;
	wire [31:0] eq_101_in1;
	wire [0:0] eq_101_out;
	eq #(.WIDTH(32)) eq_101(.in0(eq_101_in0), .in1(eq_101_in1), .out(eq_101_out));

	wire [31:0] eq_102_in0;
	wire [31:0] eq_102_in1;
	wire [0:0] eq_102_out;
	eq #(.WIDTH(32)) eq_102(.in0(eq_102_in0), .in1(eq_102_in1), .out(eq_102_out));

	wire [0:0] orOp_103_in0;
	wire [0:0] orOp_103_in1;
	wire [0:0] orOp_103_out;
	orOp #(.WIDTH(1)) orOp_103(.in0(orOp_103_in0), .in1(orOp_103_in1), .out(orOp_103_out));

	wire [31:0] eq_104_in0;
	wire [31:0] eq_104_in1;
	wire [0:0] eq_104_out;
	eq #(.WIDTH(32)) eq_104(.in0(eq_104_in0), .in1(eq_104_in1), .out(eq_104_out));

	wire [31:0] eq_105_in0;
	wire [31:0] eq_105_in1;
	wire [0:0] eq_105_out;
	eq #(.WIDTH(32)) eq_105(.in0(eq_105_in0), .in1(eq_105_in1), .out(eq_105_out));

	wire [31:0] eq_106_in0;
	wire [31:0] eq_106_in1;
	wire [0:0] eq_106_out;
	eq #(.WIDTH(32)) eq_106(.in0(eq_106_in0), .in1(eq_106_in1), .out(eq_106_out));

	wire [31:0] eq_107_in0;
	wire [31:0] eq_107_in1;
	wire [0:0] eq_107_out;
	eq #(.WIDTH(32)) eq_107(.in0(eq_107_in0), .in1(eq_107_in1), .out(eq_107_out));

	wire [31:0] eq_108_in0;
	wire [31:0] eq_108_in1;
	wire [0:0] eq_108_out;
	eq #(.WIDTH(32)) eq_108(.in0(eq_108_in0), .in1(eq_108_in1), .out(eq_108_out));

	wire [31:0] eq_109_in0;
	wire [31:0] eq_109_in1;
	wire [0:0] eq_109_out;
	eq #(.WIDTH(32)) eq_109(.in0(eq_109_in0), .in1(eq_109_in1), .out(eq_109_out));

	wire [31:0] eq_110_in0;
	wire [31:0] eq_110_in1;
	wire [0:0] eq_110_out;
	eq #(.WIDTH(32)) eq_110(.in0(eq_110_in0), .in1(eq_110_in1), .out(eq_110_out));

	wire [0:0] orOp_111_in0;
	wire [0:0] orOp_111_in1;
	wire [0:0] orOp_111_out;
	orOp #(.WIDTH(1)) orOp_111(.in0(orOp_111_in0), .in1(orOp_111_in1), .out(orOp_111_out));

	wire [31:0] eq_112_in0;
	wire [31:0] eq_112_in1;
	wire [0:0] eq_112_out;
	eq #(.WIDTH(32)) eq_112(.in0(eq_112_in0), .in1(eq_112_in1), .out(eq_112_out));

	wire [31:0] eq_113_in0;
	wire [31:0] eq_113_in1;
	wire [0:0] eq_113_out;
	eq #(.WIDTH(32)) eq_113(.in0(eq_113_in0), .in1(eq_113_in1), .out(eq_113_out));

	wire [31:0] eq_114_in0;
	wire [31:0] eq_114_in1;
	wire [0:0] eq_114_out;
	eq #(.WIDTH(32)) eq_114(.in0(eq_114_in0), .in1(eq_114_in1), .out(eq_114_out));

	wire [0:0] notOp_115_in0;
	wire [0:0] notOp_115_out;
	notOp #(.WIDTH(1)) notOp_115(.in(notOp_115_in0), .out(notOp_115_out));

	wire [0:0] andOp_116_in0;
	wire [0:0] andOp_116_in1;
	wire [0:0] andOp_116_out;
	andOp #(.WIDTH(1)) andOp_116(.in0(andOp_116_in0), .in1(andOp_116_in1), .out(andOp_116_out));

	wire [31:0] eq_117_in0;
	wire [31:0] eq_117_in1;
	wire [0:0] eq_117_out;
	eq #(.WIDTH(32)) eq_117(.in0(eq_117_in0), .in1(eq_117_in1), .out(eq_117_out));

	wire [31:0] eq_118_in0;
	wire [31:0] eq_118_in1;
	wire [0:0] eq_118_out;
	eq #(.WIDTH(32)) eq_118(.in0(eq_118_in0), .in1(eq_118_in1), .out(eq_118_out));

	wire [31:0] eq_119_in0;
	wire [31:0] eq_119_in1;
	wire [0:0] eq_119_out;
	eq #(.WIDTH(32)) eq_119(.in0(eq_119_in0), .in1(eq_119_in1), .out(eq_119_out));

	wire [31:0] eq_120_in0;
	wire [31:0] eq_120_in1;
	wire [0:0] eq_120_out;
	eq #(.WIDTH(32)) eq_120(.in0(eq_120_in0), .in1(eq_120_in1), .out(eq_120_out));

	wire [31:0] eq_121_in0;
	wire [31:0] eq_121_in1;
	wire [0:0] eq_121_out;
	eq #(.WIDTH(32)) eq_121(.in0(eq_121_in0), .in1(eq_121_in1), .out(eq_121_out));

	wire [31:0] eq_122_in0;
	wire [31:0] eq_122_in1;
	wire [0:0] eq_122_out;
	eq #(.WIDTH(32)) eq_122(.in0(eq_122_in0), .in1(eq_122_in1), .out(eq_122_out));

	wire [31:0] eq_123_in0;
	wire [31:0] eq_123_in1;
	wire [0:0] eq_123_out;
	eq #(.WIDTH(32)) eq_123(.in0(eq_123_in0), .in1(eq_123_in1), .out(eq_123_out));

	wire [0:0] notOp_124_in0;
	wire [0:0] notOp_124_out;
	notOp #(.WIDTH(1)) notOp_124(.in(notOp_124_in0), .out(notOp_124_out));

	wire [0:0] andOp_125_in0;
	wire [0:0] andOp_125_in1;
	wire [0:0] andOp_125_out;
	andOp #(.WIDTH(1)) andOp_125(.in0(andOp_125_in0), .in1(andOp_125_in1), .out(andOp_125_out));

	wire [31:0] eq_126_in0;
	wire [31:0] eq_126_in1;
	wire [0:0] eq_126_out;
	eq #(.WIDTH(32)) eq_126(.in0(eq_126_in0), .in1(eq_126_in1), .out(eq_126_out));

	wire [0:0] andOp_127_in0;
	wire [0:0] andOp_127_in1;
	wire [0:0] andOp_127_out;
	andOp #(.WIDTH(1)) andOp_127(.in0(andOp_127_in0), .in1(andOp_127_in1), .out(andOp_127_out));

	wire [31:0] concat_128_in0;
	wire [31:0] concat_128_in1;
	wire [63:0] concat_128_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_128(.in0(concat_128_in0), .in1(concat_128_in1), .out(concat_128_out));

	wire [31:0] concat_129_in0;
	wire [31:0] concat_129_in1;
	wire [63:0] concat_129_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_129(.in0(concat_129_in0), .in1(concat_129_in1), .out(concat_129_out));

	wire [0:0] andOp_130_in0;
	wire [0:0] andOp_130_in1;
	wire [0:0] andOp_130_out;
	andOp #(.WIDTH(1)) andOp_130(.in0(andOp_130_in0), .in1(andOp_130_in1), .out(andOp_130_out));

	reg [31:0] tmp_output_131_in_data;
	wire [31:0] tmp_output_131_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_131(.in_data(tmp_output_131_in_data), .out_data(tmp_output_131_out_data));

	wire [31:0] eq_132_in0;
	wire [31:0] eq_132_in1;
	wire [0:0] eq_132_out;
	eq #(.WIDTH(32)) eq_132(.in0(eq_132_in0), .in1(eq_132_in1), .out(eq_132_out));

	wire [31:0] eq_133_in0;
	wire [31:0] eq_133_in1;
	wire [0:0] eq_133_out;
	eq #(.WIDTH(32)) eq_133(.in0(eq_133_in0), .in1(eq_133_in1), .out(eq_133_out));

	wire [0:0] andOp_134_in0;
	wire [0:0] andOp_134_in1;
	wire [0:0] andOp_134_out;
	andOp #(.WIDTH(1)) andOp_134(.in0(andOp_134_in0), .in1(andOp_134_in1), .out(andOp_134_out));

	wire [0:0] andOp_135_in0;
	wire [0:0] andOp_135_in1;
	wire [0:0] andOp_135_out;
	andOp #(.WIDTH(1)) andOp_135(.in0(andOp_135_in0), .in1(andOp_135_in1), .out(andOp_135_out));

	wire [0:0] andOp_136_in0;
	wire [0:0] andOp_136_in1;
	wire [0:0] andOp_136_out;
	andOp #(.WIDTH(1)) andOp_136(.in0(andOp_136_in0), .in1(andOp_136_in1), .out(andOp_136_out));

	wire [31:0] concat_137_in0;
	wire [31:0] concat_137_in1;
	wire [63:0] concat_137_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_137(.in0(concat_137_in0), .in1(concat_137_in1), .out(concat_137_out));

	wire [31:0] concat_138_in0;
	wire [31:0] concat_138_in1;
	wire [63:0] concat_138_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_138(.in0(concat_138_in0), .in1(concat_138_in1), .out(concat_138_out));

	wire [0:0] andOp_139_in0;
	wire [0:0] andOp_139_in1;
	wire [0:0] andOp_139_out;
	andOp #(.WIDTH(1)) andOp_139(.in0(andOp_139_in0), .in1(andOp_139_in1), .out(andOp_139_out));

	wire [0:0] andOp_140_in0;
	wire [0:0] andOp_140_in1;
	wire [0:0] andOp_140_out;
	andOp #(.WIDTH(1)) andOp_140(.in0(andOp_140_in0), .in1(andOp_140_in1), .out(andOp_140_out));

	wire [0:0] andOp_141_in0;
	wire [0:0] andOp_141_in1;
	wire [0:0] andOp_141_out;
	andOp #(.WIDTH(1)) andOp_141(.in0(andOp_141_in0), .in1(andOp_141_in1), .out(andOp_141_out));

	wire [0:0] andOp_142_in0;
	wire [0:0] andOp_142_in1;
	wire [0:0] andOp_142_out;
	andOp #(.WIDTH(1)) andOp_142(.in0(andOp_142_in0), .in1(andOp_142_in1), .out(andOp_142_out));

	wire [0:0] andOp_143_in0;
	wire [0:0] andOp_143_in1;
	wire [0:0] andOp_143_out;
	andOp #(.WIDTH(1)) andOp_143(.in0(andOp_143_in0), .in1(andOp_143_in1), .out(andOp_143_out));

	wire [0:0] andOp_144_in0;
	wire [0:0] andOp_144_in1;
	wire [0:0] andOp_144_out;
	andOp #(.WIDTH(1)) andOp_144(.in0(andOp_144_in0), .in1(andOp_144_in1), .out(andOp_144_out));

	wire [0:0] andOp_145_in0;
	wire [0:0] andOp_145_in1;
	wire [0:0] andOp_145_out;
	andOp #(.WIDTH(1)) andOp_145(.in0(andOp_145_in0), .in1(andOp_145_in1), .out(andOp_145_out));

	wire [0:0] andOp_146_in0;
	wire [0:0] andOp_146_in1;
	wire [0:0] andOp_146_out;
	andOp #(.WIDTH(1)) andOp_146(.in0(andOp_146_in0), .in1(andOp_146_in1), .out(andOp_146_out));

	wire [0:0] andOp_147_in0;
	wire [0:0] andOp_147_in1;
	wire [0:0] andOp_147_out;
	andOp #(.WIDTH(1)) andOp_147(.in0(andOp_147_in0), .in1(andOp_147_in1), .out(andOp_147_out));

	wire [0:0] andOp_148_in0;
	wire [0:0] andOp_148_in1;
	wire [0:0] andOp_148_out;
	andOp #(.WIDTH(1)) andOp_148(.in0(andOp_148_in0), .in1(andOp_148_in1), .out(andOp_148_out));

	wire [0:0] andOp_149_in0;
	wire [0:0] andOp_149_in1;
	wire [0:0] andOp_149_out;
	andOp #(.WIDTH(1)) andOp_149(.in0(andOp_149_in0), .in1(andOp_149_in1), .out(andOp_149_out));

	wire [0:0] andOp_150_in0;
	wire [0:0] andOp_150_in1;
	wire [0:0] andOp_150_out;
	andOp #(.WIDTH(1)) andOp_150(.in0(andOp_150_in0), .in1(andOp_150_in1), .out(andOp_150_out));

	wire [0:0] andOp_151_in0;
	wire [0:0] andOp_151_in1;
	wire [0:0] andOp_151_out;
	andOp #(.WIDTH(1)) andOp_151(.in0(andOp_151_in0), .in1(andOp_151_in1), .out(andOp_151_out));

	wire [0:0] andOp_152_in0;
	wire [0:0] andOp_152_in1;
	wire [0:0] andOp_152_out;
	andOp #(.WIDTH(1)) andOp_152(.in0(andOp_152_in0), .in1(andOp_152_in1), .out(andOp_152_out));

	wire [0:0] andOp_153_in0;
	wire [0:0] andOp_153_in1;
	wire [0:0] andOp_153_out;
	andOp #(.WIDTH(1)) andOp_153(.in0(andOp_153_in0), .in1(andOp_153_in1), .out(andOp_153_out));

	wire [0:0] andOp_154_in0;
	wire [0:0] andOp_154_in1;
	wire [0:0] andOp_154_out;
	andOp #(.WIDTH(1)) andOp_154(.in0(andOp_154_in0), .in1(andOp_154_in1), .out(andOp_154_out));

	wire [0:0] andOp_155_in0;
	wire [0:0] andOp_155_in1;
	wire [0:0] andOp_155_out;
	andOp #(.WIDTH(1)) andOp_155(.in0(andOp_155_in0), .in1(andOp_155_in1), .out(andOp_155_out));

	wire [0:0] notOp_156_in0;
	wire [0:0] notOp_156_out;
	notOp #(.WIDTH(1)) notOp_156(.in(notOp_156_in0), .out(notOp_156_out));

	wire [0:0] andOp_157_in0;
	wire [0:0] andOp_157_in1;
	wire [0:0] andOp_157_out;
	andOp #(.WIDTH(1)) andOp_157(.in0(andOp_157_in0), .in1(andOp_157_in1), .out(andOp_157_out));

	wire [0:0] notOp_158_in0;
	wire [0:0] notOp_158_out;
	notOp #(.WIDTH(1)) notOp_158(.in(notOp_158_in0), .out(notOp_158_out));

	wire [0:0] andOp_159_in0;
	wire [0:0] andOp_159_in1;
	wire [0:0] andOp_159_out;
	andOp #(.WIDTH(1)) andOp_159(.in0(andOp_159_in0), .in1(andOp_159_in1), .out(andOp_159_out));

	wire [0:0] notOp_160_in0;
	wire [0:0] notOp_160_out;
	notOp #(.WIDTH(1)) notOp_160(.in(notOp_160_in0), .out(notOp_160_out));

	wire [0:0] andOp_161_in0;
	wire [0:0] andOp_161_in1;
	wire [0:0] andOp_161_out;
	andOp #(.WIDTH(1)) andOp_161(.in0(andOp_161_in0), .in1(andOp_161_in1), .out(andOp_161_out));

	wire [0:0] notOp_162_in0;
	wire [0:0] notOp_162_out;
	notOp #(.WIDTH(1)) notOp_162(.in(notOp_162_in0), .out(notOp_162_out));

	wire [0:0] andOp_163_in0;
	wire [0:0] andOp_163_in1;
	wire [0:0] andOp_163_out;
	andOp #(.WIDTH(1)) andOp_163(.in0(andOp_163_in0), .in1(andOp_163_in1), .out(andOp_163_out));

	wire [0:0] notOp_164_in0;
	wire [0:0] notOp_164_out;
	notOp #(.WIDTH(1)) notOp_164(.in(notOp_164_in0), .out(notOp_164_out));

	wire [0:0] andOp_165_in0;
	wire [0:0] andOp_165_in1;
	wire [0:0] andOp_165_out;
	andOp #(.WIDTH(1)) andOp_165(.in0(andOp_165_in0), .in1(andOp_165_in1), .out(andOp_165_out));

	wire [0:0] andOp_166_in0;
	wire [0:0] andOp_166_in1;
	wire [0:0] andOp_166_out;
	andOp #(.WIDTH(1)) andOp_166(.in0(andOp_166_in0), .in1(andOp_166_in1), .out(andOp_166_out));

	wire [0:0] andOp_167_in0;
	wire [0:0] andOp_167_in1;
	wire [0:0] andOp_167_out;
	andOp #(.WIDTH(1)) andOp_167(.in0(andOp_167_in0), .in1(andOp_167_in1), .out(andOp_167_out));

	wire [0:0] andOp_168_in0;
	wire [0:0] andOp_168_in1;
	wire [0:0] andOp_168_out;
	andOp #(.WIDTH(1)) andOp_168(.in0(andOp_168_in0), .in1(andOp_168_in1), .out(andOp_168_out));

	wire [0:0] notOp_169_in0;
	wire [0:0] notOp_169_out;
	notOp #(.WIDTH(1)) notOp_169(.in(notOp_169_in0), .out(notOp_169_out));

	wire [0:0] andOp_170_in0;
	wire [0:0] andOp_170_in1;
	wire [0:0] andOp_170_out;
	andOp #(.WIDTH(1)) andOp_170(.in0(andOp_170_in0), .in1(andOp_170_in1), .out(andOp_170_out));

	wire [0:0] notOp_171_in0;
	wire [0:0] notOp_171_out;
	notOp #(.WIDTH(1)) notOp_171(.in(notOp_171_in0), .out(notOp_171_out));

	wire [0:0] andOp_172_in0;
	wire [0:0] andOp_172_in1;
	wire [0:0] andOp_172_out;
	andOp #(.WIDTH(1)) andOp_172(.in0(andOp_172_in0), .in1(andOp_172_in1), .out(andOp_172_out));

	wire [0:0] notOp_173_in0;
	wire [0:0] notOp_173_out;
	notOp #(.WIDTH(1)) notOp_173(.in(notOp_173_in0), .out(notOp_173_out));

	wire [0:0] andOp_174_in0;
	wire [0:0] andOp_174_in1;
	wire [0:0] andOp_174_out;
	andOp #(.WIDTH(1)) andOp_174(.in0(andOp_174_in0), .in1(andOp_174_in1), .out(andOp_174_out));

	wire [0:0] notOp_175_in0;
	wire [0:0] notOp_175_out;
	notOp #(.WIDTH(1)) notOp_175(.in(notOp_175_in0), .out(notOp_175_out));

	wire [0:0] andOp_176_in0;
	wire [0:0] andOp_176_in1;
	wire [0:0] andOp_176_out;
	andOp #(.WIDTH(1)) andOp_176(.in0(andOp_176_in0), .in1(andOp_176_in1), .out(andOp_176_out));

	wire [0:0] notOp_177_in0;
	wire [0:0] notOp_177_out;
	notOp #(.WIDTH(1)) notOp_177(.in(notOp_177_in0), .out(notOp_177_out));

	wire [0:0] andOp_178_in0;
	wire [0:0] andOp_178_in1;
	wire [0:0] andOp_178_out;
	andOp #(.WIDTH(1)) andOp_178(.in0(andOp_178_in0), .in1(andOp_178_in1), .out(andOp_178_out));

	wire [0:0] andOp_179_in0;
	wire [0:0] andOp_179_in1;
	wire [0:0] andOp_179_out;
	andOp #(.WIDTH(1)) andOp_179(.in0(andOp_179_in0), .in1(andOp_179_in1), .out(andOp_179_out));

	wire [0:0] andOp_180_in0;
	wire [0:0] andOp_180_in1;
	wire [0:0] andOp_180_out;
	andOp #(.WIDTH(1)) andOp_180(.in0(andOp_180_in0), .in1(andOp_180_in1), .out(andOp_180_out));

	wire [0:0] andOp_181_in0;
	wire [0:0] andOp_181_in1;
	wire [0:0] andOp_181_out;
	andOp #(.WIDTH(1)) andOp_181(.in0(andOp_181_in0), .in1(andOp_181_in1), .out(andOp_181_out));

	wire [0:0] notOp_182_in0;
	wire [0:0] notOp_182_out;
	notOp #(.WIDTH(1)) notOp_182(.in(notOp_182_in0), .out(notOp_182_out));

	wire [0:0] andOp_183_in0;
	wire [0:0] andOp_183_in1;
	wire [0:0] andOp_183_out;
	andOp #(.WIDTH(1)) andOp_183(.in0(andOp_183_in0), .in1(andOp_183_in1), .out(andOp_183_out));

	wire [0:0] notOp_184_in0;
	wire [0:0] notOp_184_out;
	notOp #(.WIDTH(1)) notOp_184(.in(notOp_184_in0), .out(notOp_184_out));

	wire [0:0] andOp_185_in0;
	wire [0:0] andOp_185_in1;
	wire [0:0] andOp_185_out;
	andOp #(.WIDTH(1)) andOp_185(.in0(andOp_185_in0), .in1(andOp_185_in1), .out(andOp_185_out));

	wire [0:0] notOp_186_in0;
	wire [0:0] notOp_186_out;
	notOp #(.WIDTH(1)) notOp_186(.in(notOp_186_in0), .out(notOp_186_out));

	wire [0:0] andOp_187_in0;
	wire [0:0] andOp_187_in1;
	wire [0:0] andOp_187_out;
	andOp #(.WIDTH(1)) andOp_187(.in0(andOp_187_in0), .in1(andOp_187_in1), .out(andOp_187_out));

	wire [0:0] notOp_188_in0;
	wire [0:0] notOp_188_out;
	notOp #(.WIDTH(1)) notOp_188(.in(notOp_188_in0), .out(notOp_188_out));

	wire [0:0] andOp_189_in0;
	wire [0:0] andOp_189_in1;
	wire [0:0] andOp_189_out;
	andOp #(.WIDTH(1)) andOp_189(.in0(andOp_189_in0), .in1(andOp_189_in1), .out(andOp_189_out));

	wire [0:0] notOp_190_in0;
	wire [0:0] notOp_190_out;
	notOp #(.WIDTH(1)) notOp_190(.in(notOp_190_in0), .out(notOp_190_out));

	wire [0:0] andOp_191_in0;
	wire [0:0] andOp_191_in1;
	wire [0:0] andOp_191_out;
	andOp #(.WIDTH(1)) andOp_191(.in0(andOp_191_in0), .in1(andOp_191_in1), .out(andOp_191_out));

	wire [0:0] notOp_192_in0;
	wire [0:0] notOp_192_out;
	notOp #(.WIDTH(1)) notOp_192(.in(notOp_192_in0), .out(notOp_192_out));

	wire [0:0] andOp_193_in0;
	wire [0:0] andOp_193_in1;
	wire [0:0] andOp_193_out;
	andOp #(.WIDTH(1)) andOp_193(.in0(andOp_193_in0), .in1(andOp_193_in1), .out(andOp_193_out));

	wire [0:0] notOp_194_in0;
	wire [0:0] notOp_194_out;
	notOp #(.WIDTH(1)) notOp_194(.in(notOp_194_in0), .out(notOp_194_out));

	wire [0:0] andOp_195_in0;
	wire [0:0] andOp_195_in1;
	wire [0:0] andOp_195_out;
	andOp #(.WIDTH(1)) andOp_195(.in0(andOp_195_in0), .in1(andOp_195_in1), .out(andOp_195_out));

	wire [0:0] notOp_196_in0;
	wire [0:0] notOp_196_out;
	notOp #(.WIDTH(1)) notOp_196(.in(notOp_196_in0), .out(notOp_196_out));

	wire [0:0] andOp_197_in0;
	wire [0:0] andOp_197_in1;
	wire [0:0] andOp_197_out;
	andOp #(.WIDTH(1)) andOp_197(.in0(andOp_197_in0), .in1(andOp_197_in1), .out(andOp_197_out));

	wire [0:0] notOp_198_in0;
	wire [0:0] notOp_198_out;
	notOp #(.WIDTH(1)) notOp_198(.in(notOp_198_in0), .out(notOp_198_out));

	wire [0:0] andOp_199_in0;
	wire [0:0] andOp_199_in1;
	wire [0:0] andOp_199_out;
	andOp #(.WIDTH(1)) andOp_199(.in0(andOp_199_in0), .in1(andOp_199_in1), .out(andOp_199_out));

	wire [0:0] notOp_200_in0;
	wire [0:0] notOp_200_out;
	notOp #(.WIDTH(1)) notOp_200(.in(notOp_200_in0), .out(notOp_200_out));

	wire [0:0] andOp_201_in0;
	wire [0:0] andOp_201_in1;
	wire [0:0] andOp_201_out;
	andOp #(.WIDTH(1)) andOp_201(.in0(andOp_201_in0), .in1(andOp_201_in1), .out(andOp_201_out));

	wire [0:0] notOp_202_in0;
	wire [0:0] notOp_202_out;
	notOp #(.WIDTH(1)) notOp_202(.in(notOp_202_in0), .out(notOp_202_out));

	wire [0:0] andOp_203_in0;
	wire [0:0] andOp_203_in1;
	wire [0:0] andOp_203_out;
	andOp #(.WIDTH(1)) andOp_203(.in0(andOp_203_in0), .in1(andOp_203_in1), .out(andOp_203_out));

	reg [0:0] in_pipeline_0_in_data;
	wire [0:0] in_pipeline_0_out_data;
	hls_wire #(.WIDTH(1)) in_pipeline_0(.in_data(in_pipeline_0_in_data), .out_data(in_pipeline_0_out_data));

	wire [0:0] orOp_204_in0;
	wire [0:0] orOp_204_in1;
	wire [0:0] orOp_204_out;
	orOp #(.WIDTH(1)) orOp_204(.in0(orOp_204_in0), .in1(orOp_204_in1), .out(orOp_204_out));

	wire [0:0] orOp_205_in0;
	wire [0:0] orOp_205_in1;
	wire [0:0] orOp_205_out;
	orOp #(.WIDTH(1)) orOp_205(.in0(orOp_205_in0), .in1(orOp_205_in1), .out(orOp_205_out));

	wire [0:0] orOp_206_in0;
	wire [0:0] orOp_206_in1;
	wire [0:0] orOp_206_out;
	orOp #(.WIDTH(1)) orOp_206(.in0(orOp_206_in0), .in1(orOp_206_in1), .out(orOp_206_out));

	wire [0:0] orOp_207_in0;
	wire [0:0] orOp_207_in1;
	wire [0:0] orOp_207_out;
	orOp #(.WIDTH(1)) orOp_207(.in0(orOp_207_in0), .in1(orOp_207_in1), .out(orOp_207_out));

	wire [0:0] orOp_208_in0;
	wire [0:0] orOp_208_in1;
	wire [0:0] orOp_208_out;
	orOp #(.WIDTH(1)) orOp_208(.in0(orOp_208_in0), .in1(orOp_208_in1), .out(orOp_208_out));

	wire [0:0] orOp_209_in0;
	wire [0:0] orOp_209_in1;
	wire [0:0] orOp_209_out;
	orOp #(.WIDTH(1)) orOp_209(.in0(orOp_209_in0), .in1(orOp_209_in1), .out(orOp_209_out));

	wire [31:0] eq_210_in0;
	wire [31:0] eq_210_in1;
	wire [0:0] eq_210_out;
	eq #(.WIDTH(32)) eq_210(.in0(eq_210_in0), .in1(eq_210_in1), .out(eq_210_out));

	wire [31:0] eq_211_in0;
	wire [31:0] eq_211_in1;
	wire [0:0] eq_211_out;
	eq #(.WIDTH(32)) eq_211(.in0(eq_211_in0), .in1(eq_211_in1), .out(eq_211_out));

	wire [31:0] eq_212_in0;
	wire [31:0] eq_212_in1;
	wire [0:0] eq_212_out;
	eq #(.WIDTH(32)) eq_212(.in0(eq_212_in0), .in1(eq_212_in1), .out(eq_212_out));

	wire [31:0] eq_213_in0;
	wire [31:0] eq_213_in1;
	wire [0:0] eq_213_out;
	eq #(.WIDTH(32)) eq_213(.in0(eq_213_in0), .in1(eq_213_in1), .out(eq_213_out));

	wire [0:0] andOp_214_in0;
	wire [0:0] andOp_214_in1;
	wire [0:0] andOp_214_out;
	andOp #(.WIDTH(1)) andOp_214(.in0(andOp_214_in0), .in1(andOp_214_in1), .out(andOp_214_out));

	wire [0:0] andOp_215_in0;
	wire [0:0] andOp_215_in1;
	wire [0:0] andOp_215_out;
	andOp #(.WIDTH(1)) andOp_215(.in0(andOp_215_in0), .in1(andOp_215_in1), .out(andOp_215_out));

	wire [0:0] andOp_216_in0;
	wire [0:0] andOp_216_in1;
	wire [0:0] andOp_216_out;
	andOp #(.WIDTH(1)) andOp_216(.in0(andOp_216_in0), .in1(andOp_216_in1), .out(andOp_216_out));

	wire [0:0] andOp_217_in0;
	wire [0:0] andOp_217_in1;
	wire [0:0] andOp_217_out;
	andOp #(.WIDTH(1)) andOp_217(.in0(andOp_217_in0), .in1(andOp_217_in1), .out(andOp_217_out));

	wire [31:0] eq_218_in0;
	wire [31:0] eq_218_in1;
	wire [0:0] eq_218_out;
	eq #(.WIDTH(32)) eq_218(.in0(eq_218_in0), .in1(eq_218_in1), .out(eq_218_out));

	wire [31:0] eq_219_in0;
	wire [31:0] eq_219_in1;
	wire [0:0] eq_219_out;
	eq #(.WIDTH(32)) eq_219(.in0(eq_219_in0), .in1(eq_219_in1), .out(eq_219_out));

	wire [0:0] andOp_220_in0;
	wire [0:0] andOp_220_in1;
	wire [0:0] andOp_220_out;
	andOp #(.WIDTH(1)) andOp_220(.in0(andOp_220_in0), .in1(andOp_220_in1), .out(andOp_220_out));

	wire [31:0] eq_221_in0;
	wire [31:0] eq_221_in1;
	wire [0:0] eq_221_out;
	eq #(.WIDTH(32)) eq_221(.in0(eq_221_in0), .in1(eq_221_in1), .out(eq_221_out));

	wire [31:0] eq_222_in0;
	wire [31:0] eq_222_in1;
	wire [0:0] eq_222_out;
	eq #(.WIDTH(32)) eq_222(.in0(eq_222_in0), .in1(eq_222_in1), .out(eq_222_out));

	wire [31:0] eq_223_in0;
	wire [31:0] eq_223_in1;
	wire [0:0] eq_223_out;
	eq #(.WIDTH(32)) eq_223(.in0(eq_223_in0), .in1(eq_223_in1), .out(eq_223_out));

	wire [31:0] eq_224_in0;
	wire [31:0] eq_224_in1;
	wire [0:0] eq_224_out;
	eq #(.WIDTH(32)) eq_224(.in0(eq_224_in0), .in1(eq_224_in1), .out(eq_224_out));

	wire [31:0] eq_225_in0;
	wire [31:0] eq_225_in1;
	wire [0:0] eq_225_out;
	eq #(.WIDTH(32)) eq_225(.in0(eq_225_in0), .in1(eq_225_in1), .out(eq_225_out));

	wire [31:0] eq_226_in0;
	wire [31:0] eq_226_in1;
	wire [0:0] eq_226_out;
	eq #(.WIDTH(32)) eq_226(.in0(eq_226_in0), .in1(eq_226_in1), .out(eq_226_out));

	wire [31:0] eq_227_in0;
	wire [31:0] eq_227_in1;
	wire [0:0] eq_227_out;
	eq #(.WIDTH(32)) eq_227(.in0(eq_227_in0), .in1(eq_227_in1), .out(eq_227_out));

	wire [31:0] eq_228_in0;
	wire [31:0] eq_228_in1;
	wire [0:0] eq_228_out;
	eq #(.WIDTH(32)) eq_228(.in0(eq_228_in0), .in1(eq_228_in1), .out(eq_228_out));

	wire [31:0] eq_229_in0;
	wire [31:0] eq_229_in1;
	wire [0:0] eq_229_out;
	eq #(.WIDTH(32)) eq_229(.in0(eq_229_in0), .in1(eq_229_in1), .out(eq_229_out));

	wire [0:0] andOp_230_in0;
	wire [0:0] andOp_230_in1;
	wire [0:0] andOp_230_out;
	andOp #(.WIDTH(1)) andOp_230(.in0(andOp_230_in0), .in1(andOp_230_in1), .out(andOp_230_out));

	wire [31:0] eq_231_in0;
	wire [31:0] eq_231_in1;
	wire [0:0] eq_231_out;
	eq #(.WIDTH(32)) eq_231(.in0(eq_231_in0), .in1(eq_231_in1), .out(eq_231_out));

	wire [31:0] eq_232_in0;
	wire [31:0] eq_232_in1;
	wire [0:0] eq_232_out;
	eq #(.WIDTH(32)) eq_232(.in0(eq_232_in0), .in1(eq_232_in1), .out(eq_232_out));

	// End Functional Units

	reg [31:0] data_store_0_0;
	reg [31:0] data_store_0_2;
	reg [31:0] data_store_0_4;
	reg [31:0] data_store_0_6;
	reg [31:0] data_store_1_10;
	reg [31:0] data_store_1_11;
	reg [31:0] data_store_1_13;
	reg [31:0] data_store_1_15;
	reg [31:0] data_store_1_8;
	reg [31:0] data_store_2_17;
	reg [31:0] data_store_2_19;
	reg [31:0] data_store_2_21;
	reg [31:0] data_store_2_23;
	reg [31:0] data_store_2_25;
	reg [31:0] data_store_2_27;
	reg [31:0] data_store_3_28;
	reg [31:0] data_store_3_31;
	reg [31:0] data_store_3_33;
	reg [31:0] data_store_3_35;
	reg [31:0] data_store_4_38;
	reg [31:0] data_store_4_40;
	reg [31:0] data_store_4_42;
	reg [31:0] data_store_4_44;
	reg [31:0] data_store_5_46;
	reg [31:0] data_store_5_48;
	reg [31:0] data_store_5_50;
	reg [31:0] data_store_5_52;
	reg [31:0] data_store_6_54;
	reg [31:0] data_store_6_56;
	reg [31:0] data_store_6_58;
	reg [31:0] data_store_6_60;
	reg [31:0] global_state;
	reg [0:0] out_of_pipe_6_7;
	reg [0:0] out_of_pipe_bb_6_7;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_3_last_state;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;
	reg [31:0] state_4_last_state;
	reg [31:0] state_5_entry_BB_reg;
	reg [0:0] state_5_is_active;
	reg [31:0] state_5_last_BB_reg;
	reg [31:0] state_5_last_state;
	reg [31:0] state_6_entry_BB_reg;
	reg [0:0] state_6_is_active;
	reg [31:0] state_6_last_BB_reg;
	reg [31:0] state_6_last_state;
	reg [31:0] state_7_entry_BB_reg;
	reg [0:0] state_7_is_active;
	reg [31:0] state_7_last_BB_reg;
	reg [31:0] state_7_last_state;

	// controller for a.a_raddr_0_reg
	always @(*) begin
		if (andOp_140_out) begin 
			a_raddr_0_reg = add_add3_out;
		end else begin
			a_raddr_0_reg = 0;
		end
	end
	// controller for add_add15.add_add15_in0
	// controller for add_add15.add_add15_in1
	// Insensitive connections
	assign add_add15_in0 = b_rdata_0;
	assign add_add15_in1 = data_in_3_37_out_data;
	// controller for add_add17.add_add17_in0
	// controller for add_add17.add_add17_in1
	// Insensitive connections
	assign add_add17_in0 = data_in_6_59_out_data;
	assign add_add17_in1 = 32'd1;
	// controller for add_add3.add_add3_in0
	// controller for add_add3.add_add3_in1
	// Insensitive connections
	assign add_add3_in0 = phi_phi2_out;
	assign add_add3_in1 = tmp_output_131_out_data;
	// controller for add_add4.add_add4_in0
	// controller for add_add4.add_add4_in1
	// Insensitive connections
	assign add_add4_in0 = phi_phi2_out;
	assign add_add4_in1 = 32'd1;
	// controller for andOp_100.andOp_100_in0
	// controller for andOp_100.andOp_100_in1
	// Insensitive connections
	assign andOp_100_in0 = andOp_96_out;
	assign andOp_100_in1 = notOp_99_out;
	// controller for andOp_116.andOp_116_in0
	// controller for andOp_116.andOp_116_in1
	// Insensitive connections
	assign andOp_116_in0 = notOp_115_out;
	assign andOp_116_in1 = andOp_69_out;
	// controller for andOp_125.andOp_125_in0
	// controller for andOp_125.andOp_125_in1
	// Insensitive connections
	assign andOp_125_in0 = notOp_124_out;
	assign andOp_125_in1 = andOp_66_out;
	// controller for andOp_127.andOp_127_in0
	// controller for andOp_127.andOp_127_in1
	// Insensitive connections
	assign andOp_127_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_127_in1 = state_1_is_active;
	// controller for andOp_130.andOp_130_in0
	// controller for andOp_130.andOp_130_in1
	// Insensitive connections
	assign andOp_130_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_130_in1 = state_1_is_active;
	// controller for andOp_134.andOp_134_in0
	// controller for andOp_134.andOp_134_in1
	// Insensitive connections
	assign andOp_134_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_134_in1 = state_1_is_active;
	// controller for andOp_135.andOp_135_in0
	// controller for andOp_135.andOp_135_in1
	// Insensitive connections
	assign andOp_135_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_135_in1 = state_1_is_active;
	// controller for andOp_136.andOp_136_in0
	// controller for andOp_136.andOp_136_in1
	// Insensitive connections
	assign andOp_136_in0 = bb_1_active_in_state_1_out_data;
	assign andOp_136_in1 = state_1_is_active;
	// controller for andOp_139.andOp_139_in0
	// controller for andOp_139.andOp_139_in1
	// Insensitive connections
	assign andOp_139_in0 = bb_1_active_in_state_1_out_data;
	assign andOp_139_in1 = state_1_is_active;
	// controller for andOp_140.andOp_140_in0
	// controller for andOp_140.andOp_140_in1
	// Insensitive connections
	assign andOp_140_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_140_in1 = state_1_is_active;
	// controller for andOp_141.andOp_141_in0
	// controller for andOp_141.andOp_141_in1
	// Insensitive connections
	assign andOp_141_in0 = bb_4_active_in_state_2_out_data;
	assign andOp_141_in1 = state_2_is_active;
	// controller for andOp_142.andOp_142_in0
	// controller for andOp_142.andOp_142_in1
	// Insensitive connections
	assign andOp_142_in0 = bb_4_active_in_state_2_out_data;
	assign andOp_142_in1 = state_2_is_active;
	// controller for andOp_143.andOp_143_in0
	// controller for andOp_143.andOp_143_in1
	// Insensitive connections
	assign andOp_143_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_143_in1 = state_3_is_active;
	// controller for andOp_144.andOp_144_in0
	// controller for andOp_144.andOp_144_in1
	// Insensitive connections
	assign andOp_144_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_144_in1 = state_3_is_active;
	// controller for andOp_145.andOp_145_in0
	// controller for andOp_145.andOp_145_in1
	// Insensitive connections
	assign andOp_145_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_145_in1 = state_3_is_active;
	// controller for andOp_146.andOp_146_in0
	// controller for andOp_146.andOp_146_in1
	// Insensitive connections
	assign andOp_146_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_146_in1 = state_3_is_active;
	// controller for andOp_147.andOp_147_in0
	// controller for andOp_147.andOp_147_in1
	// Insensitive connections
	assign andOp_147_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_147_in1 = state_3_is_active;
	// controller for andOp_148.andOp_148_in0
	// controller for andOp_148.andOp_148_in1
	// Insensitive connections
	assign andOp_148_in0 = bb_3_active_in_state_6_out_data;
	assign andOp_148_in1 = state_6_is_active;
	// controller for andOp_149.andOp_149_in0
	// controller for andOp_149.andOp_149_in1
	// Insensitive connections
	assign andOp_149_in0 = bb_3_active_in_state_6_out_data;
	assign andOp_149_in1 = state_6_is_active;
	// controller for andOp_150.andOp_150_in0
	// controller for andOp_150.andOp_150_in1
	// Insensitive connections
	assign andOp_150_in0 = bb_2_active_in_state_7_out_data;
	assign andOp_150_in1 = state_7_is_active;
	// controller for andOp_151.andOp_151_in0
	// controller for andOp_151.andOp_151_in1
	// Insensitive connections
	assign andOp_151_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_151_in1 = state_1_is_active;
	// controller for andOp_152.andOp_152_in0
	// controller for andOp_152.andOp_152_in1
	// Insensitive connections
	assign andOp_152_in0 = bb_4_active_in_state_2_out_data;
	assign andOp_152_in1 = state_2_is_active;
	// controller for andOp_153.andOp_153_in0
	// controller for andOp_153.andOp_153_in1
	// Insensitive connections
	assign andOp_153_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_153_in1 = state_3_is_active;
	// controller for andOp_154.andOp_154_in0
	// controller for andOp_154.andOp_154_in1
	// Insensitive connections
	assign andOp_154_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_154_in1 = state_4_is_active;
	// controller for andOp_155.andOp_155_in0
	// controller for andOp_155.andOp_155_in1
	// Insensitive connections
	assign andOp_155_in0 = bb_4_active_in_state_5_out_data;
	assign andOp_155_in1 = state_5_is_active;
	// controller for andOp_157.andOp_157_in0
	// controller for andOp_157.andOp_157_in1
	// Insensitive connections
	assign andOp_157_in0 = 1'd1;
	assign andOp_157_in1 = notOp_156_out;
	// controller for andOp_159.andOp_159_in0
	// controller for andOp_159.andOp_159_in1
	// Insensitive connections
	assign andOp_159_in0 = andOp_157_out;
	assign andOp_159_in1 = notOp_158_out;
	// controller for andOp_161.andOp_161_in0
	// controller for andOp_161.andOp_161_in1
	// Insensitive connections
	assign andOp_161_in0 = andOp_159_out;
	assign andOp_161_in1 = notOp_160_out;
	// controller for andOp_163.andOp_163_in0
	// controller for andOp_163.andOp_163_in1
	// Insensitive connections
	assign andOp_163_in0 = andOp_161_out;
	assign andOp_163_in1 = notOp_162_out;
	// controller for andOp_165.andOp_165_in0
	// controller for andOp_165.andOp_165_in1
	// Insensitive connections
	assign andOp_165_in0 = andOp_163_out;
	assign andOp_165_in1 = notOp_164_out;
	// controller for andOp_166.andOp_166_in0
	// controller for andOp_166.andOp_166_in1
	// Insensitive connections
	assign andOp_166_in0 = in_pipeline_0_out_data;
	assign andOp_166_in1 = andOp_165_out;
	// controller for andOp_167.andOp_167_in0
	// controller for andOp_167.andOp_167_in1
	// Insensitive connections
	assign andOp_167_in0 = andOp_166_out;
	assign andOp_167_in1 = out_of_pipe_6_7;
	// controller for andOp_168.andOp_168_in0
	// controller for andOp_168.andOp_168_in1
	// Insensitive connections
	assign andOp_168_in0 = andOp_166_out;
	assign andOp_168_in1 = out_of_pipe_6_7;
	// controller for andOp_170.andOp_170_in0
	// controller for andOp_170.andOp_170_in1
	// Insensitive connections
	assign andOp_170_in0 = 1'd1;
	assign andOp_170_in1 = notOp_169_out;
	// controller for andOp_172.andOp_172_in0
	// controller for andOp_172.andOp_172_in1
	// Insensitive connections
	assign andOp_172_in0 = andOp_170_out;
	assign andOp_172_in1 = notOp_171_out;
	// controller for andOp_174.andOp_174_in0
	// controller for andOp_174.andOp_174_in1
	// Insensitive connections
	assign andOp_174_in0 = andOp_172_out;
	assign andOp_174_in1 = notOp_173_out;
	// controller for andOp_176.andOp_176_in0
	// controller for andOp_176.andOp_176_in1
	// Insensitive connections
	assign andOp_176_in0 = andOp_174_out;
	assign andOp_176_in1 = notOp_175_out;
	// controller for andOp_178.andOp_178_in0
	// controller for andOp_178.andOp_178_in1
	// Insensitive connections
	assign andOp_178_in0 = andOp_176_out;
	assign andOp_178_in1 = notOp_177_out;
	// controller for andOp_179.andOp_179_in0
	// controller for andOp_179.andOp_179_in1
	// Insensitive connections
	assign andOp_179_in0 = in_pipeline_0_out_data;
	assign andOp_179_in1 = andOp_178_out;
	// controller for andOp_180.andOp_180_in0
	// controller for andOp_180.andOp_180_in1
	// Insensitive connections
	assign andOp_180_in0 = andOp_179_out;
	assign andOp_180_in1 = out_of_pipe_bb_6_7;
	// controller for andOp_181.andOp_181_in0
	// controller for andOp_181.andOp_181_in1
	// Insensitive connections
	assign andOp_181_in0 = bb_2_active_in_state_7_out_data;
	assign andOp_181_in1 = state_7_is_active;
	// controller for andOp_183.andOp_183_in0
	// controller for andOp_183.andOp_183_in1
	// Insensitive connections
	assign andOp_183_in0 = notOp_182_out;
	assign andOp_183_in1 = 1'd1;
	// controller for andOp_185.andOp_185_in0
	// controller for andOp_185.andOp_185_in1
	// Insensitive connections
	assign andOp_185_in0 = notOp_184_out;
	assign andOp_185_in1 = andOp_183_out;
	// controller for andOp_187.andOp_187_in0
	// controller for andOp_187.andOp_187_in1
	// Insensitive connections
	assign andOp_187_in0 = notOp_186_out;
	assign andOp_187_in1 = andOp_185_out;
	// controller for andOp_189.andOp_189_in0
	// controller for andOp_189.andOp_189_in1
	// Insensitive connections
	assign andOp_189_in0 = notOp_188_out;
	assign andOp_189_in1 = 1'd1;
	// controller for andOp_191.andOp_191_in0
	// controller for andOp_191.andOp_191_in1
	// Insensitive connections
	assign andOp_191_in0 = notOp_190_out;
	assign andOp_191_in1 = 1'd1;
	// controller for andOp_193.andOp_193_in0
	// controller for andOp_193.andOp_193_in1
	// Insensitive connections
	assign andOp_193_in0 = notOp_192_out;
	assign andOp_193_in1 = 1'd1;
	// controller for andOp_195.andOp_195_in0
	// controller for andOp_195.andOp_195_in1
	// Insensitive connections
	assign andOp_195_in0 = notOp_194_out;
	assign andOp_195_in1 = 1'd1;
	// controller for andOp_197.andOp_197_in0
	// controller for andOp_197.andOp_197_in1
	// Insensitive connections
	assign andOp_197_in0 = notOp_196_out;
	assign andOp_197_in1 = 1'd1;
	// controller for andOp_199.andOp_199_in0
	// controller for andOp_199.andOp_199_in1
	// Insensitive connections
	assign andOp_199_in0 = notOp_198_out;
	assign andOp_199_in1 = andOp_197_out;
	// controller for andOp_201.andOp_201_in0
	// controller for andOp_201.andOp_201_in1
	// Insensitive connections
	assign andOp_201_in0 = notOp_200_out;
	assign andOp_201_in1 = 1'd1;
	// controller for andOp_203.andOp_203_in0
	// controller for andOp_203.andOp_203_in1
	// Insensitive connections
	assign andOp_203_in0 = notOp_202_out;
	assign andOp_203_in1 = andOp_201_out;
	// controller for andOp_214.andOp_214_in0
	// controller for andOp_214.andOp_214_in1
	// Insensitive connections
	assign andOp_214_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_214_in1 = state_1_is_active;
	// controller for andOp_215.andOp_215_in0
	// controller for andOp_215.andOp_215_in1
	// Insensitive connections
	assign andOp_215_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_215_in1 = state_1_is_active;
	// controller for andOp_216.andOp_216_in0
	// controller for andOp_216.andOp_216_in1
	// Insensitive connections
	assign andOp_216_in0 = bb_1_active_in_state_1_out_data;
	assign andOp_216_in1 = state_1_is_active;
	// controller for andOp_217.andOp_217_in0
	// controller for andOp_217.andOp_217_in1
	// Insensitive connections
	assign andOp_217_in0 = bb_1_active_in_state_1_out_data;
	assign andOp_217_in1 = state_1_is_active;
	// controller for andOp_220.andOp_220_in0
	// controller for andOp_220.andOp_220_in1
	// Insensitive connections
	assign andOp_220_in0 = bb_4_active_in_state_2_out_data;
	assign andOp_220_in1 = state_2_is_active;
	// controller for andOp_230.andOp_230_in0
	// controller for andOp_230.andOp_230_in1
	// Insensitive connections
	assign andOp_230_in0 = bb_3_active_in_state_6_out_data;
	assign andOp_230_in1 = state_6_is_active;
	// controller for andOp_62.andOp_62_in0
	// controller for andOp_62.andOp_62_in1
	// Insensitive connections
	assign andOp_62_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_62_in1 = state_0_is_active;
	// controller for andOp_64.andOp_64_in0
	// controller for andOp_64.andOp_64_in1
	// Insensitive connections
	assign andOp_64_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_64_in1 = state_1_is_active;
	// controller for andOp_66.andOp_66_in0
	// controller for andOp_66.andOp_66_in1
	// Insensitive connections
	assign andOp_66_in0 = andOp_64_out;
	assign andOp_66_in1 = icmp_icmp5_out;
	// controller for andOp_68.andOp_68_in0
	// controller for andOp_68.andOp_68_in1
	// Insensitive connections
	assign andOp_68_in0 = andOp_64_out;
	assign andOp_68_in1 = notOp_67_out;
	// controller for andOp_69.andOp_69_in0
	// controller for andOp_69.andOp_69_in1
	// Insensitive connections
	assign andOp_69_in0 = bb_1_active_in_state_1_out_data;
	assign andOp_69_in1 = state_1_is_active;
	// controller for andOp_71.andOp_71_in0
	// controller for andOp_71.andOp_71_in1
	// Insensitive connections
	assign andOp_71_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_71_in1 = state_1_is_active;
	// controller for andOp_73.andOp_73_in0
	// controller for andOp_73.andOp_73_in1
	// Insensitive connections
	assign andOp_73_in0 = andOp_71_out;
	assign andOp_73_in1 = icmp_icmp5_out;
	// controller for andOp_75.andOp_75_in0
	// controller for andOp_75.andOp_75_in1
	// Insensitive connections
	assign andOp_75_in0 = andOp_71_out;
	assign andOp_75_in1 = notOp_74_out;
	// controller for andOp_76.andOp_76_in0
	// controller for andOp_76.andOp_76_in1
	// Insensitive connections
	assign andOp_76_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_76_in1 = state_1_is_active;
	// controller for andOp_78.andOp_78_in0
	// controller for andOp_78.andOp_78_in1
	// Insensitive connections
	assign andOp_78_in0 = andOp_76_out;
	assign andOp_78_in1 = icmp_icmp5_out;
	// controller for andOp_80.andOp_80_in0
	// controller for andOp_80.andOp_80_in1
	// Insensitive connections
	assign andOp_80_in0 = andOp_76_out;
	assign andOp_80_in1 = notOp_79_out;
	// controller for andOp_81.andOp_81_in0
	// controller for andOp_81.andOp_81_in1
	// Insensitive connections
	assign andOp_81_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_81_in1 = state_1_is_active;
	// controller for andOp_83.andOp_83_in0
	// controller for andOp_83.andOp_83_in1
	// Insensitive connections
	assign andOp_83_in0 = andOp_81_out;
	assign andOp_83_in1 = icmp_icmp5_out;
	// controller for andOp_85.andOp_85_in0
	// controller for andOp_85.andOp_85_in1
	// Insensitive connections
	assign andOp_85_in0 = andOp_81_out;
	assign andOp_85_in1 = notOp_84_out;
	// controller for andOp_86.andOp_86_in0
	// controller for andOp_86.andOp_86_in1
	// Insensitive connections
	assign andOp_86_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_86_in1 = state_1_is_active;
	// controller for andOp_88.andOp_88_in0
	// controller for andOp_88.andOp_88_in1
	// Insensitive connections
	assign andOp_88_in0 = andOp_86_out;
	assign andOp_88_in1 = icmp_icmp5_out;
	// controller for andOp_90.andOp_90_in0
	// controller for andOp_90.andOp_90_in1
	// Insensitive connections
	assign andOp_90_in0 = andOp_86_out;
	assign andOp_90_in1 = notOp_89_out;
	// controller for andOp_91.andOp_91_in0
	// controller for andOp_91.andOp_91_in1
	// Insensitive connections
	assign andOp_91_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_91_in1 = state_1_is_active;
	// controller for andOp_93.andOp_93_in0
	// controller for andOp_93.andOp_93_in1
	// Insensitive connections
	assign andOp_93_in0 = andOp_91_out;
	assign andOp_93_in1 = icmp_icmp5_out;
	// controller for andOp_95.andOp_95_in0
	// controller for andOp_95.andOp_95_in1
	// Insensitive connections
	assign andOp_95_in0 = andOp_91_out;
	assign andOp_95_in1 = notOp_94_out;
	// controller for andOp_96.andOp_96_in0
	// controller for andOp_96.andOp_96_in1
	// Insensitive connections
	assign andOp_96_in0 = bb_3_active_in_state_6_out_data;
	assign andOp_96_in1 = state_6_is_active;
	// controller for andOp_98.andOp_98_in0
	// controller for andOp_98.andOp_98_in1
	// Insensitive connections
	assign andOp_98_in0 = andOp_96_out;
	assign andOp_98_in1 = icmp_icmp18_out;
	// controller for b.b_raddr_0_reg
	always @(*) begin
		if (andOp_142_out) begin 
			b_raddr_0_reg = data_in_2_20_out_data;
		end else begin
			b_raddr_0_reg = 0;
		end
	end
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_101_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_113_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_1.bb_1_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_1_in_data = eq_104_out;
		end else begin
			bb_1_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_1.bb_1_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_117_out) begin 
			bb_1_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_7.bb_2_active_in_state_7_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_7_in_data = eq_112_out;
		end else begin
			bb_2_active_in_state_7_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_7.bb_2_predecessor_in_state_7_in_data
	always @(*) begin
		if (eq_126_out) begin 
			bb_2_predecessor_in_state_7_in_data = state_7_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_7_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_6.bb_3_active_in_state_6_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_6_in_data = orOp_111_out;
		end else begin
			bb_3_active_in_state_6_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_6.bb_3_predecessor_in_state_6_in_data
	always @(*) begin
		if (andOp_125_out) begin 
			bb_3_predecessor_in_state_6_in_data = 32'd4;
		end else if (eq_123_out) begin 
			bb_3_predecessor_in_state_6_in_data = state_6_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_6_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_1.bb_4_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_1_in_data = orOp_103_out;
		end else begin
			bb_4_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_2.bb_4_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_2_in_data = eq_105_out;
		end else begin
			bb_4_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_3.bb_4_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_3_in_data = eq_106_out;
		end else begin
			bb_4_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_4.bb_4_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_4_in_data = eq_107_out;
		end else begin
			bb_4_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_5.bb_4_active_in_state_5_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_5_in_data = eq_108_out;
		end else begin
			bb_4_active_in_state_5_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_6.bb_4_active_in_state_6_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_6_in_data = eq_109_out;
		end else begin
			bb_4_active_in_state_6_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_1.bb_4_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_116_out) begin 
			bb_4_predecessor_in_state_1_in_data = 32'd1;
		end else if (eq_114_out) begin 
			bb_4_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_2.bb_4_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_118_out) begin 
			bb_4_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_3.bb_4_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_119_out) begin 
			bb_4_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_4.bb_4_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_120_out) begin 
			bb_4_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_5.bb_4_predecessor_in_state_5_in_data
	always @(*) begin
		if (eq_121_out) begin 
			bb_4_predecessor_in_state_5_in_data = state_5_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_5_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_6.bb_4_predecessor_in_state_6_in_data
	always @(*) begin
		if (eq_122_out) begin 
			bb_4_predecessor_in_state_6_in_data = state_6_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_6_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_62_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_63_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_1_happened_in_state_1.br_1_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_69_out) begin 
			br_1_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_70_out) begin 
			br_1_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_1_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_6.br_3_happened_in_state_6_in_data
	always @(*) begin
		if (andOp_96_out) begin 
			br_3_happened_in_state_6_in_data = 1'd1;
		end else if (notOp_97_out) begin 
			br_3_happened_in_state_6_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_6_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_1.br_4_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_64_out) begin 
			br_4_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_65_out) begin 
			br_4_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_2.br_4_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_71_out) begin 
			br_4_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_72_out) begin 
			br_4_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_3.br_4_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_76_out) begin 
			br_4_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_77_out) begin 
			br_4_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_4.br_4_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_81_out) begin 
			br_4_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_82_out) begin 
			br_4_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_5.br_4_happened_in_state_5_in_data
	always @(*) begin
		if (andOp_86_out) begin 
			br_4_happened_in_state_5_in_data = 1'd1;
		end else if (notOp_87_out) begin 
			br_4_happened_in_state_5_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_5_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_6.br_4_happened_in_state_6_in_data
	always @(*) begin
		if (andOp_91_out) begin 
			br_4_happened_in_state_6_in_data = 1'd1;
		end else if (notOp_92_out) begin 
			br_4_happened_in_state_6_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_6_in_data = 0;
		end
	end
	// controller for c.c_waddr_0_reg
	always @(*) begin
		if (andOp_145_out) begin 
			c_waddr_0_reg = data_in_3_30_out_data;
		end else begin
			c_waddr_0_reg = 0;
		end
	end
	// controller for c.c_wdata_0_reg
	always @(*) begin
		if (andOp_146_out) begin 
			c_wdata_0_reg = add_add15_out;
		end else begin
			c_wdata_0_reg = 0;
		end
	end
	// controller for c.c_wen_0_reg
	always @(*) begin
		if (andOp_144_out) begin 
			c_wen_0_reg = -(1'd1);
		end else begin
			c_wen_0_reg = 0;
		end
	end
	// controller for concat_128.concat_128_in0
	// controller for concat_128.concat_128_in1
	// Insensitive connections
	assign concat_128_in0 = data_in_1_12_out_data;
	assign concat_128_in1 = 32'd0;
	// controller for concat_129.concat_129_in0
	// controller for concat_129.concat_129_in1
	// Insensitive connections
	assign concat_129_in0 = 32'd4;
	assign concat_129_in1 = 32'd1;
	// controller for concat_137.concat_137_in0
	// controller for concat_137.concat_137_in1
	// Insensitive connections
	assign concat_137_in0 = data_in_1_9_out_data;
	assign concat_137_in1 = 32'd0;
	// controller for concat_138.concat_138_in0
	// controller for concat_138.concat_138_in1
	// Insensitive connections
	assign concat_138_in0 = 32'd3;
	assign concat_138_in1 = 32'd0;
	// controller for data_in_0_1.data_in_0_1_in_data
	always @(*) begin
		if (eq_210_out) begin 
			data_in_0_1_in_data = data_store_0_0;
		end else begin
			data_in_0_1_in_data = 0;
		end
	end
	// controller for data_in_0_3.data_in_0_3_in_data
	always @(*) begin
		if (eq_210_out) begin 
			data_in_0_3_in_data = data_store_0_2;
		end else begin
			data_in_0_3_in_data = 0;
		end
	end
	// controller for data_in_0_5.data_in_0_5_in_data
	always @(*) begin
		if (eq_210_out) begin 
			data_in_0_5_in_data = data_store_0_4;
		end else begin
			data_in_0_5_in_data = 0;
		end
	end
	// controller for data_in_0_7.data_in_0_7_in_data
	always @(*) begin
		if (eq_210_out) begin 
			data_in_0_7_in_data = data_store_0_6;
		end else begin
			data_in_0_7_in_data = 0;
		end
	end
	// controller for data_in_1_12.data_in_1_12_in_data
	always @(*) begin
		if (eq_211_out) begin 
			data_in_1_12_in_data = data_store_0_2;
		end else if (eq_212_out) begin 
			data_in_1_12_in_data = data_store_1_11;
		end else if (eq_213_out) begin 
			data_in_1_12_in_data = data_store_6_56;
		end else begin
			data_in_1_12_in_data = 0;
		end
	end
	// controller for data_in_1_14.data_in_1_14_in_data
	always @(*) begin
		if (eq_211_out) begin 
			data_in_1_14_in_data = data_store_0_4;
		end else if (eq_212_out) begin 
			data_in_1_14_in_data = data_store_1_13;
		end else if (eq_213_out) begin 
			data_in_1_14_in_data = data_store_6_58;
		end else begin
			data_in_1_14_in_data = 0;
		end
	end
	// controller for data_in_1_16.data_in_1_16_in_data
	always @(*) begin
		if (eq_211_out) begin 
			data_in_1_16_in_data = data_store_0_6;
		end else if (eq_212_out) begin 
			data_in_1_16_in_data = data_store_1_15;
		end else if (eq_213_out) begin 
			data_in_1_16_in_data = data_store_6_60;
		end else begin
			data_in_1_16_in_data = 0;
		end
	end
	// controller for data_in_1_9.data_in_1_9_in_data
	always @(*) begin
		if (eq_211_out) begin 
			data_in_1_9_in_data = data_store_0_0;
		end else if (eq_212_out) begin 
			data_in_1_9_in_data = data_store_1_8;
		end else if (eq_213_out) begin 
			data_in_1_9_in_data = data_store_6_54;
		end else begin
			data_in_1_9_in_data = 0;
		end
	end
	// controller for data_in_2_18.data_in_2_18_in_data
	always @(*) begin
		if (eq_218_out) begin 
			data_in_2_18_in_data = data_store_1_8;
		end else if (eq_219_out) begin 
			data_in_2_18_in_data = data_store_2_17;
		end else begin
			data_in_2_18_in_data = 0;
		end
	end
	// controller for data_in_2_20.data_in_2_20_in_data
	always @(*) begin
		if (eq_218_out) begin 
			data_in_2_20_in_data = data_store_1_10;
		end else if (eq_219_out) begin 
			data_in_2_20_in_data = data_store_2_19;
		end else begin
			data_in_2_20_in_data = 0;
		end
	end
	// controller for data_in_2_22.data_in_2_22_in_data
	always @(*) begin
		if (eq_218_out) begin 
			data_in_2_22_in_data = data_store_1_11;
		end else if (eq_219_out) begin 
			data_in_2_22_in_data = data_store_2_21;
		end else begin
			data_in_2_22_in_data = 0;
		end
	end
	// controller for data_in_2_24.data_in_2_24_in_data
	always @(*) begin
		if (eq_218_out) begin 
			data_in_2_24_in_data = data_store_1_13;
		end else if (eq_219_out) begin 
			data_in_2_24_in_data = data_store_2_23;
		end else begin
			data_in_2_24_in_data = 0;
		end
	end
	// controller for data_in_2_26.data_in_2_26_in_data
	always @(*) begin
		if (eq_218_out) begin 
			data_in_2_26_in_data = data_store_1_15;
		end else if (eq_219_out) begin 
			data_in_2_26_in_data = data_store_2_25;
		end else begin
			data_in_2_26_in_data = 0;
		end
	end
	// controller for data_in_3_29.data_in_3_29_in_data
	always @(*) begin
		if (eq_221_out) begin 
			data_in_3_29_in_data = data_store_2_17;
		end else if (eq_222_out) begin 
			data_in_3_29_in_data = data_store_3_28;
		end else begin
			data_in_3_29_in_data = 0;
		end
	end
	// controller for data_in_3_30.data_in_3_30_in_data
	always @(*) begin
		if (eq_221_out) begin 
			data_in_3_30_in_data = data_store_2_19;
		end else if (eq_222_out) begin 
			data_in_3_30_in_data = 32'd0;
		end else begin
			data_in_3_30_in_data = 0;
		end
	end
	// controller for data_in_3_32.data_in_3_32_in_data
	always @(*) begin
		if (eq_221_out) begin 
			data_in_3_32_in_data = data_store_2_21;
		end else if (eq_222_out) begin 
			data_in_3_32_in_data = data_store_3_31;
		end else begin
			data_in_3_32_in_data = 0;
		end
	end
	// controller for data_in_3_34.data_in_3_34_in_data
	always @(*) begin
		if (eq_221_out) begin 
			data_in_3_34_in_data = data_store_2_23;
		end else if (eq_222_out) begin 
			data_in_3_34_in_data = data_store_3_33;
		end else begin
			data_in_3_34_in_data = 0;
		end
	end
	// controller for data_in_3_36.data_in_3_36_in_data
	always @(*) begin
		if (eq_221_out) begin 
			data_in_3_36_in_data = data_store_2_25;
		end else if (eq_222_out) begin 
			data_in_3_36_in_data = data_store_3_35;
		end else begin
			data_in_3_36_in_data = 0;
		end
	end
	// controller for data_in_3_37.data_in_3_37_in_data
	always @(*) begin
		if (eq_221_out) begin 
			data_in_3_37_in_data = data_store_2_27;
		end else if (eq_222_out) begin 
			data_in_3_37_in_data = 32'd0;
		end else begin
			data_in_3_37_in_data = 0;
		end
	end
	// controller for data_in_4_39.data_in_4_39_in_data
	always @(*) begin
		if (eq_223_out) begin 
			data_in_4_39_in_data = data_store_3_28;
		end else if (eq_224_out) begin 
			data_in_4_39_in_data = data_store_4_38;
		end else begin
			data_in_4_39_in_data = 0;
		end
	end
	// controller for data_in_4_41.data_in_4_41_in_data
	always @(*) begin
		if (eq_223_out) begin 
			data_in_4_41_in_data = data_store_3_31;
		end else if (eq_224_out) begin 
			data_in_4_41_in_data = data_store_4_40;
		end else begin
			data_in_4_41_in_data = 0;
		end
	end
	// controller for data_in_4_43.data_in_4_43_in_data
	always @(*) begin
		if (eq_223_out) begin 
			data_in_4_43_in_data = data_store_3_33;
		end else if (eq_224_out) begin 
			data_in_4_43_in_data = data_store_4_42;
		end else begin
			data_in_4_43_in_data = 0;
		end
	end
	// controller for data_in_4_45.data_in_4_45_in_data
	always @(*) begin
		if (eq_223_out) begin 
			data_in_4_45_in_data = data_store_3_35;
		end else if (eq_224_out) begin 
			data_in_4_45_in_data = data_store_4_44;
		end else begin
			data_in_4_45_in_data = 0;
		end
	end
	// controller for data_in_5_47.data_in_5_47_in_data
	always @(*) begin
		if (eq_225_out) begin 
			data_in_5_47_in_data = data_store_4_38;
		end else if (eq_226_out) begin 
			data_in_5_47_in_data = data_store_5_46;
		end else begin
			data_in_5_47_in_data = 0;
		end
	end
	// controller for data_in_5_49.data_in_5_49_in_data
	always @(*) begin
		if (eq_225_out) begin 
			data_in_5_49_in_data = data_store_4_40;
		end else if (eq_226_out) begin 
			data_in_5_49_in_data = data_store_5_48;
		end else begin
			data_in_5_49_in_data = 0;
		end
	end
	// controller for data_in_5_51.data_in_5_51_in_data
	always @(*) begin
		if (eq_225_out) begin 
			data_in_5_51_in_data = data_store_4_42;
		end else if (eq_226_out) begin 
			data_in_5_51_in_data = data_store_5_50;
		end else begin
			data_in_5_51_in_data = 0;
		end
	end
	// controller for data_in_5_53.data_in_5_53_in_data
	always @(*) begin
		if (eq_225_out) begin 
			data_in_5_53_in_data = data_store_4_44;
		end else if (eq_226_out) begin 
			data_in_5_53_in_data = data_store_5_52;
		end else begin
			data_in_5_53_in_data = 0;
		end
	end
	// controller for data_in_6_55.data_in_6_55_in_data
	always @(*) begin
		if (eq_227_out) begin 
			data_in_6_55_in_data = data_store_1_8;
		end else if (eq_228_out) begin 
			data_in_6_55_in_data = data_store_5_46;
		end else if (eq_229_out) begin 
			data_in_6_55_in_data = data_store_6_54;
		end else begin
			data_in_6_55_in_data = 0;
		end
	end
	// controller for data_in_6_57.data_in_6_57_in_data
	always @(*) begin
		if (eq_227_out) begin 
			data_in_6_57_in_data = data_store_1_11;
		end else if (eq_228_out) begin 
			data_in_6_57_in_data = data_store_5_48;
		end else if (eq_229_out) begin 
			data_in_6_57_in_data = data_store_6_56;
		end else begin
			data_in_6_57_in_data = 0;
		end
	end
	// controller for data_in_6_59.data_in_6_59_in_data
	always @(*) begin
		if (eq_227_out) begin 
			data_in_6_59_in_data = data_store_1_13;
		end else if (eq_228_out) begin 
			data_in_6_59_in_data = data_store_5_50;
		end else if (eq_229_out) begin 
			data_in_6_59_in_data = data_store_6_58;
		end else begin
			data_in_6_59_in_data = 0;
		end
	end
	// controller for data_in_6_61.data_in_6_61_in_data
	always @(*) begin
		if (eq_227_out) begin 
			data_in_6_61_in_data = data_store_1_15;
		end else if (eq_228_out) begin 
			data_in_6_61_in_data = data_store_5_52;
		end else if (eq_229_out) begin 
			data_in_6_61_in_data = data_store_6_60;
		end else begin
			data_in_6_61_in_data = 0;
		end
	end
	// controller for eq_101.eq_101_in0
	// controller for eq_101.eq_101_in1
	// Insensitive connections
	assign eq_101_in0 = 32'd0;
	assign eq_101_in1 = state_0_entry_BB_reg;
	// controller for eq_102.eq_102_in0
	// controller for eq_102.eq_102_in1
	// Insensitive connections
	assign eq_102_in0 = 32'd4;
	assign eq_102_in1 = state_1_entry_BB_reg;
	// controller for eq_104.eq_104_in0
	// controller for eq_104.eq_104_in1
	// Insensitive connections
	assign eq_104_in0 = 32'd1;
	assign eq_104_in1 = state_1_entry_BB_reg;
	// controller for eq_105.eq_105_in0
	// controller for eq_105.eq_105_in1
	// Insensitive connections
	assign eq_105_in0 = 32'd4;
	assign eq_105_in1 = state_2_entry_BB_reg;
	// controller for eq_106.eq_106_in0
	// controller for eq_106.eq_106_in1
	// Insensitive connections
	assign eq_106_in0 = 32'd4;
	assign eq_106_in1 = state_3_entry_BB_reg;
	// controller for eq_107.eq_107_in0
	// controller for eq_107.eq_107_in1
	// Insensitive connections
	assign eq_107_in0 = 32'd4;
	assign eq_107_in1 = state_4_entry_BB_reg;
	// controller for eq_108.eq_108_in0
	// controller for eq_108.eq_108_in1
	// Insensitive connections
	assign eq_108_in0 = 32'd4;
	assign eq_108_in1 = state_5_entry_BB_reg;
	// controller for eq_109.eq_109_in0
	// controller for eq_109.eq_109_in1
	// Insensitive connections
	assign eq_109_in0 = 32'd4;
	assign eq_109_in1 = state_6_entry_BB_reg;
	// controller for eq_110.eq_110_in0
	// controller for eq_110.eq_110_in1
	// Insensitive connections
	assign eq_110_in0 = 32'd3;
	assign eq_110_in1 = state_6_entry_BB_reg;
	// controller for eq_112.eq_112_in0
	// controller for eq_112.eq_112_in1
	// Insensitive connections
	assign eq_112_in0 = 32'd2;
	assign eq_112_in1 = state_7_entry_BB_reg;
	// controller for eq_113.eq_113_in0
	// controller for eq_113.eq_113_in1
	// Insensitive connections
	assign eq_113_in0 = 32'd0;
	assign eq_113_in1 = state_0_entry_BB_reg;
	// controller for eq_114.eq_114_in0
	// controller for eq_114.eq_114_in1
	// Insensitive connections
	assign eq_114_in0 = 32'd4;
	assign eq_114_in1 = state_1_entry_BB_reg;
	// controller for eq_117.eq_117_in0
	// controller for eq_117.eq_117_in1
	// Insensitive connections
	assign eq_117_in0 = 32'd1;
	assign eq_117_in1 = state_1_entry_BB_reg;
	// controller for eq_118.eq_118_in0
	// controller for eq_118.eq_118_in1
	// Insensitive connections
	assign eq_118_in0 = 32'd4;
	assign eq_118_in1 = state_2_entry_BB_reg;
	// controller for eq_119.eq_119_in0
	// controller for eq_119.eq_119_in1
	// Insensitive connections
	assign eq_119_in0 = 32'd4;
	assign eq_119_in1 = state_3_entry_BB_reg;
	// controller for eq_120.eq_120_in0
	// controller for eq_120.eq_120_in1
	// Insensitive connections
	assign eq_120_in0 = 32'd4;
	assign eq_120_in1 = state_4_entry_BB_reg;
	// controller for eq_121.eq_121_in0
	// controller for eq_121.eq_121_in1
	// Insensitive connections
	assign eq_121_in0 = 32'd4;
	assign eq_121_in1 = state_5_entry_BB_reg;
	// controller for eq_122.eq_122_in0
	// controller for eq_122.eq_122_in1
	// Insensitive connections
	assign eq_122_in0 = 32'd4;
	assign eq_122_in1 = state_6_entry_BB_reg;
	// controller for eq_123.eq_123_in0
	// controller for eq_123.eq_123_in1
	// Insensitive connections
	assign eq_123_in0 = 32'd3;
	assign eq_123_in1 = state_6_entry_BB_reg;
	// controller for eq_126.eq_126_in0
	// controller for eq_126.eq_126_in1
	// Insensitive connections
	assign eq_126_in0 = 32'd2;
	assign eq_126_in1 = state_7_entry_BB_reg;
	// controller for eq_132.eq_132_in0
	// controller for eq_132.eq_132_in1
	// Insensitive connections
	assign eq_132_in0 = 32'd4;
	assign eq_132_in1 = state_1_entry_BB_reg;
	// controller for eq_133.eq_133_in0
	// controller for eq_133.eq_133_in1
	// Insensitive connections
	assign eq_133_in0 = 32'd1;
	assign eq_133_in1 = state_1_entry_BB_reg;
	// controller for eq_210.eq_210_in0
	// controller for eq_210.eq_210_in1
	// Insensitive connections
	assign eq_210_in0 = 32'd0;
	assign eq_210_in1 = state_0_last_state;
	// controller for eq_211.eq_211_in0
	// controller for eq_211.eq_211_in1
	// Insensitive connections
	assign eq_211_in0 = 32'd0;
	assign eq_211_in1 = state_1_last_state;
	// controller for eq_212.eq_212_in0
	// controller for eq_212.eq_212_in1
	// Insensitive connections
	assign eq_212_in0 = 32'd1;
	assign eq_212_in1 = state_1_last_state;
	// controller for eq_213.eq_213_in0
	// controller for eq_213.eq_213_in1
	// Insensitive connections
	assign eq_213_in0 = 32'd6;
	assign eq_213_in1 = state_1_last_state;
	// controller for eq_218.eq_218_in0
	// controller for eq_218.eq_218_in1
	// Insensitive connections
	assign eq_218_in0 = 32'd1;
	assign eq_218_in1 = state_2_last_state;
	// controller for eq_219.eq_219_in0
	// controller for eq_219.eq_219_in1
	// Insensitive connections
	assign eq_219_in0 = 32'd2;
	assign eq_219_in1 = state_2_last_state;
	// controller for eq_221.eq_221_in0
	// controller for eq_221.eq_221_in1
	// Insensitive connections
	assign eq_221_in0 = 32'd2;
	assign eq_221_in1 = state_3_last_state;
	// controller for eq_222.eq_222_in0
	// controller for eq_222.eq_222_in1
	// Insensitive connections
	assign eq_222_in0 = 32'd3;
	assign eq_222_in1 = state_3_last_state;
	// controller for eq_223.eq_223_in0
	// controller for eq_223.eq_223_in1
	// Insensitive connections
	assign eq_223_in0 = 32'd3;
	assign eq_223_in1 = state_4_last_state;
	// controller for eq_224.eq_224_in0
	// controller for eq_224.eq_224_in1
	// Insensitive connections
	assign eq_224_in0 = 32'd4;
	assign eq_224_in1 = state_4_last_state;
	// controller for eq_225.eq_225_in0
	// controller for eq_225.eq_225_in1
	// Insensitive connections
	assign eq_225_in0 = 32'd4;
	assign eq_225_in1 = state_5_last_state;
	// controller for eq_226.eq_226_in0
	// controller for eq_226.eq_226_in1
	// Insensitive connections
	assign eq_226_in0 = 32'd5;
	assign eq_226_in1 = state_5_last_state;
	// controller for eq_227.eq_227_in0
	// controller for eq_227.eq_227_in1
	// Insensitive connections
	assign eq_227_in0 = 32'd1;
	assign eq_227_in1 = state_6_last_state;
	// controller for eq_228.eq_228_in0
	// controller for eq_228.eq_228_in1
	// Insensitive connections
	assign eq_228_in0 = 32'd5;
	assign eq_228_in1 = state_6_last_state;
	// controller for eq_229.eq_229_in0
	// controller for eq_229.eq_229_in1
	// Insensitive connections
	assign eq_229_in0 = 32'd6;
	assign eq_229_in1 = state_6_last_state;
	// controller for eq_231.eq_231_in0
	// controller for eq_231.eq_231_in1
	// Insensitive connections
	assign eq_231_in0 = 32'd6;
	assign eq_231_in1 = state_7_last_state;
	// controller for eq_232.eq_232_in0
	// controller for eq_232.eq_232_in1
	// Insensitive connections
	assign eq_232_in0 = 32'd7;
	assign eq_232_in1 = state_7_last_state;
	// controller for icmp_icmp18.icmp_icmp18_in0
	// controller for icmp_icmp18.icmp_icmp18_in1
	// Insensitive connections
	assign icmp_icmp18_in0 = add_add17_out;
	assign icmp_icmp18_in1 = 32'd16;
	// controller for icmp_icmp5.icmp_icmp5_in0
	// controller for icmp_icmp5.icmp_icmp5_in1
	// Insensitive connections
	assign icmp_icmp5_in0 = add_add4_out;
	assign icmp_icmp5_in1 = 32'd16;
	// controller for in_pipeline_0.in_pipeline_0_in_data
	always @(*) begin
		if (1'd1) begin 
			in_pipeline_0_in_data = orOp_209_out;
		end else begin
			in_pipeline_0_in_data = 0;
		end
	end
	// controller for notOp_115.notOp_115_in0
	// Insensitive connections
	assign notOp_115_in0 = eq_114_out;
	// controller for notOp_124.notOp_124_in0
	// Insensitive connections
	assign notOp_124_in0 = eq_123_out;
	// controller for notOp_156.notOp_156_in0
	// Insensitive connections
	assign notOp_156_in0 = state_1_is_active;
	// controller for notOp_158.notOp_158_in0
	// Insensitive connections
	assign notOp_158_in0 = state_2_is_active;
	// controller for notOp_160.notOp_160_in0
	// Insensitive connections
	assign notOp_160_in0 = state_3_is_active;
	// controller for notOp_162.notOp_162_in0
	// Insensitive connections
	assign notOp_162_in0 = state_4_is_active;
	// controller for notOp_164.notOp_164_in0
	// Insensitive connections
	assign notOp_164_in0 = state_5_is_active;
	// controller for notOp_169.notOp_169_in0
	// Insensitive connections
	assign notOp_169_in0 = state_1_is_active;
	// controller for notOp_171.notOp_171_in0
	// Insensitive connections
	assign notOp_171_in0 = state_2_is_active;
	// controller for notOp_173.notOp_173_in0
	// Insensitive connections
	assign notOp_173_in0 = state_3_is_active;
	// controller for notOp_175.notOp_175_in0
	// Insensitive connections
	assign notOp_175_in0 = state_4_is_active;
	// controller for notOp_177.notOp_177_in0
	// Insensitive connections
	assign notOp_177_in0 = state_5_is_active;
	// controller for notOp_182.notOp_182_in0
	// Insensitive connections
	assign notOp_182_in0 = andOp_100_out;
	// controller for notOp_184.notOp_184_in0
	// Insensitive connections
	assign notOp_184_in0 = andOp_62_out;
	// controller for notOp_186.notOp_186_in0
	// Insensitive connections
	assign notOp_186_in0 = andOp_68_out;
	// controller for notOp_188.notOp_188_in0
	// Insensitive connections
	assign notOp_188_in0 = andOp_151_out;
	// controller for notOp_190.notOp_190_in0
	// Insensitive connections
	assign notOp_190_in0 = andOp_152_out;
	// controller for notOp_192.notOp_192_in0
	// Insensitive connections
	assign notOp_192_in0 = andOp_153_out;
	// controller for notOp_194.notOp_194_in0
	// Insensitive connections
	assign notOp_194_in0 = andOp_154_out;
	// controller for notOp_196.notOp_196_in0
	// Insensitive connections
	assign notOp_196_in0 = andOp_155_out;
	// controller for notOp_198.notOp_198_in0
	// Insensitive connections
	assign notOp_198_in0 = andOp_66_out;
	// controller for notOp_200.notOp_200_in0
	// Insensitive connections
	assign notOp_200_in0 = andOp_168_out;
	// controller for notOp_202.notOp_202_in0
	// Insensitive connections
	assign notOp_202_in0 = andOp_181_out;
	// controller for notOp_63.notOp_63_in0
	// Insensitive connections
	assign notOp_63_in0 = andOp_62_out;
	// controller for notOp_65.notOp_65_in0
	// Insensitive connections
	assign notOp_65_in0 = andOp_64_out;
	// controller for notOp_67.notOp_67_in0
	// Insensitive connections
	assign notOp_67_in0 = icmp_icmp5_out;
	// controller for notOp_70.notOp_70_in0
	// Insensitive connections
	assign notOp_70_in0 = andOp_69_out;
	// controller for notOp_72.notOp_72_in0
	// Insensitive connections
	assign notOp_72_in0 = andOp_71_out;
	// controller for notOp_74.notOp_74_in0
	// Insensitive connections
	assign notOp_74_in0 = icmp_icmp5_out;
	// controller for notOp_77.notOp_77_in0
	// Insensitive connections
	assign notOp_77_in0 = andOp_76_out;
	// controller for notOp_79.notOp_79_in0
	// Insensitive connections
	assign notOp_79_in0 = icmp_icmp5_out;
	// controller for notOp_82.notOp_82_in0
	// Insensitive connections
	assign notOp_82_in0 = andOp_81_out;
	// controller for notOp_84.notOp_84_in0
	// Insensitive connections
	assign notOp_84_in0 = icmp_icmp5_out;
	// controller for notOp_87.notOp_87_in0
	// Insensitive connections
	assign notOp_87_in0 = andOp_86_out;
	// controller for notOp_89.notOp_89_in0
	// Insensitive connections
	assign notOp_89_in0 = icmp_icmp5_out;
	// controller for notOp_92.notOp_92_in0
	// Insensitive connections
	assign notOp_92_in0 = andOp_91_out;
	// controller for notOp_94.notOp_94_in0
	// Insensitive connections
	assign notOp_94_in0 = icmp_icmp5_out;
	// controller for notOp_97.notOp_97_in0
	// Insensitive connections
	assign notOp_97_in0 = andOp_96_out;
	// controller for notOp_99.notOp_99_in0
	// Insensitive connections
	assign notOp_99_in0 = icmp_icmp18_out;
	// controller for orOp_103.orOp_103_in0
	// controller for orOp_103.orOp_103_in1
	// Insensitive connections
	assign orOp_103_in0 = eq_102_out;
	assign orOp_103_in1 = andOp_69_out;
	// controller for orOp_111.orOp_111_in0
	// controller for orOp_111.orOp_111_in1
	// Insensitive connections
	assign orOp_111_in0 = eq_110_out;
	assign orOp_111_in1 = andOp_66_out;
	// controller for orOp_204.orOp_204_in0
	// controller for orOp_204.orOp_204_in1
	// Insensitive connections
	assign orOp_204_in0 = state_1_is_active;
	assign orOp_204_in1 = 1'd0;
	// controller for orOp_205.orOp_205_in0
	// controller for orOp_205.orOp_205_in1
	// Insensitive connections
	assign orOp_205_in0 = state_2_is_active;
	assign orOp_205_in1 = orOp_204_out;
	// controller for orOp_206.orOp_206_in0
	// controller for orOp_206.orOp_206_in1
	// Insensitive connections
	assign orOp_206_in0 = state_3_is_active;
	assign orOp_206_in1 = orOp_205_out;
	// controller for orOp_207.orOp_207_in0
	// controller for orOp_207.orOp_207_in1
	// Insensitive connections
	assign orOp_207_in0 = state_4_is_active;
	assign orOp_207_in1 = orOp_206_out;
	// controller for orOp_208.orOp_208_in0
	// controller for orOp_208.orOp_208_in1
	// Insensitive connections
	assign orOp_208_in0 = state_5_is_active;
	assign orOp_208_in1 = orOp_207_out;
	// controller for orOp_209.orOp_209_in0
	// controller for orOp_209.orOp_209_in1
	// Insensitive connections
	assign orOp_209_in0 = state_6_is_active;
	assign orOp_209_in1 = orOp_208_out;
	// controller for phi_phi2.phi_phi2_in
	// controller for phi_phi2.phi_phi2_last_block
	// controller for phi_phi2.phi_phi2_s
	// Insensitive connections
	assign phi_phi2_in = concat_128_out;
	assign phi_phi2_last_block = bb_4_predecessor_in_state_1_out_data;
	assign phi_phi2_s = concat_129_out;
	// controller for phi_phi7.phi_phi7_in
	// controller for phi_phi7.phi_phi7_last_block
	// controller for phi_phi7.phi_phi7_s
	// Insensitive connections
	assign phi_phi7_in = concat_137_out;
	assign phi_phi7_last_block = bb_1_predecessor_in_state_1_out_data;
	assign phi_phi7_s = concat_138_out;
	// controller for ret20.valid_reg
	always @(*) begin
		if (andOp_150_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// controller for shl_shl8.shl_shl8_in0
	// controller for shl_shl8.shl_shl8_in1
	// Insensitive connections
	assign shl_shl8_in0 = phi_phi7_out;
	assign shl_shl8_in1 = 32'd4;
	// controller for tmp_output_131.tmp_output_131_in_data
	always @(*) begin
		if (eq_132_out) begin 
			tmp_output_131_in_data = data_in_1_16_out_data;
		end else if (eq_133_out) begin 
			tmp_output_131_in_data = shl_shl8_out;
		end else begin
			tmp_output_131_in_data = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			data_store_0_0 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_0 <= data_in_0_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_2 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_2 <= data_in_0_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_4 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_4 <= data_in_0_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_6 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_6 <= data_in_0_7_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_10 <= 0;
		end else begin
			if (andOp_214_out) begin
				data_store_1_10 <= add_add3_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_11 <= 0;
		end else begin
			if (andOp_215_out) begin
				data_store_1_11 <= add_add4_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_13 <= 0;
		end else begin
			if (andOp_216_out) begin
				data_store_1_13 <= phi_phi7_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_15 <= 0;
		end else begin
			if (andOp_217_out) begin
				data_store_1_15 <= shl_shl8_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_8 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_8 <= data_in_1_9_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_17 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_17 <= data_in_2_18_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_19 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_19 <= data_in_2_20_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_21 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_21 <= data_in_2_22_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_23 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_23 <= data_in_2_24_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_25 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_25 <= data_in_2_26_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_27 <= 0;
		end else begin
			if (andOp_220_out) begin
				data_store_2_27 <= a_rdata_0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_28 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_28 <= data_in_3_29_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_31 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_31 <= data_in_3_32_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_33 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_33 <= data_in_3_34_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_35 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_35 <= data_in_3_36_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_38 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_38 <= data_in_4_39_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_40 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_40 <= data_in_4_41_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_42 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_42 <= data_in_4_43_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_44 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_44 <= data_in_4_45_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_46 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_46 <= data_in_5_47_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_48 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_48 <= data_in_5_49_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_50 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_50 <= data_in_5_51_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_52 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_52 <= data_in_5_53_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_54 <= 0;
		end else begin
			if (andOp_230_out) begin
				data_store_6_54 <= add_add17_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_56 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_56 <= data_in_6_57_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_58 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_58 <= data_in_6_59_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_60 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_60 <= data_in_6_61_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_167_out) begin
				global_state <= 32'd7;
			end
			if (andOp_181_out) begin
				global_state <= 32'd7;
			end
			if (andOp_62_out) begin
				global_state <= 32'd200000;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			out_of_pipe_6_7 <= 0;
		end else begin
			if (andOp_98_out) begin
				out_of_pipe_6_7 <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			out_of_pipe_bb_6_7 <= 0;
		end else begin
			if (andOp_98_out) begin
				out_of_pipe_bb_6_7 <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (1'd1) begin
				state_0_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_100_out) begin
				state_1_entry_BB_reg <= 32'd1;
			end
			if (andOp_62_out) begin
				state_1_entry_BB_reg <= 32'd1;
			end
			if (andOp_68_out) begin
				state_1_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_100_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_187_out) begin
				state_1_is_active <= 1'd0;
			end
			if (andOp_62_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_68_out) begin
				state_1_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_100_out) begin
				state_1_last_BB_reg <= 32'd3;
			end
			if (andOp_62_out) begin
				state_1_last_BB_reg <= 32'd0;
			end
			if (andOp_68_out) begin
				state_1_last_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_100_out) begin
				state_1_last_state <= 32'd6;
			end
			if (andOp_62_out) begin
				state_1_last_state <= 32'd0;
			end
			if (andOp_68_out) begin
				state_1_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_151_out) begin
				state_2_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_151_out) begin
				state_2_is_active <= 1'd1;
			end
			if (andOp_189_out) begin
				state_2_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_151_out) begin
				state_2_last_BB_reg <= bb_4_predecessor_in_state_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_151_out) begin
				state_2_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_152_out) begin
				state_3_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_152_out) begin
				state_3_is_active <= 1'd1;
			end
			if (andOp_191_out) begin
				state_3_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_152_out) begin
				state_3_last_BB_reg <= bb_4_predecessor_in_state_2_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_state <= 0;
		end else begin
			if (andOp_152_out) begin
				state_3_last_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_153_out) begin
				state_4_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_153_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_193_out) begin
				state_4_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_153_out) begin
				state_4_last_BB_reg <= bb_4_predecessor_in_state_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_state <= 0;
		end else begin
			if (andOp_153_out) begin
				state_4_last_state <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_entry_BB_reg <= 0;
		end else begin
			if (andOp_154_out) begin
				state_5_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_is_active <= 0;
		end else begin
			if (andOp_154_out) begin
				state_5_is_active <= 1'd1;
			end
			if (andOp_195_out) begin
				state_5_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_last_BB_reg <= 0;
		end else begin
			if (andOp_154_out) begin
				state_5_last_BB_reg <= bb_4_predecessor_in_state_4_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_last_state <= 0;
		end else begin
			if (andOp_154_out) begin
				state_5_last_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_entry_BB_reg <= 0;
		end else begin
			if (andOp_155_out) begin
				state_6_entry_BB_reg <= 32'd4;
			end
			if (andOp_66_out) begin
				state_6_entry_BB_reg <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_is_active <= 0;
		end else begin
			if (andOp_155_out) begin
				state_6_is_active <= 1'd1;
			end
			if (andOp_199_out) begin
				state_6_is_active <= 1'd0;
			end
			if (andOp_66_out) begin
				state_6_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_last_BB_reg <= 0;
		end else begin
			if (andOp_155_out) begin
				state_6_last_BB_reg <= bb_4_predecessor_in_state_5_out_data;
			end
			if (andOp_66_out) begin
				state_6_last_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_last_state <= 0;
		end else begin
			if (andOp_155_out) begin
				state_6_last_state <= 32'd5;
			end
			if (andOp_66_out) begin
				state_6_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_entry_BB_reg <= 0;
		end else begin
			if (andOp_180_out) begin
				state_7_entry_BB_reg <= 32'd2;
			end
			if (andOp_181_out) begin
				state_7_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_is_active <= 0;
		end else begin
			if (andOp_168_out) begin
				state_7_is_active <= 1'd1;
			end
			if (andOp_181_out) begin
				state_7_is_active <= 1'd1;
			end
			if (andOp_203_out) begin
				state_7_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_last_BB_reg <= 0;
		end else begin
			if (andOp_181_out) begin
				state_7_last_BB_reg <= bb_2_predecessor_in_state_7_out_data;
			end
			if (andOp_98_out) begin
				state_7_last_BB_reg <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_last_state <= 0;
		end else begin
			if (andOp_181_out) begin
				state_7_last_state <= 32'd7;
			end
			if (andOp_98_out) begin
				state_7_last_state <= 32'd6;
			end
		end
	end

endmodule

