module channel_reduce_4(input [0:0] clk, input [0:0] rst, output [31:0] out_in_data, output [0:0] out_read_valid, output [0:0] out_rst, output [0:0] out_write_valid, input [31:0] out_out_data, input [0:0] out_read_ready, input [0:0] out_write_ready, output [31:0] in_in_data, output [0:0] in_read_valid, output [0:0] in_rst, output [0:0] in_write_valid, input [31:0] in_out_data, input [0:0] in_read_ready, input [0:0] in_write_ready, output [0:0] valid);

	reg [31:0] out_in_data_reg;
	reg [0:0] out_read_valid_reg;
	reg [0:0] out_rst_reg;
	reg [0:0] out_write_valid_reg;
	reg [31:0] in_in_data_reg;
	reg [0:0] in_read_valid_reg;
	reg [0:0] in_rst_reg;
	reg [0:0] in_write_valid_reg;
	reg [0:0] valid_reg;

	assign out_in_data = out_in_data_reg;
	assign out_read_valid = out_read_valid_reg;
	assign out_rst = out_rst_reg;
	assign out_write_valid = out_write_valid_reg;
	assign in_in_data = in_in_data_reg;
	assign in_read_valid = in_read_valid_reg;
	assign in_rst = in_rst_reg;
	assign in_write_valid = in_write_valid_reg;
	assign valid = valid_reg;

	// Start debug wires and ports

	initial begin
	end





	// End debug wires and ports

	// Start Functional Units
	br_dummy br_unit();

	add alloca_0();

	add bitcast_1();

	add call_2();

	reg [31:0] raddr_ram_0_reg;
	reg [31:0] waddr_ram_0_reg;
	reg [31:0] wdata_ram_0_reg;
	reg [0:0] wen_ram_0_reg;
	wire [31:0] rdata_ram_0;
	register #(.WIDTH(32)) ram_0(.clk(clk), .raddr(raddr_ram_0_reg), .rdata(rdata_ram_0), .rst(rst), .waddr(waddr_ram_0_reg), .wdata(wdata_ram_0_reg), .wen(wen_ram_0_reg));

	add call_20();

	reg [63:0] phi_in_phi_8;
	reg [31:0] phi_last_block_phi_8;
	reg [63:0] phi_s_phi_8;
	wire [31:0] phi_out_phi_8;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_8(.in(phi_in_phi_8), .last_block(phi_last_block_phi_8), .out(phi_out_phi_8), .s(phi_s_phi_8));

	reg [31:0] add_in0_add_14;
	reg [31:0] add_in1_add_14;
	wire [31:0] add_out_add_14;
	add #(.WIDTH(32)) add_add_14(.in0(add_in0_add_14), .in1(add_in1_add_14), .out(add_out_add_14));

	reg [31:0] add_in0_add_16;
	reg [31:0] add_in1_add_16;
	wire [31:0] add_out_add_16;
	add #(.WIDTH(32)) add_add_16(.in0(add_in0_add_16), .in1(add_in1_add_16), .out(add_out_add_16));

	reg [31:0] cmp_in0_icmp_17;
	reg [31:0] cmp_in1_icmp_17;
	wire [0:0] cmp_out_icmp_17;
	eq #(.WIDTH(32)) icmp_17(.in0(cmp_in0_icmp_17), .in1(cmp_in1_icmp_17), .out(cmp_out_icmp_17));

	reg [31:0] data_in_0_1_in_data;
	wire [31:0] data_in_0_1_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_1(.in_data(data_in_0_1_in_data), .out_data(data_in_0_1_out_data));

	reg [31:0] data_in_0_3_in_data;
	wire [31:0] data_in_0_3_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_3(.in_data(data_in_0_3_in_data), .out_data(data_in_0_3_out_data));

	reg [0:0] data_in_0_5_in_data;
	wire [0:0] data_in_0_5_out_data;
	hls_wire #(.WIDTH(1)) data_in_0_5(.in_data(data_in_0_5_in_data), .out_data(data_in_0_5_out_data));

	reg [31:0] data_in_1_7_in_data;
	wire [31:0] data_in_1_7_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_7(.in_data(data_in_1_7_in_data), .out_data(data_in_1_7_out_data));

	reg [31:0] data_in_1_9_in_data;
	wire [31:0] data_in_1_9_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_9(.in_data(data_in_1_9_in_data), .out_data(data_in_1_9_out_data));

	reg [0:0] data_in_1_11_in_data;
	wire [0:0] data_in_1_11_out_data;
	hls_wire #(.WIDTH(1)) data_in_1_11(.in_data(data_in_1_11_in_data), .out_data(data_in_1_11_out_data));

	reg [31:0] data_in_2_13_in_data;
	wire [31:0] data_in_2_13_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_13(.in_data(data_in_2_13_in_data), .out_data(data_in_2_13_out_data));

	reg [31:0] data_in_2_15_in_data;
	wire [31:0] data_in_2_15_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_15(.in_data(data_in_2_15_in_data), .out_data(data_in_2_15_out_data));

	reg [0:0] data_in_2_17_in_data;
	wire [0:0] data_in_2_17_out_data;
	hls_wire #(.WIDTH(1)) data_in_2_17(.in_data(data_in_2_17_in_data), .out_data(data_in_2_17_out_data));

	reg [31:0] data_in_3_19_in_data;
	wire [31:0] data_in_3_19_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_19(.in_data(data_in_3_19_in_data), .out_data(data_in_3_19_out_data));

	reg [31:0] data_in_3_21_in_data;
	wire [31:0] data_in_3_21_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_21(.in_data(data_in_3_21_in_data), .out_data(data_in_3_21_out_data));

	reg [0:0] data_in_3_23_in_data;
	wire [0:0] data_in_3_23_out_data;
	hls_wire #(.WIDTH(1)) data_in_3_23(.in_data(data_in_3_23_in_data), .out_data(data_in_3_23_out_data));

	reg [31:0] data_in_4_25_in_data;
	wire [31:0] data_in_4_25_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_25(.in_data(data_in_4_25_in_data), .out_data(data_in_4_25_out_data));

	reg [31:0] data_in_4_27_in_data;
	wire [31:0] data_in_4_27_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_27(.in_data(data_in_4_27_in_data), .out_data(data_in_4_27_out_data));

	reg [0:0] data_in_4_29_in_data;
	wire [0:0] data_in_4_29_out_data;
	hls_wire #(.WIDTH(1)) data_in_4_29(.in_data(data_in_4_29_in_data), .out_data(data_in_4_29_out_data));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] bb_0_active_in_state_1_in_data;
	wire [0:0] bb_0_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_1(.in_data(bb_0_active_in_state_1_in_data), .out_data(bb_0_active_in_state_1_out_data));

	reg [31:0] bb_0_predecessor_in_state_1_in_data;
	wire [31:0] bb_0_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_1(.in_data(bb_0_predecessor_in_state_1_in_data), .out_data(bb_0_predecessor_in_state_1_out_data));

	reg [0:0] bb_3_active_in_state_1_in_data;
	wire [0:0] bb_3_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_1(.in_data(bb_3_active_in_state_1_in_data), .out_data(bb_3_active_in_state_1_out_data));

	reg [31:0] bb_3_predecessor_in_state_1_in_data;
	wire [31:0] bb_3_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_1(.in_data(bb_3_predecessor_in_state_1_in_data), .out_data(bb_3_predecessor_in_state_1_out_data));

	reg [0:0] bb_9_active_in_state_1_in_data;
	wire [0:0] bb_9_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_9_active_in_state_1(.in_data(bb_9_active_in_state_1_in_data), .out_data(bb_9_active_in_state_1_out_data));

	reg [31:0] bb_9_predecessor_in_state_1_in_data;
	wire [31:0] bb_9_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_9_predecessor_in_state_1(.in_data(bb_9_predecessor_in_state_1_in_data), .out_data(bb_9_predecessor_in_state_1_out_data));

	reg [0:0] bb_8_active_in_state_1_in_data;
	wire [0:0] bb_8_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active_in_state_1(.in_data(bb_8_active_in_state_1_in_data), .out_data(bb_8_active_in_state_1_out_data));

	reg [31:0] bb_8_predecessor_in_state_1_in_data;
	wire [31:0] bb_8_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor_in_state_1(.in_data(bb_8_predecessor_in_state_1_in_data), .out_data(bb_8_predecessor_in_state_1_out_data));

	reg [0:0] bb_10_active_in_state_2_in_data;
	wire [0:0] bb_10_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_2(.in_data(bb_10_active_in_state_2_in_data), .out_data(bb_10_active_in_state_2_out_data));

	reg [31:0] bb_10_predecessor_in_state_2_in_data;
	wire [31:0] bb_10_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_2(.in_data(bb_10_predecessor_in_state_2_in_data), .out_data(bb_10_predecessor_in_state_2_out_data));

	reg [0:0] bb_4_active_in_state_3_in_data;
	wire [0:0] bb_4_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_3(.in_data(bb_4_active_in_state_3_in_data), .out_data(bb_4_active_in_state_3_out_data));

	reg [31:0] bb_4_predecessor_in_state_3_in_data;
	wire [31:0] bb_4_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_3(.in_data(bb_4_predecessor_in_state_3_in_data), .out_data(bb_4_predecessor_in_state_3_out_data));

	reg [0:0] bb_10_active_in_state_3_in_data;
	wire [0:0] bb_10_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_3(.in_data(bb_10_active_in_state_3_in_data), .out_data(bb_10_active_in_state_3_out_data));

	reg [31:0] bb_10_predecessor_in_state_3_in_data;
	wire [31:0] bb_10_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_3(.in_data(bb_10_predecessor_in_state_3_in_data), .out_data(bb_10_predecessor_in_state_3_out_data));

	reg [0:0] bb_5_active_in_state_4_in_data;
	wire [0:0] bb_5_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_5_active_in_state_4(.in_data(bb_5_active_in_state_4_in_data), .out_data(bb_5_active_in_state_4_out_data));

	reg [31:0] bb_5_predecessor_in_state_4_in_data;
	wire [31:0] bb_5_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_5_predecessor_in_state_4(.in_data(bb_5_predecessor_in_state_4_in_data), .out_data(bb_5_predecessor_in_state_4_out_data));

	reg [0:0] bb_6_active_in_state_4_in_data;
	wire [0:0] bb_6_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_6_active_in_state_4(.in_data(bb_6_active_in_state_4_in_data), .out_data(bb_6_active_in_state_4_out_data));

	reg [31:0] bb_6_predecessor_in_state_4_in_data;
	wire [31:0] bb_6_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_6_predecessor_in_state_4(.in_data(bb_6_predecessor_in_state_4_in_data), .out_data(bb_6_predecessor_in_state_4_out_data));

	reg [0:0] bb_7_active_in_state_4_in_data;
	wire [0:0] bb_7_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_7_active_in_state_4(.in_data(bb_7_active_in_state_4_in_data), .out_data(bb_7_active_in_state_4_out_data));

	reg [31:0] bb_7_predecessor_in_state_4_in_data;
	wire [31:0] bb_7_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_7_predecessor_in_state_4(.in_data(bb_7_predecessor_in_state_4_in_data), .out_data(bb_7_predecessor_in_state_4_out_data));

	reg [0:0] bb_2_active_in_state_4_in_data;
	wire [0:0] bb_2_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_4(.in_data(bb_2_active_in_state_4_in_data), .out_data(bb_2_active_in_state_4_out_data));

	reg [31:0] bb_2_predecessor_in_state_4_in_data;
	wire [31:0] bb_2_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_4(.in_data(bb_2_predecessor_in_state_4_in_data), .out_data(bb_2_predecessor_in_state_4_out_data));

	reg [0:0] bb_1_active_in_state_4_in_data;
	wire [0:0] bb_1_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_4(.in_data(bb_1_active_in_state_4_in_data), .out_data(bb_1_active_in_state_4_out_data));

	reg [31:0] bb_1_predecessor_in_state_4_in_data;
	wire [31:0] bb_1_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_4(.in_data(bb_1_predecessor_in_state_4_in_data), .out_data(bb_1_predecessor_in_state_4_out_data));

	reg [0:0] bb_4_active_in_state_4_in_data;
	wire [0:0] bb_4_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_4(.in_data(bb_4_active_in_state_4_in_data), .out_data(bb_4_active_in_state_4_out_data));

	reg [31:0] bb_4_predecessor_in_state_4_in_data;
	wire [31:0] bb_4_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_4(.in_data(bb_4_predecessor_in_state_4_in_data), .out_data(bb_4_predecessor_in_state_4_out_data));

	reg [0:0] andOp_30_in0;
	reg [0:0] andOp_30_in1;
	wire [0:0] andOp_30_out;
	andOp #(.WIDTH(1)) andOp_30(.in0(andOp_30_in0), .in1(andOp_30_in1), .out(andOp_30_out));

	reg [0:0] andOp_31_in0;
	reg [0:0] andOp_31_in1;
	wire [0:0] andOp_31_out;
	andOp #(.WIDTH(1)) andOp_31(.in0(andOp_31_in0), .in1(andOp_31_in1), .out(andOp_31_out));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] notOp_32_in0;
	wire [0:0] notOp_32_out;
	notOp #(.WIDTH(1)) notOp_32(.in(notOp_32_in0), .out(notOp_32_out));

	reg [0:0] andOp_33_in0;
	reg [0:0] andOp_33_in1;
	wire [0:0] andOp_33_out;
	andOp #(.WIDTH(1)) andOp_33(.in0(andOp_33_in0), .in1(andOp_33_in1), .out(andOp_33_out));

	reg [0:0] andOp_34_in0;
	reg [0:0] andOp_34_in1;
	wire [0:0] andOp_34_out;
	andOp #(.WIDTH(1)) andOp_34(.in0(andOp_34_in0), .in1(andOp_34_in1), .out(andOp_34_out));

	reg [0:0] br_0_happened_in_state_1_in_data;
	wire [0:0] br_0_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_1(.in_data(br_0_happened_in_state_1_in_data), .out_data(br_0_happened_in_state_1_out_data));

	reg [0:0] notOp_35_in0;
	wire [0:0] notOp_35_out;
	notOp #(.WIDTH(1)) notOp_35(.in(notOp_35_in0), .out(notOp_35_out));

	reg [0:0] andOp_36_in0;
	reg [0:0] andOp_36_in1;
	wire [0:0] andOp_36_out;
	andOp #(.WIDTH(1)) andOp_36(.in0(andOp_36_in0), .in1(andOp_36_in1), .out(andOp_36_out));

	reg [0:0] andOp_37_in0;
	reg [0:0] andOp_37_in1;
	wire [0:0] andOp_37_out;
	andOp #(.WIDTH(1)) andOp_37(.in0(andOp_37_in0), .in1(andOp_37_in1), .out(andOp_37_out));

	reg [0:0] br_3_happened_in_state_1_in_data;
	wire [0:0] br_3_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_1(.in_data(br_3_happened_in_state_1_in_data), .out_data(br_3_happened_in_state_1_out_data));

	reg [0:0] notOp_38_in0;
	wire [0:0] notOp_38_out;
	notOp #(.WIDTH(1)) notOp_38(.in(notOp_38_in0), .out(notOp_38_out));

	reg [0:0] andOp_39_in0;
	reg [0:0] andOp_39_in1;
	wire [0:0] andOp_39_out;
	andOp #(.WIDTH(1)) andOp_39(.in0(andOp_39_in0), .in1(andOp_39_in1), .out(andOp_39_out));

	reg [0:0] andOp_40_in0;
	reg [0:0] andOp_40_in1;
	wire [0:0] andOp_40_out;
	andOp #(.WIDTH(1)) andOp_40(.in0(andOp_40_in0), .in1(andOp_40_in1), .out(andOp_40_out));

	reg [0:0] br_9_happened_in_state_1_in_data;
	wire [0:0] br_9_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_9_happened_in_state_1(.in_data(br_9_happened_in_state_1_in_data), .out_data(br_9_happened_in_state_1_out_data));

	reg [0:0] notOp_41_in0;
	wire [0:0] notOp_41_out;
	notOp #(.WIDTH(1)) notOp_41(.in(notOp_41_in0), .out(notOp_41_out));

	reg [0:0] andOp_42_in0;
	reg [0:0] andOp_42_in1;
	wire [0:0] andOp_42_out;
	andOp #(.WIDTH(1)) andOp_42(.in0(andOp_42_in0), .in1(andOp_42_in1), .out(andOp_42_out));

	reg [0:0] notOp_43_in0;
	wire [0:0] notOp_43_out;
	notOp #(.WIDTH(1)) notOp_43(.in(notOp_43_in0), .out(notOp_43_out));

	reg [0:0] andOp_44_in0;
	reg [0:0] andOp_44_in1;
	wire [0:0] andOp_44_out;
	andOp #(.WIDTH(1)) andOp_44(.in0(andOp_44_in0), .in1(andOp_44_in1), .out(andOp_44_out));

	reg [0:0] andOp_45_in0;
	reg [0:0] andOp_45_in1;
	wire [0:0] andOp_45_out;
	andOp #(.WIDTH(1)) andOp_45(.in0(andOp_45_in0), .in1(andOp_45_in1), .out(andOp_45_out));

	reg [0:0] andOp_46_in0;
	reg [0:0] andOp_46_in1;
	wire [0:0] andOp_46_out;
	andOp #(.WIDTH(1)) andOp_46(.in0(andOp_46_in0), .in1(andOp_46_in1), .out(andOp_46_out));

	reg [0:0] br_8_happened_in_state_1_in_data;
	wire [0:0] br_8_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_8_happened_in_state_1(.in_data(br_8_happened_in_state_1_in_data), .out_data(br_8_happened_in_state_1_out_data));

	reg [0:0] notOp_47_in0;
	wire [0:0] notOp_47_out;
	notOp #(.WIDTH(1)) notOp_47(.in(notOp_47_in0), .out(notOp_47_out));

	reg [0:0] andOp_48_in0;
	reg [0:0] andOp_48_in1;
	wire [0:0] andOp_48_out;
	andOp #(.WIDTH(1)) andOp_48(.in0(andOp_48_in0), .in1(andOp_48_in1), .out(andOp_48_out));

	reg [0:0] andOp_49_in0;
	reg [0:0] andOp_49_in1;
	wire [0:0] andOp_49_out;
	andOp #(.WIDTH(1)) andOp_49(.in0(andOp_49_in0), .in1(andOp_49_in1), .out(andOp_49_out));

	reg [0:0] br_10_happened_in_state_2_in_data;
	wire [0:0] br_10_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_2(.in_data(br_10_happened_in_state_2_in_data), .out_data(br_10_happened_in_state_2_out_data));

	reg [0:0] notOp_50_in0;
	wire [0:0] notOp_50_out;
	notOp #(.WIDTH(1)) notOp_50(.in(notOp_50_in0), .out(notOp_50_out));

	reg [0:0] andOp_51_in0;
	reg [0:0] andOp_51_in1;
	wire [0:0] andOp_51_out;
	andOp #(.WIDTH(1)) andOp_51(.in0(andOp_51_in0), .in1(andOp_51_in1), .out(andOp_51_out));

	reg [0:0] andOp_52_in0;
	reg [0:0] andOp_52_in1;
	wire [0:0] andOp_52_out;
	andOp #(.WIDTH(1)) andOp_52(.in0(andOp_52_in0), .in1(andOp_52_in1), .out(andOp_52_out));

	reg [0:0] br_4_happened_in_state_3_in_data;
	wire [0:0] br_4_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_3(.in_data(br_4_happened_in_state_3_in_data), .out_data(br_4_happened_in_state_3_out_data));

	reg [0:0] notOp_53_in0;
	wire [0:0] notOp_53_out;
	notOp #(.WIDTH(1)) notOp_53(.in(notOp_53_in0), .out(notOp_53_out));

	reg [0:0] andOp_54_in0;
	reg [0:0] andOp_54_in1;
	wire [0:0] andOp_54_out;
	andOp #(.WIDTH(1)) andOp_54(.in0(andOp_54_in0), .in1(andOp_54_in1), .out(andOp_54_out));

	reg [0:0] notOp_55_in0;
	wire [0:0] notOp_55_out;
	notOp #(.WIDTH(1)) notOp_55(.in(notOp_55_in0), .out(notOp_55_out));

	reg [0:0] andOp_56_in0;
	reg [0:0] andOp_56_in1;
	wire [0:0] andOp_56_out;
	andOp #(.WIDTH(1)) andOp_56(.in0(andOp_56_in0), .in1(andOp_56_in1), .out(andOp_56_out));

	reg [0:0] andOp_57_in0;
	reg [0:0] andOp_57_in1;
	wire [0:0] andOp_57_out;
	andOp #(.WIDTH(1)) andOp_57(.in0(andOp_57_in0), .in1(andOp_57_in1), .out(andOp_57_out));

	reg [0:0] andOp_58_in0;
	reg [0:0] andOp_58_in1;
	wire [0:0] andOp_58_out;
	andOp #(.WIDTH(1)) andOp_58(.in0(andOp_58_in0), .in1(andOp_58_in1), .out(andOp_58_out));

	reg [0:0] br_10_happened_in_state_3_in_data;
	wire [0:0] br_10_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_3(.in_data(br_10_happened_in_state_3_in_data), .out_data(br_10_happened_in_state_3_out_data));

	reg [0:0] notOp_59_in0;
	wire [0:0] notOp_59_out;
	notOp #(.WIDTH(1)) notOp_59(.in(notOp_59_in0), .out(notOp_59_out));

	reg [0:0] andOp_60_in0;
	reg [0:0] andOp_60_in1;
	wire [0:0] andOp_60_out;
	andOp #(.WIDTH(1)) andOp_60(.in0(andOp_60_in0), .in1(andOp_60_in1), .out(andOp_60_out));

	reg [0:0] andOp_61_in0;
	reg [0:0] andOp_61_in1;
	wire [0:0] andOp_61_out;
	andOp #(.WIDTH(1)) andOp_61(.in0(andOp_61_in0), .in1(andOp_61_in1), .out(andOp_61_out));

	reg [0:0] br_5_happened_in_state_4_in_data;
	wire [0:0] br_5_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_5_happened_in_state_4(.in_data(br_5_happened_in_state_4_in_data), .out_data(br_5_happened_in_state_4_out_data));

	reg [0:0] notOp_62_in0;
	wire [0:0] notOp_62_out;
	notOp #(.WIDTH(1)) notOp_62(.in(notOp_62_in0), .out(notOp_62_out));

	reg [0:0] andOp_63_in0;
	reg [0:0] andOp_63_in1;
	wire [0:0] andOp_63_out;
	andOp #(.WIDTH(1)) andOp_63(.in0(andOp_63_in0), .in1(andOp_63_in1), .out(andOp_63_out));

	reg [0:0] andOp_64_in0;
	reg [0:0] andOp_64_in1;
	wire [0:0] andOp_64_out;
	andOp #(.WIDTH(1)) andOp_64(.in0(andOp_64_in0), .in1(andOp_64_in1), .out(andOp_64_out));

	reg [0:0] br_6_happened_in_state_4_in_data;
	wire [0:0] br_6_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_6_happened_in_state_4(.in_data(br_6_happened_in_state_4_in_data), .out_data(br_6_happened_in_state_4_out_data));

	reg [0:0] notOp_65_in0;
	wire [0:0] notOp_65_out;
	notOp #(.WIDTH(1)) notOp_65(.in(notOp_65_in0), .out(notOp_65_out));

	reg [0:0] andOp_66_in0;
	reg [0:0] andOp_66_in1;
	wire [0:0] andOp_66_out;
	andOp #(.WIDTH(1)) andOp_66(.in0(andOp_66_in0), .in1(andOp_66_in1), .out(andOp_66_out));

	reg [0:0] notOp_67_in0;
	wire [0:0] notOp_67_out;
	notOp #(.WIDTH(1)) notOp_67(.in(notOp_67_in0), .out(notOp_67_out));

	reg [0:0] andOp_68_in0;
	reg [0:0] andOp_68_in1;
	wire [0:0] andOp_68_out;
	andOp #(.WIDTH(1)) andOp_68(.in0(andOp_68_in0), .in1(andOp_68_in1), .out(andOp_68_out));

	reg [0:0] andOp_69_in0;
	reg [0:0] andOp_69_in1;
	wire [0:0] andOp_69_out;
	andOp #(.WIDTH(1)) andOp_69(.in0(andOp_69_in0), .in1(andOp_69_in1), .out(andOp_69_out));

	reg [0:0] andOp_70_in0;
	reg [0:0] andOp_70_in1;
	wire [0:0] andOp_70_out;
	andOp #(.WIDTH(1)) andOp_70(.in0(andOp_70_in0), .in1(andOp_70_in1), .out(andOp_70_out));

	reg [0:0] br_7_happened_in_state_4_in_data;
	wire [0:0] br_7_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_7_happened_in_state_4(.in_data(br_7_happened_in_state_4_in_data), .out_data(br_7_happened_in_state_4_out_data));

	reg [0:0] notOp_71_in0;
	wire [0:0] notOp_71_out;
	notOp #(.WIDTH(1)) notOp_71(.in(notOp_71_in0), .out(notOp_71_out));

	reg [0:0] andOp_72_in0;
	reg [0:0] andOp_72_in1;
	wire [0:0] andOp_72_out;
	andOp #(.WIDTH(1)) andOp_72(.in0(andOp_72_in0), .in1(andOp_72_in1), .out(andOp_72_out));

	reg [0:0] andOp_73_in0;
	reg [0:0] andOp_73_in1;
	wire [0:0] andOp_73_out;
	andOp #(.WIDTH(1)) andOp_73(.in0(andOp_73_in0), .in1(andOp_73_in1), .out(andOp_73_out));

	reg [0:0] br_1_happened_in_state_4_in_data;
	wire [0:0] br_1_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened_in_state_4(.in_data(br_1_happened_in_state_4_in_data), .out_data(br_1_happened_in_state_4_out_data));

	reg [0:0] notOp_74_in0;
	wire [0:0] notOp_74_out;
	notOp #(.WIDTH(1)) notOp_74(.in(notOp_74_in0), .out(notOp_74_out));

	reg [0:0] andOp_75_in0;
	reg [0:0] andOp_75_in1;
	wire [0:0] andOp_75_out;
	andOp #(.WIDTH(1)) andOp_75(.in0(andOp_75_in0), .in1(andOp_75_in1), .out(andOp_75_out));

	reg [0:0] andOp_76_in0;
	reg [0:0] andOp_76_in1;
	wire [0:0] andOp_76_out;
	andOp #(.WIDTH(1)) andOp_76(.in0(andOp_76_in0), .in1(andOp_76_in1), .out(andOp_76_out));

	reg [0:0] br_4_happened_in_state_4_in_data;
	wire [0:0] br_4_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_4(.in_data(br_4_happened_in_state_4_in_data), .out_data(br_4_happened_in_state_4_out_data));

	reg [0:0] notOp_77_in0;
	wire [0:0] notOp_77_out;
	notOp #(.WIDTH(1)) notOp_77(.in(notOp_77_in0), .out(notOp_77_out));

	reg [0:0] andOp_78_in0;
	reg [0:0] andOp_78_in1;
	wire [0:0] andOp_78_out;
	andOp #(.WIDTH(1)) andOp_78(.in0(andOp_78_in0), .in1(andOp_78_in1), .out(andOp_78_out));

	reg [0:0] notOp_79_in0;
	wire [0:0] notOp_79_out;
	notOp #(.WIDTH(1)) notOp_79(.in(notOp_79_in0), .out(notOp_79_out));

	reg [0:0] andOp_80_in0;
	reg [0:0] andOp_80_in1;
	wire [0:0] andOp_80_out;
	andOp #(.WIDTH(1)) andOp_80(.in0(andOp_80_in0), .in1(andOp_80_in1), .out(andOp_80_out));

	reg [31:0] eq_81_in0;
	reg [31:0] eq_81_in1;
	wire [0:0] eq_81_out;
	eq #(.WIDTH(32)) eq_81(.in0(eq_81_in0), .in1(eq_81_in1), .out(eq_81_out));

	reg [31:0] eq_82_in0;
	reg [31:0] eq_82_in1;
	wire [0:0] eq_82_out;
	eq #(.WIDTH(32)) eq_82(.in0(eq_82_in0), .in1(eq_82_in1), .out(eq_82_out));

	reg [31:0] eq_83_in0;
	reg [31:0] eq_83_in1;
	wire [0:0] eq_83_out;
	eq #(.WIDTH(32)) eq_83(.in0(eq_83_in0), .in1(eq_83_in1), .out(eq_83_out));

	reg [0:0] orOp_84_in0;
	reg [0:0] orOp_84_in1;
	wire [0:0] orOp_84_out;
	orOp #(.WIDTH(1)) orOp_84(.in0(orOp_84_in0), .in1(orOp_84_in1), .out(orOp_84_out));

	reg [31:0] eq_85_in0;
	reg [31:0] eq_85_in1;
	wire [0:0] eq_85_out;
	eq #(.WIDTH(32)) eq_85(.in0(eq_85_in0), .in1(eq_85_in1), .out(eq_85_out));

	reg [0:0] orOp_86_in0;
	reg [0:0] orOp_86_in1;
	wire [0:0] orOp_86_out;
	orOp #(.WIDTH(1)) orOp_86(.in0(orOp_86_in0), .in1(orOp_86_in1), .out(orOp_86_out));

	reg [31:0] eq_87_in0;
	reg [31:0] eq_87_in1;
	wire [0:0] eq_87_out;
	eq #(.WIDTH(32)) eq_87(.in0(eq_87_in0), .in1(eq_87_in1), .out(eq_87_out));

	reg [0:0] orOp_88_in0;
	reg [0:0] orOp_88_in1;
	wire [0:0] orOp_88_out;
	orOp #(.WIDTH(1)) orOp_88(.in0(orOp_88_in0), .in1(orOp_88_in1), .out(orOp_88_out));

	reg [31:0] eq_89_in0;
	reg [31:0] eq_89_in1;
	wire [0:0] eq_89_out;
	eq #(.WIDTH(32)) eq_89(.in0(eq_89_in0), .in1(eq_89_in1), .out(eq_89_out));

	reg [31:0] eq_90_in0;
	reg [31:0] eq_90_in1;
	wire [0:0] eq_90_out;
	eq #(.WIDTH(32)) eq_90(.in0(eq_90_in0), .in1(eq_90_in1), .out(eq_90_out));

	reg [0:0] orOp_91_in0;
	reg [0:0] orOp_91_in1;
	wire [0:0] orOp_91_out;
	orOp #(.WIDTH(1)) orOp_91(.in0(orOp_91_in0), .in1(orOp_91_in1), .out(orOp_91_out));

	reg [31:0] eq_92_in0;
	reg [31:0] eq_92_in1;
	wire [0:0] eq_92_out;
	eq #(.WIDTH(32)) eq_92(.in0(eq_92_in0), .in1(eq_92_in1), .out(eq_92_out));

	reg [31:0] eq_93_in0;
	reg [31:0] eq_93_in1;
	wire [0:0] eq_93_out;
	eq #(.WIDTH(32)) eq_93(.in0(eq_93_in0), .in1(eq_93_in1), .out(eq_93_out));

	reg [0:0] orOp_94_in0;
	reg [0:0] orOp_94_in1;
	wire [0:0] orOp_94_out;
	orOp #(.WIDTH(1)) orOp_94(.in0(orOp_94_in0), .in1(orOp_94_in1), .out(orOp_94_out));

	reg [31:0] eq_95_in0;
	reg [31:0] eq_95_in1;
	wire [0:0] eq_95_out;
	eq #(.WIDTH(32)) eq_95(.in0(eq_95_in0), .in1(eq_95_in1), .out(eq_95_out));

	reg [0:0] orOp_96_in0;
	reg [0:0] orOp_96_in1;
	wire [0:0] orOp_96_out;
	orOp #(.WIDTH(1)) orOp_96(.in0(orOp_96_in0), .in1(orOp_96_in1), .out(orOp_96_out));

	reg [31:0] eq_97_in0;
	reg [31:0] eq_97_in1;
	wire [0:0] eq_97_out;
	eq #(.WIDTH(32)) eq_97(.in0(eq_97_in0), .in1(eq_97_in1), .out(eq_97_out));

	reg [0:0] orOp_98_in0;
	reg [0:0] orOp_98_in1;
	wire [0:0] orOp_98_out;
	orOp #(.WIDTH(1)) orOp_98(.in0(orOp_98_in0), .in1(orOp_98_in1), .out(orOp_98_out));

	reg [31:0] eq_99_in0;
	reg [31:0] eq_99_in1;
	wire [0:0] eq_99_out;
	eq #(.WIDTH(32)) eq_99(.in0(eq_99_in0), .in1(eq_99_in1), .out(eq_99_out));

	reg [0:0] orOp_100_in0;
	reg [0:0] orOp_100_in1;
	wire [0:0] orOp_100_out;
	orOp #(.WIDTH(1)) orOp_100(.in0(orOp_100_in0), .in1(orOp_100_in1), .out(orOp_100_out));

	reg [31:0] eq_101_in0;
	reg [31:0] eq_101_in1;
	wire [0:0] eq_101_out;
	eq #(.WIDTH(32)) eq_101(.in0(eq_101_in0), .in1(eq_101_in1), .out(eq_101_out));

	reg [0:0] orOp_102_in0;
	reg [0:0] orOp_102_in1;
	wire [0:0] orOp_102_out;
	orOp #(.WIDTH(1)) orOp_102(.in0(orOp_102_in0), .in1(orOp_102_in1), .out(orOp_102_out));

	reg [31:0] eq_103_in0;
	reg [31:0] eq_103_in1;
	wire [0:0] eq_103_out;
	eq #(.WIDTH(32)) eq_103(.in0(eq_103_in0), .in1(eq_103_in1), .out(eq_103_out));

	reg [31:0] eq_104_in0;
	reg [31:0] eq_104_in1;
	wire [0:0] eq_104_out;
	eq #(.WIDTH(32)) eq_104(.in0(eq_104_in0), .in1(eq_104_in1), .out(eq_104_out));

	reg [31:0] eq_105_in0;
	reg [31:0] eq_105_in1;
	wire [0:0] eq_105_out;
	eq #(.WIDTH(32)) eq_105(.in0(eq_105_in0), .in1(eq_105_in1), .out(eq_105_out));

	reg [31:0] eq_106_in0;
	reg [31:0] eq_106_in1;
	wire [0:0] eq_106_out;
	eq #(.WIDTH(32)) eq_106(.in0(eq_106_in0), .in1(eq_106_in1), .out(eq_106_out));

	reg [0:0] notOp_107_in0;
	wire [0:0] notOp_107_out;
	notOp #(.WIDTH(1)) notOp_107(.in(notOp_107_in0), .out(notOp_107_out));

	reg [0:0] andOp_108_in0;
	reg [0:0] andOp_108_in1;
	wire [0:0] andOp_108_out;
	andOp #(.WIDTH(1)) andOp_108(.in0(andOp_108_in0), .in1(andOp_108_in1), .out(andOp_108_out));

	reg [31:0] eq_109_in0;
	reg [31:0] eq_109_in1;
	wire [0:0] eq_109_out;
	eq #(.WIDTH(32)) eq_109(.in0(eq_109_in0), .in1(eq_109_in1), .out(eq_109_out));

	reg [0:0] notOp_110_in0;
	wire [0:0] notOp_110_out;
	notOp #(.WIDTH(1)) notOp_110(.in(notOp_110_in0), .out(notOp_110_out));

	reg [0:0] andOp_111_in0;
	reg [0:0] andOp_111_in1;
	wire [0:0] andOp_111_out;
	andOp #(.WIDTH(1)) andOp_111(.in0(andOp_111_in0), .in1(andOp_111_in1), .out(andOp_111_out));

	reg [31:0] eq_112_in0;
	reg [31:0] eq_112_in1;
	wire [0:0] eq_112_out;
	eq #(.WIDTH(32)) eq_112(.in0(eq_112_in0), .in1(eq_112_in1), .out(eq_112_out));

	reg [0:0] notOp_113_in0;
	wire [0:0] notOp_113_out;
	notOp #(.WIDTH(1)) notOp_113(.in(notOp_113_in0), .out(notOp_113_out));

	reg [0:0] andOp_114_in0;
	reg [0:0] andOp_114_in1;
	wire [0:0] andOp_114_out;
	andOp #(.WIDTH(1)) andOp_114(.in0(andOp_114_in0), .in1(andOp_114_in1), .out(andOp_114_out));

	reg [31:0] eq_115_in0;
	reg [31:0] eq_115_in1;
	wire [0:0] eq_115_out;
	eq #(.WIDTH(32)) eq_115(.in0(eq_115_in0), .in1(eq_115_in1), .out(eq_115_out));

	reg [31:0] eq_116_in0;
	reg [31:0] eq_116_in1;
	wire [0:0] eq_116_out;
	eq #(.WIDTH(32)) eq_116(.in0(eq_116_in0), .in1(eq_116_in1), .out(eq_116_out));

	reg [0:0] notOp_117_in0;
	wire [0:0] notOp_117_out;
	notOp #(.WIDTH(1)) notOp_117(.in(notOp_117_in0), .out(notOp_117_out));

	reg [0:0] andOp_118_in0;
	reg [0:0] andOp_118_in1;
	wire [0:0] andOp_118_out;
	andOp #(.WIDTH(1)) andOp_118(.in0(andOp_118_in0), .in1(andOp_118_in1), .out(andOp_118_out));

	reg [31:0] eq_119_in0;
	reg [31:0] eq_119_in1;
	wire [0:0] eq_119_out;
	eq #(.WIDTH(32)) eq_119(.in0(eq_119_in0), .in1(eq_119_in1), .out(eq_119_out));

	reg [31:0] eq_120_in0;
	reg [31:0] eq_120_in1;
	wire [0:0] eq_120_out;
	eq #(.WIDTH(32)) eq_120(.in0(eq_120_in0), .in1(eq_120_in1), .out(eq_120_out));

	reg [0:0] notOp_121_in0;
	wire [0:0] notOp_121_out;
	notOp #(.WIDTH(1)) notOp_121(.in(notOp_121_in0), .out(notOp_121_out));

	reg [0:0] andOp_122_in0;
	reg [0:0] andOp_122_in1;
	wire [0:0] andOp_122_out;
	andOp #(.WIDTH(1)) andOp_122(.in0(andOp_122_in0), .in1(andOp_122_in1), .out(andOp_122_out));

	reg [31:0] eq_123_in0;
	reg [31:0] eq_123_in1;
	wire [0:0] eq_123_out;
	eq #(.WIDTH(32)) eq_123(.in0(eq_123_in0), .in1(eq_123_in1), .out(eq_123_out));

	reg [0:0] notOp_124_in0;
	wire [0:0] notOp_124_out;
	notOp #(.WIDTH(1)) notOp_124(.in(notOp_124_in0), .out(notOp_124_out));

	reg [0:0] andOp_125_in0;
	reg [0:0] andOp_125_in1;
	wire [0:0] andOp_125_out;
	andOp #(.WIDTH(1)) andOp_125(.in0(andOp_125_in0), .in1(andOp_125_in1), .out(andOp_125_out));

	reg [31:0] eq_126_in0;
	reg [31:0] eq_126_in1;
	wire [0:0] eq_126_out;
	eq #(.WIDTH(32)) eq_126(.in0(eq_126_in0), .in1(eq_126_in1), .out(eq_126_out));

	reg [0:0] notOp_127_in0;
	wire [0:0] notOp_127_out;
	notOp #(.WIDTH(1)) notOp_127(.in(notOp_127_in0), .out(notOp_127_out));

	reg [0:0] andOp_128_in0;
	reg [0:0] andOp_128_in1;
	wire [0:0] andOp_128_out;
	andOp #(.WIDTH(1)) andOp_128(.in0(andOp_128_in0), .in1(andOp_128_in1), .out(andOp_128_out));

	reg [31:0] eq_129_in0;
	reg [31:0] eq_129_in1;
	wire [0:0] eq_129_out;
	eq #(.WIDTH(32)) eq_129(.in0(eq_129_in0), .in1(eq_129_in1), .out(eq_129_out));

	reg [0:0] notOp_130_in0;
	wire [0:0] notOp_130_out;
	notOp #(.WIDTH(1)) notOp_130(.in(notOp_130_in0), .out(notOp_130_out));

	reg [0:0] andOp_131_in0;
	reg [0:0] andOp_131_in1;
	wire [0:0] andOp_131_out;
	andOp #(.WIDTH(1)) andOp_131(.in0(andOp_131_in0), .in1(andOp_131_in1), .out(andOp_131_out));

	reg [31:0] eq_132_in0;
	reg [31:0] eq_132_in1;
	wire [0:0] eq_132_out;
	eq #(.WIDTH(32)) eq_132(.in0(eq_132_in0), .in1(eq_132_in1), .out(eq_132_out));

	reg [0:0] notOp_133_in0;
	wire [0:0] notOp_133_out;
	notOp #(.WIDTH(1)) notOp_133(.in(notOp_133_in0), .out(notOp_133_out));

	reg [0:0] andOp_134_in0;
	reg [0:0] andOp_134_in1;
	wire [0:0] andOp_134_out;
	andOp #(.WIDTH(1)) andOp_134(.in0(andOp_134_in0), .in1(andOp_134_in1), .out(andOp_134_out));

	reg [31:0] eq_135_in0;
	reg [31:0] eq_135_in1;
	wire [0:0] eq_135_out;
	eq #(.WIDTH(32)) eq_135(.in0(eq_135_in0), .in1(eq_135_in1), .out(eq_135_out));

	reg [0:0] andOp_136_in0;
	reg [0:0] andOp_136_in1;
	wire [0:0] andOp_136_out;
	andOp #(.WIDTH(1)) andOp_136(.in0(andOp_136_in0), .in1(andOp_136_in1), .out(andOp_136_out));

	reg [0:0] andOp_137_in0;
	reg [0:0] andOp_137_in1;
	wire [0:0] andOp_137_out;
	andOp #(.WIDTH(1)) andOp_137(.in0(andOp_137_in0), .in1(andOp_137_in1), .out(andOp_137_out));

	reg [0:0] andOp_138_in0;
	reg [0:0] andOp_138_in1;
	wire [0:0] andOp_138_out;
	andOp #(.WIDTH(1)) andOp_138(.in0(andOp_138_in0), .in1(andOp_138_in1), .out(andOp_138_out));

	reg [0:0] andOp_139_in0;
	reg [0:0] andOp_139_in1;
	wire [0:0] andOp_139_out;
	andOp #(.WIDTH(1)) andOp_139(.in0(andOp_139_in0), .in1(andOp_139_in1), .out(andOp_139_out));

	reg [0:0] andOp_140_in0;
	reg [0:0] andOp_140_in1;
	wire [0:0] andOp_140_out;
	andOp #(.WIDTH(1)) andOp_140(.in0(andOp_140_in0), .in1(andOp_140_in1), .out(andOp_140_out));

	reg [0:0] andOp_141_in0;
	reg [0:0] andOp_141_in1;
	wire [0:0] andOp_141_out;
	andOp #(.WIDTH(1)) andOp_141(.in0(andOp_141_in0), .in1(andOp_141_in1), .out(andOp_141_out));

	reg [0:0] andOp_142_in0;
	reg [0:0] andOp_142_in1;
	wire [0:0] andOp_142_out;
	andOp #(.WIDTH(1)) andOp_142(.in0(andOp_142_in0), .in1(andOp_142_in1), .out(andOp_142_out));

	reg [0:0] andOp_143_in0;
	reg [0:0] andOp_143_in1;
	wire [0:0] andOp_143_out;
	andOp #(.WIDTH(1)) andOp_143(.in0(andOp_143_in0), .in1(andOp_143_in1), .out(andOp_143_out));

	reg [0:0] andOp_144_in0;
	reg [0:0] andOp_144_in1;
	wire [0:0] andOp_144_out;
	andOp #(.WIDTH(1)) andOp_144(.in0(andOp_144_in0), .in1(andOp_144_in1), .out(andOp_144_out));

	reg [0:0] andOp_145_in0;
	reg [0:0] andOp_145_in1;
	wire [0:0] andOp_145_out;
	andOp #(.WIDTH(1)) andOp_145(.in0(andOp_145_in0), .in1(andOp_145_in1), .out(andOp_145_out));

	reg [0:0] andOp_146_in0;
	reg [0:0] andOp_146_in1;
	wire [0:0] andOp_146_out;
	andOp #(.WIDTH(1)) andOp_146(.in0(andOp_146_in0), .in1(andOp_146_in1), .out(andOp_146_out));

	reg [31:0] concat_147_in0;
	reg [31:0] concat_147_in1;
	wire [63:0] concat_147_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_147(.in0(concat_147_in0), .in1(concat_147_in1), .out(concat_147_out));

	reg [31:0] concat_148_in0;
	reg [31:0] concat_148_in1;
	wire [63:0] concat_148_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_148(.in0(concat_148_in0), .in1(concat_148_in1), .out(concat_148_out));

	reg [0:0] andOp_149_in0;
	reg [0:0] andOp_149_in1;
	wire [0:0] andOp_149_out;
	andOp #(.WIDTH(1)) andOp_149(.in0(andOp_149_in0), .in1(andOp_149_in1), .out(andOp_149_out));

	reg [31:0] tmp_output_150_in_data;
	wire [31:0] tmp_output_150_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_150(.in_data(tmp_output_150_in_data), .out_data(tmp_output_150_out_data));

	reg [31:0] eq_151_in0;
	reg [31:0] eq_151_in1;
	wire [0:0] eq_151_out;
	eq #(.WIDTH(32)) eq_151(.in0(eq_151_in0), .in1(eq_151_in1), .out(eq_151_out));

	reg [0:0] andOp_152_in0;
	reg [0:0] andOp_152_in1;
	wire [0:0] andOp_152_out;
	andOp #(.WIDTH(1)) andOp_152(.in0(andOp_152_in0), .in1(andOp_152_in1), .out(andOp_152_out));

	reg [0:0] andOp_153_in0;
	reg [0:0] andOp_153_in1;
	wire [0:0] andOp_153_out;
	andOp #(.WIDTH(1)) andOp_153(.in0(andOp_153_in0), .in1(andOp_153_in1), .out(andOp_153_out));

	reg [0:0] andOp_154_in0;
	reg [0:0] andOp_154_in1;
	wire [0:0] andOp_154_out;
	andOp #(.WIDTH(1)) andOp_154(.in0(andOp_154_in0), .in1(andOp_154_in1), .out(andOp_154_out));

	reg [0:0] andOp_155_in0;
	reg [0:0] andOp_155_in1;
	wire [0:0] andOp_155_out;
	andOp #(.WIDTH(1)) andOp_155(.in0(andOp_155_in0), .in1(andOp_155_in1), .out(andOp_155_out));

	reg [0:0] andOp_156_in0;
	reg [0:0] andOp_156_in1;
	wire [0:0] andOp_156_out;
	andOp #(.WIDTH(1)) andOp_156(.in0(andOp_156_in0), .in1(andOp_156_in1), .out(andOp_156_out));

	reg [0:0] andOp_157_in0;
	reg [0:0] andOp_157_in1;
	wire [0:0] andOp_157_out;
	andOp #(.WIDTH(1)) andOp_157(.in0(andOp_157_in0), .in1(andOp_157_in1), .out(andOp_157_out));

	reg [0:0] andOp_158_in0;
	reg [0:0] andOp_158_in1;
	wire [0:0] andOp_158_out;
	andOp #(.WIDTH(1)) andOp_158(.in0(andOp_158_in0), .in1(andOp_158_in1), .out(andOp_158_out));

	reg [0:0] andOp_159_in0;
	reg [0:0] andOp_159_in1;
	wire [0:0] andOp_159_out;
	andOp #(.WIDTH(1)) andOp_159(.in0(andOp_159_in0), .in1(andOp_159_in1), .out(andOp_159_out));

	reg [0:0] andOp_160_in0;
	reg [0:0] andOp_160_in1;
	wire [0:0] andOp_160_out;
	andOp #(.WIDTH(1)) andOp_160(.in0(andOp_160_in0), .in1(andOp_160_in1), .out(andOp_160_out));

	reg [0:0] andOp_161_in0;
	reg [0:0] andOp_161_in1;
	wire [0:0] andOp_161_out;
	andOp #(.WIDTH(1)) andOp_161(.in0(andOp_161_in0), .in1(andOp_161_in1), .out(andOp_161_out));

	reg [0:0] andOp_162_in0;
	reg [0:0] andOp_162_in1;
	wire [0:0] andOp_162_out;
	andOp #(.WIDTH(1)) andOp_162(.in0(andOp_162_in0), .in1(andOp_162_in1), .out(andOp_162_out));

	reg [0:0] notOp_163_in0;
	wire [0:0] notOp_163_out;
	notOp #(.WIDTH(1)) notOp_163(.in(notOp_163_in0), .out(notOp_163_out));

	reg [0:0] andOp_164_in0;
	reg [0:0] andOp_164_in1;
	wire [0:0] andOp_164_out;
	andOp #(.WIDTH(1)) andOp_164(.in0(andOp_164_in0), .in1(andOp_164_in1), .out(andOp_164_out));

	reg [0:0] notOp_165_in0;
	wire [0:0] notOp_165_out;
	notOp #(.WIDTH(1)) notOp_165(.in(notOp_165_in0), .out(notOp_165_out));

	reg [0:0] andOp_166_in0;
	reg [0:0] andOp_166_in1;
	wire [0:0] andOp_166_out;
	andOp #(.WIDTH(1)) andOp_166(.in0(andOp_166_in0), .in1(andOp_166_in1), .out(andOp_166_out));

	reg [0:0] notOp_167_in0;
	wire [0:0] notOp_167_out;
	notOp #(.WIDTH(1)) notOp_167(.in(notOp_167_in0), .out(notOp_167_out));

	reg [0:0] andOp_168_in0;
	reg [0:0] andOp_168_in1;
	wire [0:0] andOp_168_out;
	andOp #(.WIDTH(1)) andOp_168(.in0(andOp_168_in0), .in1(andOp_168_in1), .out(andOp_168_out));

	reg [0:0] notOp_169_in0;
	wire [0:0] notOp_169_out;
	notOp #(.WIDTH(1)) notOp_169(.in(notOp_169_in0), .out(notOp_169_out));

	reg [0:0] andOp_170_in0;
	reg [0:0] andOp_170_in1;
	wire [0:0] andOp_170_out;
	andOp #(.WIDTH(1)) andOp_170(.in0(andOp_170_in0), .in1(andOp_170_in1), .out(andOp_170_out));

	reg [0:0] notOp_171_in0;
	wire [0:0] notOp_171_out;
	notOp #(.WIDTH(1)) notOp_171(.in(notOp_171_in0), .out(notOp_171_out));

	reg [0:0] andOp_172_in0;
	reg [0:0] andOp_172_in1;
	wire [0:0] andOp_172_out;
	andOp #(.WIDTH(1)) andOp_172(.in0(andOp_172_in0), .in1(andOp_172_in1), .out(andOp_172_out));

	reg [0:0] notOp_173_in0;
	wire [0:0] notOp_173_out;
	notOp #(.WIDTH(1)) notOp_173(.in(notOp_173_in0), .out(notOp_173_out));

	reg [0:0] andOp_174_in0;
	reg [0:0] andOp_174_in1;
	wire [0:0] andOp_174_out;
	andOp #(.WIDTH(1)) andOp_174(.in0(andOp_174_in0), .in1(andOp_174_in1), .out(andOp_174_out));

	reg [0:0] notOp_175_in0;
	wire [0:0] notOp_175_out;
	notOp #(.WIDTH(1)) notOp_175(.in(notOp_175_in0), .out(notOp_175_out));

	reg [0:0] andOp_176_in0;
	reg [0:0] andOp_176_in1;
	wire [0:0] andOp_176_out;
	andOp #(.WIDTH(1)) andOp_176(.in0(andOp_176_in0), .in1(andOp_176_in1), .out(andOp_176_out));

	reg [0:0] notOp_177_in0;
	wire [0:0] notOp_177_out;
	notOp #(.WIDTH(1)) notOp_177(.in(notOp_177_in0), .out(notOp_177_out));

	reg [0:0] andOp_178_in0;
	reg [0:0] andOp_178_in1;
	wire [0:0] andOp_178_out;
	andOp #(.WIDTH(1)) andOp_178(.in0(andOp_178_in0), .in1(andOp_178_in1), .out(andOp_178_out));

	reg [0:0] andOp_179_in0;
	reg [0:0] andOp_179_in1;
	wire [0:0] andOp_179_out;
	andOp #(.WIDTH(1)) andOp_179(.in0(andOp_179_in0), .in1(andOp_179_in1), .out(andOp_179_out));

	reg [0:0] andOp_180_in0;
	reg [0:0] andOp_180_in1;
	wire [0:0] andOp_180_out;
	andOp #(.WIDTH(1)) andOp_180(.in0(andOp_180_in0), .in1(andOp_180_in1), .out(andOp_180_out));

	reg [0:0] andOp_181_in0;
	reg [0:0] andOp_181_in1;
	wire [0:0] andOp_181_out;
	andOp #(.WIDTH(1)) andOp_181(.in0(andOp_181_in0), .in1(andOp_181_in1), .out(andOp_181_out));

	reg [0:0] andOp_182_in0;
	reg [0:0] andOp_182_in1;
	wire [0:0] andOp_182_out;
	andOp #(.WIDTH(1)) andOp_182(.in0(andOp_182_in0), .in1(andOp_182_in1), .out(andOp_182_out));

	reg [31:0] eq_183_in0;
	reg [31:0] eq_183_in1;
	wire [0:0] eq_183_out;
	eq #(.WIDTH(32)) eq_183(.in0(eq_183_in0), .in1(eq_183_in1), .out(eq_183_out));

	reg [0:0] andOp_184_in0;
	reg [0:0] andOp_184_in1;
	wire [0:0] andOp_184_out;
	andOp #(.WIDTH(1)) andOp_184(.in0(andOp_184_in0), .in1(andOp_184_in1), .out(andOp_184_out));

	reg [31:0] eq_185_in0;
	reg [31:0] eq_185_in1;
	wire [0:0] eq_185_out;
	eq #(.WIDTH(32)) eq_185(.in0(eq_185_in0), .in1(eq_185_in1), .out(eq_185_out));

	reg [0:0] andOp_186_in0;
	reg [0:0] andOp_186_in1;
	wire [0:0] andOp_186_out;
	andOp #(.WIDTH(1)) andOp_186(.in0(andOp_186_in0), .in1(andOp_186_in1), .out(andOp_186_out));

	reg [31:0] eq_187_in0;
	reg [31:0] eq_187_in1;
	wire [0:0] eq_187_out;
	eq #(.WIDTH(32)) eq_187(.in0(eq_187_in0), .in1(eq_187_in1), .out(eq_187_out));

	reg [0:0] andOp_188_in0;
	reg [0:0] andOp_188_in1;
	wire [0:0] andOp_188_out;
	andOp #(.WIDTH(1)) andOp_188(.in0(andOp_188_in0), .in1(andOp_188_in1), .out(andOp_188_out));

	reg [31:0] eq_189_in0;
	reg [31:0] eq_189_in1;
	wire [0:0] eq_189_out;
	eq #(.WIDTH(32)) eq_189(.in0(eq_189_in0), .in1(eq_189_in1), .out(eq_189_out));

	reg [0:0] andOp_190_in0;
	reg [0:0] andOp_190_in1;
	wire [0:0] andOp_190_out;
	andOp #(.WIDTH(1)) andOp_190(.in0(andOp_190_in0), .in1(andOp_190_in1), .out(andOp_190_out));

	reg [31:0] eq_191_in0;
	reg [31:0] eq_191_in1;
	wire [0:0] eq_191_out;
	eq #(.WIDTH(32)) eq_191(.in0(eq_191_in0), .in1(eq_191_in1), .out(eq_191_out));

	reg [0:0] andOp_192_in0;
	reg [0:0] andOp_192_in1;
	wire [0:0] andOp_192_out;
	andOp #(.WIDTH(1)) andOp_192(.in0(andOp_192_in0), .in1(andOp_192_in1), .out(andOp_192_out));

	reg [0:0] andOp_193_in0;
	reg [0:0] andOp_193_in1;
	wire [0:0] andOp_193_out;
	andOp #(.WIDTH(1)) andOp_193(.in0(andOp_193_in0), .in1(andOp_193_in1), .out(andOp_193_out));

	reg [31:0] eq_194_in0;
	reg [31:0] eq_194_in1;
	wire [0:0] eq_194_out;
	eq #(.WIDTH(32)) eq_194(.in0(eq_194_in0), .in1(eq_194_in1), .out(eq_194_out));

	reg [0:0] andOp_195_in0;
	reg [0:0] andOp_195_in1;
	wire [0:0] andOp_195_out;
	andOp #(.WIDTH(1)) andOp_195(.in0(andOp_195_in0), .in1(andOp_195_in1), .out(andOp_195_out));

	reg [0:0] notOp_196_in0;
	wire [0:0] notOp_196_out;
	notOp #(.WIDTH(1)) notOp_196(.in(notOp_196_in0), .out(notOp_196_out));

	reg [0:0] andOp_197_in0;
	reg [0:0] andOp_197_in1;
	wire [0:0] andOp_197_out;
	andOp #(.WIDTH(1)) andOp_197(.in0(andOp_197_in0), .in1(andOp_197_in1), .out(andOp_197_out));

	reg [0:0] notOp_198_in0;
	wire [0:0] notOp_198_out;
	notOp #(.WIDTH(1)) notOp_198(.in(notOp_198_in0), .out(notOp_198_out));

	reg [0:0] andOp_199_in0;
	reg [0:0] andOp_199_in1;
	wire [0:0] andOp_199_out;
	andOp #(.WIDTH(1)) andOp_199(.in0(andOp_199_in0), .in1(andOp_199_in1), .out(andOp_199_out));

	reg [0:0] notOp_200_in0;
	wire [0:0] notOp_200_out;
	notOp #(.WIDTH(1)) notOp_200(.in(notOp_200_in0), .out(notOp_200_out));

	reg [0:0] andOp_201_in0;
	reg [0:0] andOp_201_in1;
	wire [0:0] andOp_201_out;
	andOp #(.WIDTH(1)) andOp_201(.in0(andOp_201_in0), .in1(andOp_201_in1), .out(andOp_201_out));

	reg [0:0] andOp_202_in0;
	reg [0:0] andOp_202_in1;
	wire [0:0] andOp_202_out;
	andOp #(.WIDTH(1)) andOp_202(.in0(andOp_202_in0), .in1(andOp_202_in1), .out(andOp_202_out));

	reg [31:0] eq_203_in0;
	reg [31:0] eq_203_in1;
	wire [0:0] eq_203_out;
	eq #(.WIDTH(32)) eq_203(.in0(eq_203_in0), .in1(eq_203_in1), .out(eq_203_out));

	reg [0:0] andOp_204_in0;
	reg [0:0] andOp_204_in1;
	wire [0:0] andOp_204_out;
	andOp #(.WIDTH(1)) andOp_204(.in0(andOp_204_in0), .in1(andOp_204_in1), .out(andOp_204_out));

	reg [0:0] notOp_205_in0;
	wire [0:0] notOp_205_out;
	notOp #(.WIDTH(1)) notOp_205(.in(notOp_205_in0), .out(notOp_205_out));

	reg [0:0] andOp_206_in0;
	reg [0:0] andOp_206_in1;
	wire [0:0] andOp_206_out;
	andOp #(.WIDTH(1)) andOp_206(.in0(andOp_206_in0), .in1(andOp_206_in1), .out(andOp_206_out));

	reg [0:0] notOp_207_in0;
	wire [0:0] notOp_207_out;
	notOp #(.WIDTH(1)) notOp_207(.in(notOp_207_in0), .out(notOp_207_out));

	reg [0:0] andOp_208_in0;
	reg [0:0] andOp_208_in1;
	wire [0:0] andOp_208_out;
	andOp #(.WIDTH(1)) andOp_208(.in0(andOp_208_in0), .in1(andOp_208_in1), .out(andOp_208_out));

	reg [0:0] notOp_209_in0;
	wire [0:0] notOp_209_out;
	notOp #(.WIDTH(1)) notOp_209(.in(notOp_209_in0), .out(notOp_209_out));

	reg [0:0] andOp_210_in0;
	reg [0:0] andOp_210_in1;
	wire [0:0] andOp_210_out;
	andOp #(.WIDTH(1)) andOp_210(.in0(andOp_210_in0), .in1(andOp_210_in1), .out(andOp_210_out));

	reg [0:0] andOp_211_in0;
	reg [0:0] andOp_211_in1;
	wire [0:0] andOp_211_out;
	andOp #(.WIDTH(1)) andOp_211(.in0(andOp_211_in0), .in1(andOp_211_in1), .out(andOp_211_out));

	reg [31:0] eq_212_in0;
	reg [31:0] eq_212_in1;
	wire [0:0] eq_212_out;
	eq #(.WIDTH(32)) eq_212(.in0(eq_212_in0), .in1(eq_212_in1), .out(eq_212_out));

	reg [0:0] andOp_213_in0;
	reg [0:0] andOp_213_in1;
	wire [0:0] andOp_213_out;
	andOp #(.WIDTH(1)) andOp_213(.in0(andOp_213_in0), .in1(andOp_213_in1), .out(andOp_213_out));

	reg [0:0] notOp_214_in0;
	wire [0:0] notOp_214_out;
	notOp #(.WIDTH(1)) notOp_214(.in(notOp_214_in0), .out(notOp_214_out));

	reg [0:0] andOp_215_in0;
	reg [0:0] andOp_215_in1;
	wire [0:0] andOp_215_out;
	andOp #(.WIDTH(1)) andOp_215(.in0(andOp_215_in0), .in1(andOp_215_in1), .out(andOp_215_out));

	reg [0:0] notOp_216_in0;
	wire [0:0] notOp_216_out;
	notOp #(.WIDTH(1)) notOp_216(.in(notOp_216_in0), .out(notOp_216_out));

	reg [0:0] andOp_217_in0;
	reg [0:0] andOp_217_in1;
	wire [0:0] andOp_217_out;
	andOp #(.WIDTH(1)) andOp_217(.in0(andOp_217_in0), .in1(andOp_217_in1), .out(andOp_217_out));

	reg [0:0] notOp_218_in0;
	wire [0:0] notOp_218_out;
	notOp #(.WIDTH(1)) notOp_218(.in(notOp_218_in0), .out(notOp_218_out));

	reg [0:0] andOp_219_in0;
	reg [0:0] andOp_219_in1;
	wire [0:0] andOp_219_out;
	andOp #(.WIDTH(1)) andOp_219(.in0(andOp_219_in0), .in1(andOp_219_in1), .out(andOp_219_out));

	reg [31:0] eq_220_in0;
	reg [31:0] eq_220_in1;
	wire [0:0] eq_220_out;
	eq #(.WIDTH(32)) eq_220(.in0(eq_220_in0), .in1(eq_220_in1), .out(eq_220_out));

	reg [0:0] andOp_221_in0;
	reg [0:0] andOp_221_in1;
	wire [0:0] andOp_221_out;
	andOp #(.WIDTH(1)) andOp_221(.in0(andOp_221_in0), .in1(andOp_221_in1), .out(andOp_221_out));

	reg [31:0] eq_222_in0;
	reg [31:0] eq_222_in1;
	wire [0:0] eq_222_out;
	eq #(.WIDTH(32)) eq_222(.in0(eq_222_in0), .in1(eq_222_in1), .out(eq_222_out));

	reg [0:0] andOp_223_in0;
	reg [0:0] andOp_223_in1;
	wire [0:0] andOp_223_out;
	andOp #(.WIDTH(1)) andOp_223(.in0(andOp_223_in0), .in1(andOp_223_in1), .out(andOp_223_out));

	reg [31:0] eq_224_in0;
	reg [31:0] eq_224_in1;
	wire [0:0] eq_224_out;
	eq #(.WIDTH(32)) eq_224(.in0(eq_224_in0), .in1(eq_224_in1), .out(eq_224_out));

	reg [0:0] andOp_225_in0;
	reg [0:0] andOp_225_in1;
	wire [0:0] andOp_225_out;
	andOp #(.WIDTH(1)) andOp_225(.in0(andOp_225_in0), .in1(andOp_225_in1), .out(andOp_225_out));

	reg [31:0] eq_226_in0;
	reg [31:0] eq_226_in1;
	wire [0:0] eq_226_out;
	eq #(.WIDTH(32)) eq_226(.in0(eq_226_in0), .in1(eq_226_in1), .out(eq_226_out));

	reg [0:0] andOp_227_in0;
	reg [0:0] andOp_227_in1;
	wire [0:0] andOp_227_out;
	andOp #(.WIDTH(1)) andOp_227(.in0(andOp_227_in0), .in1(andOp_227_in1), .out(andOp_227_out));

	reg [31:0] eq_228_in0;
	reg [31:0] eq_228_in1;
	wire [0:0] eq_228_out;
	eq #(.WIDTH(32)) eq_228(.in0(eq_228_in0), .in1(eq_228_in1), .out(eq_228_out));

	reg [0:0] andOp_229_in0;
	reg [0:0] andOp_229_in1;
	wire [0:0] andOp_229_out;
	andOp #(.WIDTH(1)) andOp_229(.in0(andOp_229_in0), .in1(andOp_229_in1), .out(andOp_229_out));

	reg [0:0] andOp_230_in0;
	reg [0:0] andOp_230_in1;
	wire [0:0] andOp_230_out;
	andOp #(.WIDTH(1)) andOp_230(.in0(andOp_230_in0), .in1(andOp_230_in1), .out(andOp_230_out));

	reg [31:0] eq_231_in0;
	reg [31:0] eq_231_in1;
	wire [0:0] eq_231_out;
	eq #(.WIDTH(32)) eq_231(.in0(eq_231_in0), .in1(eq_231_in1), .out(eq_231_out));

	reg [0:0] andOp_232_in0;
	reg [0:0] andOp_232_in1;
	wire [0:0] andOp_232_out;
	andOp #(.WIDTH(1)) andOp_232(.in0(andOp_232_in0), .in1(andOp_232_in1), .out(andOp_232_out));

	reg [0:0] notOp_233_in0;
	wire [0:0] notOp_233_out;
	notOp #(.WIDTH(1)) notOp_233(.in(notOp_233_in0), .out(notOp_233_out));

	reg [0:0] andOp_234_in0;
	reg [0:0] andOp_234_in1;
	wire [0:0] andOp_234_out;
	andOp #(.WIDTH(1)) andOp_234(.in0(andOp_234_in0), .in1(andOp_234_in1), .out(andOp_234_out));

	reg [0:0] notOp_235_in0;
	wire [0:0] notOp_235_out;
	notOp #(.WIDTH(1)) notOp_235(.in(notOp_235_in0), .out(notOp_235_out));

	reg [0:0] andOp_236_in0;
	reg [0:0] andOp_236_in1;
	wire [0:0] andOp_236_out;
	andOp #(.WIDTH(1)) andOp_236(.in0(andOp_236_in0), .in1(andOp_236_in1), .out(andOp_236_out));

	reg [0:0] notOp_237_in0;
	wire [0:0] notOp_237_out;
	notOp #(.WIDTH(1)) notOp_237(.in(notOp_237_in0), .out(notOp_237_out));

	reg [0:0] andOp_238_in0;
	reg [0:0] andOp_238_in1;
	wire [0:0] andOp_238_out;
	andOp #(.WIDTH(1)) andOp_238(.in0(andOp_238_in0), .in1(andOp_238_in1), .out(andOp_238_out));

	reg [0:0] andOp_239_in0;
	reg [0:0] andOp_239_in1;
	wire [0:0] andOp_239_out;
	andOp #(.WIDTH(1)) andOp_239(.in0(andOp_239_in0), .in1(andOp_239_in1), .out(andOp_239_out));

	reg [31:0] eq_240_in0;
	reg [31:0] eq_240_in1;
	wire [0:0] eq_240_out;
	eq #(.WIDTH(32)) eq_240(.in0(eq_240_in0), .in1(eq_240_in1), .out(eq_240_out));

	reg [0:0] andOp_241_in0;
	reg [0:0] andOp_241_in1;
	wire [0:0] andOp_241_out;
	andOp #(.WIDTH(1)) andOp_241(.in0(andOp_241_in0), .in1(andOp_241_in1), .out(andOp_241_out));

	reg [0:0] notOp_242_in0;
	wire [0:0] notOp_242_out;
	notOp #(.WIDTH(1)) notOp_242(.in(notOp_242_in0), .out(notOp_242_out));

	reg [0:0] andOp_243_in0;
	reg [0:0] andOp_243_in1;
	wire [0:0] andOp_243_out;
	andOp #(.WIDTH(1)) andOp_243(.in0(andOp_243_in0), .in1(andOp_243_in1), .out(andOp_243_out));

	reg [0:0] notOp_244_in0;
	wire [0:0] notOp_244_out;
	notOp #(.WIDTH(1)) notOp_244(.in(notOp_244_in0), .out(notOp_244_out));

	reg [0:0] andOp_245_in0;
	reg [0:0] andOp_245_in1;
	wire [0:0] andOp_245_out;
	andOp #(.WIDTH(1)) andOp_245(.in0(andOp_245_in0), .in1(andOp_245_in1), .out(andOp_245_out));

	reg [0:0] notOp_246_in0;
	wire [0:0] notOp_246_out;
	notOp #(.WIDTH(1)) notOp_246(.in(notOp_246_in0), .out(notOp_246_out));

	reg [0:0] andOp_247_in0;
	reg [0:0] andOp_247_in1;
	wire [0:0] andOp_247_out;
	andOp #(.WIDTH(1)) andOp_247(.in0(andOp_247_in0), .in1(andOp_247_in1), .out(andOp_247_out));

	reg [0:0] andOp_248_in0;
	reg [0:0] andOp_248_in1;
	wire [0:0] andOp_248_out;
	andOp #(.WIDTH(1)) andOp_248(.in0(andOp_248_in0), .in1(andOp_248_in1), .out(andOp_248_out));

	reg [31:0] eq_249_in0;
	reg [31:0] eq_249_in1;
	wire [0:0] eq_249_out;
	eq #(.WIDTH(32)) eq_249(.in0(eq_249_in0), .in1(eq_249_in1), .out(eq_249_out));

	reg [0:0] andOp_250_in0;
	reg [0:0] andOp_250_in1;
	wire [0:0] andOp_250_out;
	andOp #(.WIDTH(1)) andOp_250(.in0(andOp_250_in0), .in1(andOp_250_in1), .out(andOp_250_out));

	reg [0:0] notOp_251_in0;
	wire [0:0] notOp_251_out;
	notOp #(.WIDTH(1)) notOp_251(.in(notOp_251_in0), .out(notOp_251_out));

	reg [0:0] andOp_252_in0;
	reg [0:0] andOp_252_in1;
	wire [0:0] andOp_252_out;
	andOp #(.WIDTH(1)) andOp_252(.in0(andOp_252_in0), .in1(andOp_252_in1), .out(andOp_252_out));

	reg [0:0] notOp_253_in0;
	wire [0:0] notOp_253_out;
	notOp #(.WIDTH(1)) notOp_253(.in(notOp_253_in0), .out(notOp_253_out));

	reg [0:0] andOp_254_in0;
	reg [0:0] andOp_254_in1;
	wire [0:0] andOp_254_out;
	andOp #(.WIDTH(1)) andOp_254(.in0(andOp_254_in0), .in1(andOp_254_in1), .out(andOp_254_out));

	reg [0:0] notOp_255_in0;
	wire [0:0] notOp_255_out;
	notOp #(.WIDTH(1)) notOp_255(.in(notOp_255_in0), .out(notOp_255_out));

	reg [0:0] andOp_256_in0;
	reg [0:0] andOp_256_in1;
	wire [0:0] andOp_256_out;
	andOp #(.WIDTH(1)) andOp_256(.in0(andOp_256_in0), .in1(andOp_256_in1), .out(andOp_256_out));

	reg [31:0] eq_257_in0;
	reg [31:0] eq_257_in1;
	wire [0:0] eq_257_out;
	eq #(.WIDTH(32)) eq_257(.in0(eq_257_in0), .in1(eq_257_in1), .out(eq_257_out));

	reg [0:0] andOp_258_in0;
	reg [0:0] andOp_258_in1;
	wire [0:0] andOp_258_out;
	andOp #(.WIDTH(1)) andOp_258(.in0(andOp_258_in0), .in1(andOp_258_in1), .out(andOp_258_out));

	reg [31:0] eq_259_in0;
	reg [31:0] eq_259_in1;
	wire [0:0] eq_259_out;
	eq #(.WIDTH(32)) eq_259(.in0(eq_259_in0), .in1(eq_259_in1), .out(eq_259_out));

	reg [0:0] andOp_260_in0;
	reg [0:0] andOp_260_in1;
	wire [0:0] andOp_260_out;
	andOp #(.WIDTH(1)) andOp_260(.in0(andOp_260_in0), .in1(andOp_260_in1), .out(andOp_260_out));

	reg [31:0] eq_261_in0;
	reg [31:0] eq_261_in1;
	wire [0:0] eq_261_out;
	eq #(.WIDTH(32)) eq_261(.in0(eq_261_in0), .in1(eq_261_in1), .out(eq_261_out));

	reg [0:0] andOp_262_in0;
	reg [0:0] andOp_262_in1;
	wire [0:0] andOp_262_out;
	andOp #(.WIDTH(1)) andOp_262(.in0(andOp_262_in0), .in1(andOp_262_in1), .out(andOp_262_out));

	reg [31:0] eq_263_in0;
	reg [31:0] eq_263_in1;
	wire [0:0] eq_263_out;
	eq #(.WIDTH(32)) eq_263(.in0(eq_263_in0), .in1(eq_263_in1), .out(eq_263_out));

	reg [0:0] andOp_264_in0;
	reg [0:0] andOp_264_in1;
	wire [0:0] andOp_264_out;
	andOp #(.WIDTH(1)) andOp_264(.in0(andOp_264_in0), .in1(andOp_264_in1), .out(andOp_264_out));

	reg [31:0] eq_265_in0;
	reg [31:0] eq_265_in1;
	wire [0:0] eq_265_out;
	eq #(.WIDTH(32)) eq_265(.in0(eq_265_in0), .in1(eq_265_in1), .out(eq_265_out));

	reg [0:0] andOp_266_in0;
	reg [0:0] andOp_266_in1;
	wire [0:0] andOp_266_out;
	andOp #(.WIDTH(1)) andOp_266(.in0(andOp_266_in0), .in1(andOp_266_in1), .out(andOp_266_out));

	reg [0:0] andOp_267_in0;
	reg [0:0] andOp_267_in1;
	wire [0:0] andOp_267_out;
	andOp #(.WIDTH(1)) andOp_267(.in0(andOp_267_in0), .in1(andOp_267_in1), .out(andOp_267_out));

	reg [31:0] eq_268_in0;
	reg [31:0] eq_268_in1;
	wire [0:0] eq_268_out;
	eq #(.WIDTH(32)) eq_268(.in0(eq_268_in0), .in1(eq_268_in1), .out(eq_268_out));

	reg [0:0] andOp_269_in0;
	reg [0:0] andOp_269_in1;
	wire [0:0] andOp_269_out;
	andOp #(.WIDTH(1)) andOp_269(.in0(andOp_269_in0), .in1(andOp_269_in1), .out(andOp_269_out));

	reg [0:0] notOp_270_in0;
	wire [0:0] notOp_270_out;
	notOp #(.WIDTH(1)) notOp_270(.in(notOp_270_in0), .out(notOp_270_out));

	reg [0:0] andOp_271_in0;
	reg [0:0] andOp_271_in1;
	wire [0:0] andOp_271_out;
	andOp #(.WIDTH(1)) andOp_271(.in0(andOp_271_in0), .in1(andOp_271_in1), .out(andOp_271_out));

	reg [0:0] notOp_272_in0;
	wire [0:0] notOp_272_out;
	notOp #(.WIDTH(1)) notOp_272(.in(notOp_272_in0), .out(notOp_272_out));

	reg [0:0] andOp_273_in0;
	reg [0:0] andOp_273_in1;
	wire [0:0] andOp_273_out;
	andOp #(.WIDTH(1)) andOp_273(.in0(andOp_273_in0), .in1(andOp_273_in1), .out(andOp_273_out));

	reg [0:0] notOp_274_in0;
	wire [0:0] notOp_274_out;
	notOp #(.WIDTH(1)) notOp_274(.in(notOp_274_in0), .out(notOp_274_out));

	reg [0:0] andOp_275_in0;
	reg [0:0] andOp_275_in1;
	wire [0:0] andOp_275_out;
	andOp #(.WIDTH(1)) andOp_275(.in0(andOp_275_in0), .in1(andOp_275_in1), .out(andOp_275_out));

	reg [0:0] andOp_276_in0;
	reg [0:0] andOp_276_in1;
	wire [0:0] andOp_276_out;
	andOp #(.WIDTH(1)) andOp_276(.in0(andOp_276_in0), .in1(andOp_276_in1), .out(andOp_276_out));

	reg [31:0] eq_277_in0;
	reg [31:0] eq_277_in1;
	wire [0:0] eq_277_out;
	eq #(.WIDTH(32)) eq_277(.in0(eq_277_in0), .in1(eq_277_in1), .out(eq_277_out));

	reg [0:0] andOp_278_in0;
	reg [0:0] andOp_278_in1;
	wire [0:0] andOp_278_out;
	andOp #(.WIDTH(1)) andOp_278(.in0(andOp_278_in0), .in1(andOp_278_in1), .out(andOp_278_out));

	reg [0:0] notOp_279_in0;
	wire [0:0] notOp_279_out;
	notOp #(.WIDTH(1)) notOp_279(.in(notOp_279_in0), .out(notOp_279_out));

	reg [0:0] andOp_280_in0;
	reg [0:0] andOp_280_in1;
	wire [0:0] andOp_280_out;
	andOp #(.WIDTH(1)) andOp_280(.in0(andOp_280_in0), .in1(andOp_280_in1), .out(andOp_280_out));

	reg [0:0] notOp_281_in0;
	wire [0:0] notOp_281_out;
	notOp #(.WIDTH(1)) notOp_281(.in(notOp_281_in0), .out(notOp_281_out));

	reg [0:0] andOp_282_in0;
	reg [0:0] andOp_282_in1;
	wire [0:0] andOp_282_out;
	andOp #(.WIDTH(1)) andOp_282(.in0(andOp_282_in0), .in1(andOp_282_in1), .out(andOp_282_out));

	reg [0:0] notOp_283_in0;
	wire [0:0] notOp_283_out;
	notOp #(.WIDTH(1)) notOp_283(.in(notOp_283_in0), .out(notOp_283_out));

	reg [0:0] andOp_284_in0;
	reg [0:0] andOp_284_in1;
	wire [0:0] andOp_284_out;
	andOp #(.WIDTH(1)) andOp_284(.in0(andOp_284_in0), .in1(andOp_284_in1), .out(andOp_284_out));

	reg [0:0] andOp_285_in0;
	reg [0:0] andOp_285_in1;
	wire [0:0] andOp_285_out;
	andOp #(.WIDTH(1)) andOp_285(.in0(andOp_285_in0), .in1(andOp_285_in1), .out(andOp_285_out));

	reg [31:0] eq_286_in0;
	reg [31:0] eq_286_in1;
	wire [0:0] eq_286_out;
	eq #(.WIDTH(32)) eq_286(.in0(eq_286_in0), .in1(eq_286_in1), .out(eq_286_out));

	reg [0:0] andOp_287_in0;
	reg [0:0] andOp_287_in1;
	wire [0:0] andOp_287_out;
	andOp #(.WIDTH(1)) andOp_287(.in0(andOp_287_in0), .in1(andOp_287_in1), .out(andOp_287_out));

	reg [0:0] notOp_288_in0;
	wire [0:0] notOp_288_out;
	notOp #(.WIDTH(1)) notOp_288(.in(notOp_288_in0), .out(notOp_288_out));

	reg [0:0] andOp_289_in0;
	reg [0:0] andOp_289_in1;
	wire [0:0] andOp_289_out;
	andOp #(.WIDTH(1)) andOp_289(.in0(andOp_289_in0), .in1(andOp_289_in1), .out(andOp_289_out));

	reg [0:0] notOp_290_in0;
	wire [0:0] notOp_290_out;
	notOp #(.WIDTH(1)) notOp_290(.in(notOp_290_in0), .out(notOp_290_out));

	reg [0:0] andOp_291_in0;
	reg [0:0] andOp_291_in1;
	wire [0:0] andOp_291_out;
	andOp #(.WIDTH(1)) andOp_291(.in0(andOp_291_in0), .in1(andOp_291_in1), .out(andOp_291_out));

	reg [0:0] notOp_292_in0;
	wire [0:0] notOp_292_out;
	notOp #(.WIDTH(1)) notOp_292(.in(notOp_292_in0), .out(notOp_292_out));

	reg [0:0] andOp_293_in0;
	reg [0:0] andOp_293_in1;
	wire [0:0] andOp_293_out;
	andOp #(.WIDTH(1)) andOp_293(.in0(andOp_293_in0), .in1(andOp_293_in1), .out(andOp_293_out));

	reg [31:0] eq_294_in0;
	reg [31:0] eq_294_in1;
	wire [0:0] eq_294_out;
	eq #(.WIDTH(32)) eq_294(.in0(eq_294_in0), .in1(eq_294_in1), .out(eq_294_out));

	reg [0:0] andOp_295_in0;
	reg [0:0] andOp_295_in1;
	wire [0:0] andOp_295_out;
	andOp #(.WIDTH(1)) andOp_295(.in0(andOp_295_in0), .in1(andOp_295_in1), .out(andOp_295_out));

	reg [31:0] eq_296_in0;
	reg [31:0] eq_296_in1;
	wire [0:0] eq_296_out;
	eq #(.WIDTH(32)) eq_296(.in0(eq_296_in0), .in1(eq_296_in1), .out(eq_296_out));

	reg [0:0] andOp_297_in0;
	reg [0:0] andOp_297_in1;
	wire [0:0] andOp_297_out;
	andOp #(.WIDTH(1)) andOp_297(.in0(andOp_297_in0), .in1(andOp_297_in1), .out(andOp_297_out));

	reg [31:0] eq_298_in0;
	reg [31:0] eq_298_in1;
	wire [0:0] eq_298_out;
	eq #(.WIDTH(32)) eq_298(.in0(eq_298_in0), .in1(eq_298_in1), .out(eq_298_out));

	reg [0:0] andOp_299_in0;
	reg [0:0] andOp_299_in1;
	wire [0:0] andOp_299_out;
	andOp #(.WIDTH(1)) andOp_299(.in0(andOp_299_in0), .in1(andOp_299_in1), .out(andOp_299_out));

	reg [31:0] eq_300_in0;
	reg [31:0] eq_300_in1;
	wire [0:0] eq_300_out;
	eq #(.WIDTH(32)) eq_300(.in0(eq_300_in0), .in1(eq_300_in1), .out(eq_300_out));

	reg [0:0] andOp_301_in0;
	reg [0:0] andOp_301_in1;
	wire [0:0] andOp_301_out;
	andOp #(.WIDTH(1)) andOp_301(.in0(andOp_301_in0), .in1(andOp_301_in1), .out(andOp_301_out));

	reg [31:0] eq_302_in0;
	reg [31:0] eq_302_in1;
	wire [0:0] eq_302_out;
	eq #(.WIDTH(32)) eq_302(.in0(eq_302_in0), .in1(eq_302_in1), .out(eq_302_out));

	reg [0:0] andOp_303_in0;
	reg [0:0] andOp_303_in1;
	wire [0:0] andOp_303_out;
	andOp #(.WIDTH(1)) andOp_303(.in0(andOp_303_in0), .in1(andOp_303_in1), .out(andOp_303_out));

	reg [0:0] andOp_304_in0;
	reg [0:0] andOp_304_in1;
	wire [0:0] andOp_304_out;
	andOp #(.WIDTH(1)) andOp_304(.in0(andOp_304_in0), .in1(andOp_304_in1), .out(andOp_304_out));

	reg [31:0] eq_305_in0;
	reg [31:0] eq_305_in1;
	wire [0:0] eq_305_out;
	eq #(.WIDTH(32)) eq_305(.in0(eq_305_in0), .in1(eq_305_in1), .out(eq_305_out));

	reg [0:0] andOp_306_in0;
	reg [0:0] andOp_306_in1;
	wire [0:0] andOp_306_out;
	andOp #(.WIDTH(1)) andOp_306(.in0(andOp_306_in0), .in1(andOp_306_in1), .out(andOp_306_out));

	reg [0:0] notOp_307_in0;
	wire [0:0] notOp_307_out;
	notOp #(.WIDTH(1)) notOp_307(.in(notOp_307_in0), .out(notOp_307_out));

	reg [0:0] andOp_308_in0;
	reg [0:0] andOp_308_in1;
	wire [0:0] andOp_308_out;
	andOp #(.WIDTH(1)) andOp_308(.in0(andOp_308_in0), .in1(andOp_308_in1), .out(andOp_308_out));

	reg [0:0] notOp_309_in0;
	wire [0:0] notOp_309_out;
	notOp #(.WIDTH(1)) notOp_309(.in(notOp_309_in0), .out(notOp_309_out));

	reg [0:0] andOp_310_in0;
	reg [0:0] andOp_310_in1;
	wire [0:0] andOp_310_out;
	andOp #(.WIDTH(1)) andOp_310(.in0(andOp_310_in0), .in1(andOp_310_in1), .out(andOp_310_out));

	reg [0:0] notOp_311_in0;
	wire [0:0] notOp_311_out;
	notOp #(.WIDTH(1)) notOp_311(.in(notOp_311_in0), .out(notOp_311_out));

	reg [0:0] andOp_312_in0;
	reg [0:0] andOp_312_in1;
	wire [0:0] andOp_312_out;
	andOp #(.WIDTH(1)) andOp_312(.in0(andOp_312_in0), .in1(andOp_312_in1), .out(andOp_312_out));

	reg [0:0] andOp_313_in0;
	reg [0:0] andOp_313_in1;
	wire [0:0] andOp_313_out;
	andOp #(.WIDTH(1)) andOp_313(.in0(andOp_313_in0), .in1(andOp_313_in1), .out(andOp_313_out));

	reg [31:0] eq_314_in0;
	reg [31:0] eq_314_in1;
	wire [0:0] eq_314_out;
	eq #(.WIDTH(32)) eq_314(.in0(eq_314_in0), .in1(eq_314_in1), .out(eq_314_out));

	reg [0:0] andOp_315_in0;
	reg [0:0] andOp_315_in1;
	wire [0:0] andOp_315_out;
	andOp #(.WIDTH(1)) andOp_315(.in0(andOp_315_in0), .in1(andOp_315_in1), .out(andOp_315_out));

	reg [0:0] notOp_316_in0;
	wire [0:0] notOp_316_out;
	notOp #(.WIDTH(1)) notOp_316(.in(notOp_316_in0), .out(notOp_316_out));

	reg [0:0] andOp_317_in0;
	reg [0:0] andOp_317_in1;
	wire [0:0] andOp_317_out;
	andOp #(.WIDTH(1)) andOp_317(.in0(andOp_317_in0), .in1(andOp_317_in1), .out(andOp_317_out));

	reg [0:0] notOp_318_in0;
	wire [0:0] notOp_318_out;
	notOp #(.WIDTH(1)) notOp_318(.in(notOp_318_in0), .out(notOp_318_out));

	reg [0:0] andOp_319_in0;
	reg [0:0] andOp_319_in1;
	wire [0:0] andOp_319_out;
	andOp #(.WIDTH(1)) andOp_319(.in0(andOp_319_in0), .in1(andOp_319_in1), .out(andOp_319_out));

	reg [0:0] notOp_320_in0;
	wire [0:0] notOp_320_out;
	notOp #(.WIDTH(1)) notOp_320(.in(notOp_320_in0), .out(notOp_320_out));

	reg [0:0] andOp_321_in0;
	reg [0:0] andOp_321_in1;
	wire [0:0] andOp_321_out;
	andOp #(.WIDTH(1)) andOp_321(.in0(andOp_321_in0), .in1(andOp_321_in1), .out(andOp_321_out));

	reg [0:0] andOp_322_in0;
	reg [0:0] andOp_322_in1;
	wire [0:0] andOp_322_out;
	andOp #(.WIDTH(1)) andOp_322(.in0(andOp_322_in0), .in1(andOp_322_in1), .out(andOp_322_out));

	reg [31:0] eq_323_in0;
	reg [31:0] eq_323_in1;
	wire [0:0] eq_323_out;
	eq #(.WIDTH(32)) eq_323(.in0(eq_323_in0), .in1(eq_323_in1), .out(eq_323_out));

	reg [0:0] andOp_324_in0;
	reg [0:0] andOp_324_in1;
	wire [0:0] andOp_324_out;
	andOp #(.WIDTH(1)) andOp_324(.in0(andOp_324_in0), .in1(andOp_324_in1), .out(andOp_324_out));

	reg [0:0] notOp_325_in0;
	wire [0:0] notOp_325_out;
	notOp #(.WIDTH(1)) notOp_325(.in(notOp_325_in0), .out(notOp_325_out));

	reg [0:0] andOp_326_in0;
	reg [0:0] andOp_326_in1;
	wire [0:0] andOp_326_out;
	andOp #(.WIDTH(1)) andOp_326(.in0(andOp_326_in0), .in1(andOp_326_in1), .out(andOp_326_out));

	reg [0:0] notOp_327_in0;
	wire [0:0] notOp_327_out;
	notOp #(.WIDTH(1)) notOp_327(.in(notOp_327_in0), .out(notOp_327_out));

	reg [0:0] andOp_328_in0;
	reg [0:0] andOp_328_in1;
	wire [0:0] andOp_328_out;
	andOp #(.WIDTH(1)) andOp_328(.in0(andOp_328_in0), .in1(andOp_328_in1), .out(andOp_328_out));

	reg [0:0] notOp_329_in0;
	wire [0:0] notOp_329_out;
	notOp #(.WIDTH(1)) notOp_329(.in(notOp_329_in0), .out(notOp_329_out));

	reg [0:0] andOp_330_in0;
	reg [0:0] andOp_330_in1;
	wire [0:0] andOp_330_out;
	andOp #(.WIDTH(1)) andOp_330(.in0(andOp_330_in0), .in1(andOp_330_in1), .out(andOp_330_out));

	reg [31:0] eq_331_in0;
	reg [31:0] eq_331_in1;
	wire [0:0] eq_331_out;
	eq #(.WIDTH(32)) eq_331(.in0(eq_331_in0), .in1(eq_331_in1), .out(eq_331_out));

	reg [0:0] andOp_332_in0;
	reg [0:0] andOp_332_in1;
	wire [0:0] andOp_332_out;
	andOp #(.WIDTH(1)) andOp_332(.in0(andOp_332_in0), .in1(andOp_332_in1), .out(andOp_332_out));

	reg [31:0] eq_333_in0;
	reg [31:0] eq_333_in1;
	wire [0:0] eq_333_out;
	eq #(.WIDTH(32)) eq_333(.in0(eq_333_in0), .in1(eq_333_in1), .out(eq_333_out));

	reg [0:0] andOp_334_in0;
	reg [0:0] andOp_334_in1;
	wire [0:0] andOp_334_out;
	andOp #(.WIDTH(1)) andOp_334(.in0(andOp_334_in0), .in1(andOp_334_in1), .out(andOp_334_out));

	reg [31:0] eq_335_in0;
	reg [31:0] eq_335_in1;
	wire [0:0] eq_335_out;
	eq #(.WIDTH(32)) eq_335(.in0(eq_335_in0), .in1(eq_335_in1), .out(eq_335_out));

	reg [0:0] andOp_336_in0;
	reg [0:0] andOp_336_in1;
	wire [0:0] andOp_336_out;
	andOp #(.WIDTH(1)) andOp_336(.in0(andOp_336_in0), .in1(andOp_336_in1), .out(andOp_336_out));

	reg [31:0] eq_337_in0;
	reg [31:0] eq_337_in1;
	wire [0:0] eq_337_out;
	eq #(.WIDTH(32)) eq_337(.in0(eq_337_in0), .in1(eq_337_in1), .out(eq_337_out));

	reg [0:0] andOp_338_in0;
	reg [0:0] andOp_338_in1;
	wire [0:0] andOp_338_out;
	andOp #(.WIDTH(1)) andOp_338(.in0(andOp_338_in0), .in1(andOp_338_in1), .out(andOp_338_out));

	reg [31:0] eq_339_in0;
	reg [31:0] eq_339_in1;
	wire [0:0] eq_339_out;
	eq #(.WIDTH(32)) eq_339(.in0(eq_339_in0), .in1(eq_339_in1), .out(eq_339_out));

	reg [0:0] andOp_340_in0;
	reg [0:0] andOp_340_in1;
	wire [0:0] andOp_340_out;
	andOp #(.WIDTH(1)) andOp_340(.in0(andOp_340_in0), .in1(andOp_340_in1), .out(andOp_340_out));

	reg [0:0] andOp_341_in0;
	reg [0:0] andOp_341_in1;
	wire [0:0] andOp_341_out;
	andOp #(.WIDTH(1)) andOp_341(.in0(andOp_341_in0), .in1(andOp_341_in1), .out(andOp_341_out));

	reg [31:0] eq_342_in0;
	reg [31:0] eq_342_in1;
	wire [0:0] eq_342_out;
	eq #(.WIDTH(32)) eq_342(.in0(eq_342_in0), .in1(eq_342_in1), .out(eq_342_out));

	reg [0:0] andOp_343_in0;
	reg [0:0] andOp_343_in1;
	wire [0:0] andOp_343_out;
	andOp #(.WIDTH(1)) andOp_343(.in0(andOp_343_in0), .in1(andOp_343_in1), .out(andOp_343_out));

	reg [0:0] notOp_344_in0;
	wire [0:0] notOp_344_out;
	notOp #(.WIDTH(1)) notOp_344(.in(notOp_344_in0), .out(notOp_344_out));

	reg [0:0] andOp_345_in0;
	reg [0:0] andOp_345_in1;
	wire [0:0] andOp_345_out;
	andOp #(.WIDTH(1)) andOp_345(.in0(andOp_345_in0), .in1(andOp_345_in1), .out(andOp_345_out));

	reg [0:0] notOp_346_in0;
	wire [0:0] notOp_346_out;
	notOp #(.WIDTH(1)) notOp_346(.in(notOp_346_in0), .out(notOp_346_out));

	reg [0:0] andOp_347_in0;
	reg [0:0] andOp_347_in1;
	wire [0:0] andOp_347_out;
	andOp #(.WIDTH(1)) andOp_347(.in0(andOp_347_in0), .in1(andOp_347_in1), .out(andOp_347_out));

	reg [0:0] notOp_348_in0;
	wire [0:0] notOp_348_out;
	notOp #(.WIDTH(1)) notOp_348(.in(notOp_348_in0), .out(notOp_348_out));

	reg [0:0] andOp_349_in0;
	reg [0:0] andOp_349_in1;
	wire [0:0] andOp_349_out;
	andOp #(.WIDTH(1)) andOp_349(.in0(andOp_349_in0), .in1(andOp_349_in1), .out(andOp_349_out));

	reg [0:0] andOp_350_in0;
	reg [0:0] andOp_350_in1;
	wire [0:0] andOp_350_out;
	andOp #(.WIDTH(1)) andOp_350(.in0(andOp_350_in0), .in1(andOp_350_in1), .out(andOp_350_out));

	reg [31:0] eq_351_in0;
	reg [31:0] eq_351_in1;
	wire [0:0] eq_351_out;
	eq #(.WIDTH(32)) eq_351(.in0(eq_351_in0), .in1(eq_351_in1), .out(eq_351_out));

	reg [0:0] andOp_352_in0;
	reg [0:0] andOp_352_in1;
	wire [0:0] andOp_352_out;
	andOp #(.WIDTH(1)) andOp_352(.in0(andOp_352_in0), .in1(andOp_352_in1), .out(andOp_352_out));

	reg [0:0] notOp_353_in0;
	wire [0:0] notOp_353_out;
	notOp #(.WIDTH(1)) notOp_353(.in(notOp_353_in0), .out(notOp_353_out));

	reg [0:0] andOp_354_in0;
	reg [0:0] andOp_354_in1;
	wire [0:0] andOp_354_out;
	andOp #(.WIDTH(1)) andOp_354(.in0(andOp_354_in0), .in1(andOp_354_in1), .out(andOp_354_out));

	reg [0:0] notOp_355_in0;
	wire [0:0] notOp_355_out;
	notOp #(.WIDTH(1)) notOp_355(.in(notOp_355_in0), .out(notOp_355_out));

	reg [0:0] andOp_356_in0;
	reg [0:0] andOp_356_in1;
	wire [0:0] andOp_356_out;
	andOp #(.WIDTH(1)) andOp_356(.in0(andOp_356_in0), .in1(andOp_356_in1), .out(andOp_356_out));

	reg [0:0] notOp_357_in0;
	wire [0:0] notOp_357_out;
	notOp #(.WIDTH(1)) notOp_357(.in(notOp_357_in0), .out(notOp_357_out));

	reg [0:0] andOp_358_in0;
	reg [0:0] andOp_358_in1;
	wire [0:0] andOp_358_out;
	andOp #(.WIDTH(1)) andOp_358(.in0(andOp_358_in0), .in1(andOp_358_in1), .out(andOp_358_out));

	reg [0:0] andOp_359_in0;
	reg [0:0] andOp_359_in1;
	wire [0:0] andOp_359_out;
	andOp #(.WIDTH(1)) andOp_359(.in0(andOp_359_in0), .in1(andOp_359_in1), .out(andOp_359_out));

	reg [31:0] eq_360_in0;
	reg [31:0] eq_360_in1;
	wire [0:0] eq_360_out;
	eq #(.WIDTH(32)) eq_360(.in0(eq_360_in0), .in1(eq_360_in1), .out(eq_360_out));

	reg [0:0] andOp_361_in0;
	reg [0:0] andOp_361_in1;
	wire [0:0] andOp_361_out;
	andOp #(.WIDTH(1)) andOp_361(.in0(andOp_361_in0), .in1(andOp_361_in1), .out(andOp_361_out));

	reg [0:0] notOp_362_in0;
	wire [0:0] notOp_362_out;
	notOp #(.WIDTH(1)) notOp_362(.in(notOp_362_in0), .out(notOp_362_out));

	reg [0:0] andOp_363_in0;
	reg [0:0] andOp_363_in1;
	wire [0:0] andOp_363_out;
	andOp #(.WIDTH(1)) andOp_363(.in0(andOp_363_in0), .in1(andOp_363_in1), .out(andOp_363_out));

	reg [0:0] notOp_364_in0;
	wire [0:0] notOp_364_out;
	notOp #(.WIDTH(1)) notOp_364(.in(notOp_364_in0), .out(notOp_364_out));

	reg [0:0] andOp_365_in0;
	reg [0:0] andOp_365_in1;
	wire [0:0] andOp_365_out;
	andOp #(.WIDTH(1)) andOp_365(.in0(andOp_365_in0), .in1(andOp_365_in1), .out(andOp_365_out));

	reg [0:0] notOp_366_in0;
	wire [0:0] notOp_366_out;
	notOp #(.WIDTH(1)) notOp_366(.in(notOp_366_in0), .out(notOp_366_out));

	reg [0:0] andOp_367_in0;
	reg [0:0] andOp_367_in1;
	wire [0:0] andOp_367_out;
	andOp #(.WIDTH(1)) andOp_367(.in0(andOp_367_in0), .in1(andOp_367_in1), .out(andOp_367_out));

	// End Functional Units

	reg [31:0] add_tmp_5;
	reg [31:0] call_tmp_2;
	reg [31:0] data_store_0_0;
	reg [31:0] data_store_0_2;
	reg [0:0] data_store_0_4;
	reg [0:0] data_store_1_10;
	reg [31:0] data_store_1_6;
	reg [31:0] data_store_1_8;
	reg [31:0] data_store_2_12;
	reg [31:0] data_store_2_14;
	reg [0:0] data_store_2_16;
	reg [31:0] data_store_3_18;
	reg [31:0] data_store_3_20;
	reg [0:0] data_store_3_22;
	reg [31:0] data_store_4_24;
	reg [31:0] data_store_4_26;
	reg [0:0] data_store_4_28;
	reg [31:0] global_state;
	reg [0:0] icmp_tmp_6;
	reg [31:0] phi_tmp_1;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_3_last_state;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;
	reg [31:0] state_4_last_state;

	// controller for add_add_14.add_in0_add_14
	// controller for add_add_14.add_in1_add_14
	// Insensitive connections
	always @(*) begin
		add_in0_add_14 = valid ? rdata_ram_0 : rdata_ram_0;
		add_in1_add_14 = valid ? tmp_output_150_out_data : tmp_output_150_out_data;
	end
	// controller for add_add_16.add_in0_add_16
	// controller for add_add_16.add_in1_add_16
	// Insensitive connections
	always @(*) begin
		add_in0_add_16 = valid ? data_in_3_19_out_data : data_in_3_19_out_data;
		add_in1_add_16 = valid ? 32'd1 : 32'd1;
	end
	// controller for andOp_108.andOp_108_in0
	// controller for andOp_108.andOp_108_in1
	// Insensitive connections
	always @(*) begin
		andOp_108_in0 = valid ? notOp_107_out : notOp_107_out;
		andOp_108_in1 = valid ? andOp_31_out : andOp_31_out;
	end
	// controller for andOp_111.andOp_111_in0
	// controller for andOp_111.andOp_111_in1
	// Insensitive connections
	always @(*) begin
		andOp_111_in0 = valid ? notOp_110_out : notOp_110_out;
		andOp_111_in1 = valid ? andOp_46_out : andOp_46_out;
	end
	// controller for andOp_114.andOp_114_in0
	// controller for andOp_114.andOp_114_in1
	// Insensitive connections
	always @(*) begin
		andOp_114_in0 = valid ? notOp_113_out : notOp_113_out;
		andOp_114_in1 = valid ? andOp_37_out : andOp_37_out;
	end
	// controller for andOp_118.andOp_118_in0
	// controller for andOp_118.andOp_118_in1
	// Insensitive connections
	always @(*) begin
		andOp_118_in0 = valid ? notOp_117_out : notOp_117_out;
		andOp_118_in1 = valid ? andOp_49_out : andOp_49_out;
	end
	// controller for andOp_122.andOp_122_in0
	// controller for andOp_122.andOp_122_in1
	// Insensitive connections
	always @(*) begin
		andOp_122_in0 = valid ? notOp_121_out : notOp_121_out;
		andOp_122_in1 = valid ? andOp_73_out : andOp_73_out;
	end
	// controller for andOp_125.andOp_125_in0
	// controller for andOp_125.andOp_125_in1
	// Insensitive connections
	always @(*) begin
		andOp_125_in0 = valid ? notOp_124_out : notOp_124_out;
		andOp_125_in1 = valid ? andOp_61_out : andOp_61_out;
	end
	// controller for andOp_128.andOp_128_in0
	// controller for andOp_128.andOp_128_in1
	// Insensitive connections
	always @(*) begin
		andOp_128_in0 = valid ? notOp_127_out : notOp_127_out;
		andOp_128_in1 = valid ? andOp_66_out : andOp_66_out;
	end
	// controller for andOp_131.andOp_131_in0
	// controller for andOp_131.andOp_131_in1
	// Insensitive connections
	always @(*) begin
		andOp_131_in0 = valid ? notOp_130_out : notOp_130_out;
		andOp_131_in1 = valid ? andOp_70_out : andOp_70_out;
	end
	// controller for andOp_134.andOp_134_in0
	// controller for andOp_134.andOp_134_in1
	// Insensitive connections
	always @(*) begin
		andOp_134_in0 = valid ? notOp_133_out : notOp_133_out;
		andOp_134_in1 = valid ? andOp_54_out : andOp_54_out;
	end
	// controller for andOp_136.andOp_136_in0
	// controller for andOp_136.andOp_136_in1
	// Insensitive connections
	always @(*) begin
		andOp_136_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_136_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_137.andOp_137_in0
	// controller for andOp_137.andOp_137_in1
	// Insensitive connections
	always @(*) begin
		andOp_137_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_137_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_138.andOp_138_in0
	// controller for andOp_138.andOp_138_in1
	// Insensitive connections
	always @(*) begin
		andOp_138_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_138_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_139.andOp_139_in0
	// controller for andOp_139.andOp_139_in1
	// Insensitive connections
	always @(*) begin
		andOp_139_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_139_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_140.andOp_140_in0
	// controller for andOp_140.andOp_140_in1
	// Insensitive connections
	always @(*) begin
		andOp_140_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_140_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_141.andOp_141_in0
	// controller for andOp_141.andOp_141_in1
	// Insensitive connections
	always @(*) begin
		andOp_141_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_141_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_142.andOp_142_in0
	// controller for andOp_142.andOp_142_in1
	// Insensitive connections
	always @(*) begin
		andOp_142_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_142_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_143.andOp_143_in0
	// controller for andOp_143.andOp_143_in1
	// Insensitive connections
	always @(*) begin
		andOp_143_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
		andOp_143_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_144.andOp_144_in0
	// controller for andOp_144.andOp_144_in1
	// Insensitive connections
	always @(*) begin
		andOp_144_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_144_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_145.andOp_145_in0
	// controller for andOp_145.andOp_145_in1
	// Insensitive connections
	always @(*) begin
		andOp_145_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_145_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_146.andOp_146_in0
	// controller for andOp_146.andOp_146_in1
	// Insensitive connections
	always @(*) begin
		andOp_146_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_146_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_149.andOp_149_in0
	// controller for andOp_149.andOp_149_in1
	// Insensitive connections
	always @(*) begin
		andOp_149_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_149_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_152.andOp_152_in0
	// controller for andOp_152.andOp_152_in1
	// Insensitive connections
	always @(*) begin
		andOp_152_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_152_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_153.andOp_153_in0
	// controller for andOp_153.andOp_153_in1
	// Insensitive connections
	always @(*) begin
		andOp_153_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_153_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_154.andOp_154_in0
	// controller for andOp_154.andOp_154_in1
	// Insensitive connections
	always @(*) begin
		andOp_154_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_154_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_155.andOp_155_in0
	// controller for andOp_155.andOp_155_in1
	// Insensitive connections
	always @(*) begin
		andOp_155_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_155_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_156.andOp_156_in0
	// controller for andOp_156.andOp_156_in1
	// Insensitive connections
	always @(*) begin
		andOp_156_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
		andOp_156_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_157.andOp_157_in0
	// controller for andOp_157.andOp_157_in1
	// Insensitive connections
	always @(*) begin
		andOp_157_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_157_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_158.andOp_158_in0
	// controller for andOp_158.andOp_158_in1
	// Insensitive connections
	always @(*) begin
		andOp_158_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_158_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_159.andOp_159_in0
	// controller for andOp_159.andOp_159_in1
	// Insensitive connections
	always @(*) begin
		andOp_159_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_159_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_160.andOp_160_in0
	// controller for andOp_160.andOp_160_in1
	// Insensitive connections
	always @(*) begin
		andOp_160_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_160_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_161.andOp_161_in0
	// controller for andOp_161.andOp_161_in1
	// Insensitive connections
	always @(*) begin
		andOp_161_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_161_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_162.andOp_162_in0
	// controller for andOp_162.andOp_162_in1
	// Insensitive connections
	always @(*) begin
		andOp_162_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_162_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_164.andOp_164_in0
	// controller for andOp_164.andOp_164_in1
	// Insensitive connections
	always @(*) begin
		andOp_164_in0 = valid ? notOp_163_out : notOp_163_out;
		andOp_164_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_166.andOp_166_in0
	// controller for andOp_166.andOp_166_in1
	// Insensitive connections
	always @(*) begin
		andOp_166_in0 = valid ? notOp_165_out : notOp_165_out;
		andOp_166_in1 = valid ? andOp_164_out : andOp_164_out;
	end
	// controller for andOp_168.andOp_168_in0
	// controller for andOp_168.andOp_168_in1
	// Insensitive connections
	always @(*) begin
		andOp_168_in0 = valid ? notOp_167_out : notOp_167_out;
		andOp_168_in1 = valid ? andOp_166_out : andOp_166_out;
	end
	// controller for andOp_170.andOp_170_in0
	// controller for andOp_170.andOp_170_in1
	// Insensitive connections
	always @(*) begin
		andOp_170_in0 = valid ? notOp_169_out : notOp_169_out;
		andOp_170_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_172.andOp_172_in0
	// controller for andOp_172.andOp_172_in1
	// Insensitive connections
	always @(*) begin
		andOp_172_in0 = valid ? notOp_171_out : notOp_171_out;
		andOp_172_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_174.andOp_174_in0
	// controller for andOp_174.andOp_174_in1
	// Insensitive connections
	always @(*) begin
		andOp_174_in0 = valid ? notOp_173_out : notOp_173_out;
		andOp_174_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_176.andOp_176_in0
	// controller for andOp_176.andOp_176_in1
	// Insensitive connections
	always @(*) begin
		andOp_176_in0 = valid ? notOp_175_out : notOp_175_out;
		andOp_176_in1 = valid ? andOp_174_out : andOp_174_out;
	end
	// controller for andOp_178.andOp_178_in0
	// controller for andOp_178.andOp_178_in1
	// Insensitive connections
	always @(*) begin
		andOp_178_in0 = valid ? notOp_177_out : notOp_177_out;
		andOp_178_in1 = valid ? andOp_176_out : andOp_176_out;
	end
	// controller for andOp_179.andOp_179_in0
	// controller for andOp_179.andOp_179_in1
	// Insensitive connections
	always @(*) begin
		andOp_179_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_179_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_180.andOp_180_in0
	// controller for andOp_180.andOp_180_in1
	// Insensitive connections
	always @(*) begin
		andOp_180_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_180_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_181.andOp_181_in0
	// controller for andOp_181.andOp_181_in1
	// Insensitive connections
	always @(*) begin
		andOp_181_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_181_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_182.andOp_182_in0
	// controller for andOp_182.andOp_182_in1
	// Insensitive connections
	always @(*) begin
		andOp_182_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_182_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_184.andOp_184_in0
	// controller for andOp_184.andOp_184_in1
	// Insensitive connections
	always @(*) begin
		andOp_184_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_184_in1 = valid ? eq_183_out : eq_183_out;
	end
	// controller for andOp_186.andOp_186_in0
	// controller for andOp_186.andOp_186_in1
	// Insensitive connections
	always @(*) begin
		andOp_186_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_186_in1 = valid ? eq_185_out : eq_185_out;
	end
	// controller for andOp_188.andOp_188_in0
	// controller for andOp_188.andOp_188_in1
	// Insensitive connections
	always @(*) begin
		andOp_188_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_188_in1 = valid ? eq_187_out : eq_187_out;
	end
	// controller for andOp_190.andOp_190_in0
	// controller for andOp_190.andOp_190_in1
	// Insensitive connections
	always @(*) begin
		andOp_190_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_190_in1 = valid ? eq_189_out : eq_189_out;
	end
	// controller for andOp_192.andOp_192_in0
	// controller for andOp_192.andOp_192_in1
	// Insensitive connections
	always @(*) begin
		andOp_192_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_192_in1 = valid ? eq_191_out : eq_191_out;
	end
	// controller for andOp_193.andOp_193_in0
	// controller for andOp_193.andOp_193_in1
	// Insensitive connections
	always @(*) begin
		andOp_193_in0 = valid ? 1'd0 : 1'd0;
		andOp_193_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_195.andOp_195_in0
	// controller for andOp_195.andOp_195_in1
	// Insensitive connections
	always @(*) begin
		andOp_195_in0 = valid ? andOp_193_out : andOp_193_out;
		andOp_195_in1 = valid ? eq_194_out : eq_194_out;
	end
	// controller for andOp_197.andOp_197_in0
	// controller for andOp_197.andOp_197_in1
	// Insensitive connections
	always @(*) begin
		andOp_197_in0 = valid ? andOp_193_out : andOp_193_out;
		andOp_197_in1 = valid ? notOp_196_out : notOp_196_out;
	end
	// controller for andOp_199.andOp_199_in0
	// controller for andOp_199.andOp_199_in1
	// Insensitive connections
	always @(*) begin
		andOp_199_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_199_in1 = valid ? notOp_198_out : notOp_198_out;
	end
	// controller for andOp_201.andOp_201_in0
	// controller for andOp_201.andOp_201_in1
	// Insensitive connections
	always @(*) begin
		andOp_201_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_201_in1 = valid ? notOp_200_out : notOp_200_out;
	end
	// controller for andOp_202.andOp_202_in0
	// controller for andOp_202.andOp_202_in1
	// Insensitive connections
	always @(*) begin
		andOp_202_in0 = valid ? 1'd0 : 1'd0;
		andOp_202_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_204.andOp_204_in0
	// controller for andOp_204.andOp_204_in1
	// Insensitive connections
	always @(*) begin
		andOp_204_in0 = valid ? andOp_202_out : andOp_202_out;
		andOp_204_in1 = valid ? eq_203_out : eq_203_out;
	end
	// controller for andOp_206.andOp_206_in0
	// controller for andOp_206.andOp_206_in1
	// Insensitive connections
	always @(*) begin
		andOp_206_in0 = valid ? andOp_202_out : andOp_202_out;
		andOp_206_in1 = valid ? notOp_205_out : notOp_205_out;
	end
	// controller for andOp_208.andOp_208_in0
	// controller for andOp_208.andOp_208_in1
	// Insensitive connections
	always @(*) begin
		andOp_208_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_208_in1 = valid ? notOp_207_out : notOp_207_out;
	end
	// controller for andOp_210.andOp_210_in0
	// controller for andOp_210.andOp_210_in1
	// Insensitive connections
	always @(*) begin
		andOp_210_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_210_in1 = valid ? notOp_209_out : notOp_209_out;
	end
	// controller for andOp_211.andOp_211_in0
	// controller for andOp_211.andOp_211_in1
	// Insensitive connections
	always @(*) begin
		andOp_211_in0 = valid ? 1'd0 : 1'd0;
		andOp_211_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_213.andOp_213_in0
	// controller for andOp_213.andOp_213_in1
	// Insensitive connections
	always @(*) begin
		andOp_213_in0 = valid ? andOp_211_out : andOp_211_out;
		andOp_213_in1 = valid ? eq_212_out : eq_212_out;
	end
	// controller for andOp_215.andOp_215_in0
	// controller for andOp_215.andOp_215_in1
	// Insensitive connections
	always @(*) begin
		andOp_215_in0 = valid ? andOp_211_out : andOp_211_out;
		andOp_215_in1 = valid ? notOp_214_out : notOp_214_out;
	end
	// controller for andOp_217.andOp_217_in0
	// controller for andOp_217.andOp_217_in1
	// Insensitive connections
	always @(*) begin
		andOp_217_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_217_in1 = valid ? notOp_216_out : notOp_216_out;
	end
	// controller for andOp_219.andOp_219_in0
	// controller for andOp_219.andOp_219_in1
	// Insensitive connections
	always @(*) begin
		andOp_219_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_219_in1 = valid ? notOp_218_out : notOp_218_out;
	end
	// controller for andOp_221.andOp_221_in0
	// controller for andOp_221.andOp_221_in1
	// Insensitive connections
	always @(*) begin
		andOp_221_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_221_in1 = valid ? eq_220_out : eq_220_out;
	end
	// controller for andOp_223.andOp_223_in0
	// controller for andOp_223.andOp_223_in1
	// Insensitive connections
	always @(*) begin
		andOp_223_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_223_in1 = valid ? eq_222_out : eq_222_out;
	end
	// controller for andOp_225.andOp_225_in0
	// controller for andOp_225.andOp_225_in1
	// Insensitive connections
	always @(*) begin
		andOp_225_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_225_in1 = valid ? eq_224_out : eq_224_out;
	end
	// controller for andOp_227.andOp_227_in0
	// controller for andOp_227.andOp_227_in1
	// Insensitive connections
	always @(*) begin
		andOp_227_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_227_in1 = valid ? eq_226_out : eq_226_out;
	end
	// controller for andOp_229.andOp_229_in0
	// controller for andOp_229.andOp_229_in1
	// Insensitive connections
	always @(*) begin
		andOp_229_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_229_in1 = valid ? eq_228_out : eq_228_out;
	end
	// controller for andOp_230.andOp_230_in0
	// controller for andOp_230.andOp_230_in1
	// Insensitive connections
	always @(*) begin
		andOp_230_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_230_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_232.andOp_232_in0
	// controller for andOp_232.andOp_232_in1
	// Insensitive connections
	always @(*) begin
		andOp_232_in0 = valid ? andOp_230_out : andOp_230_out;
		andOp_232_in1 = valid ? eq_231_out : eq_231_out;
	end
	// controller for andOp_234.andOp_234_in0
	// controller for andOp_234.andOp_234_in1
	// Insensitive connections
	always @(*) begin
		andOp_234_in0 = valid ? andOp_230_out : andOp_230_out;
		andOp_234_in1 = valid ? notOp_233_out : notOp_233_out;
	end
	// controller for andOp_236.andOp_236_in0
	// controller for andOp_236.andOp_236_in1
	// Insensitive connections
	always @(*) begin
		andOp_236_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_236_in1 = valid ? notOp_235_out : notOp_235_out;
	end
	// controller for andOp_238.andOp_238_in0
	// controller for andOp_238.andOp_238_in1
	// Insensitive connections
	always @(*) begin
		andOp_238_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_238_in1 = valid ? notOp_237_out : notOp_237_out;
	end
	// controller for andOp_239.andOp_239_in0
	// controller for andOp_239.andOp_239_in1
	// Insensitive connections
	always @(*) begin
		andOp_239_in0 = valid ? 1'd0 : 1'd0;
		andOp_239_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_241.andOp_241_in0
	// controller for andOp_241.andOp_241_in1
	// Insensitive connections
	always @(*) begin
		andOp_241_in0 = valid ? andOp_239_out : andOp_239_out;
		andOp_241_in1 = valid ? eq_240_out : eq_240_out;
	end
	// controller for andOp_243.andOp_243_in0
	// controller for andOp_243.andOp_243_in1
	// Insensitive connections
	always @(*) begin
		andOp_243_in0 = valid ? andOp_239_out : andOp_239_out;
		andOp_243_in1 = valid ? notOp_242_out : notOp_242_out;
	end
	// controller for andOp_245.andOp_245_in0
	// controller for andOp_245.andOp_245_in1
	// Insensitive connections
	always @(*) begin
		andOp_245_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_245_in1 = valid ? notOp_244_out : notOp_244_out;
	end
	// controller for andOp_247.andOp_247_in0
	// controller for andOp_247.andOp_247_in1
	// Insensitive connections
	always @(*) begin
		andOp_247_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_247_in1 = valid ? notOp_246_out : notOp_246_out;
	end
	// controller for andOp_248.andOp_248_in0
	// controller for andOp_248.andOp_248_in1
	// Insensitive connections
	always @(*) begin
		andOp_248_in0 = valid ? 1'd0 : 1'd0;
		andOp_248_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_250.andOp_250_in0
	// controller for andOp_250.andOp_250_in1
	// Insensitive connections
	always @(*) begin
		andOp_250_in0 = valid ? andOp_248_out : andOp_248_out;
		andOp_250_in1 = valid ? eq_249_out : eq_249_out;
	end
	// controller for andOp_252.andOp_252_in0
	// controller for andOp_252.andOp_252_in1
	// Insensitive connections
	always @(*) begin
		andOp_252_in0 = valid ? andOp_248_out : andOp_248_out;
		andOp_252_in1 = valid ? notOp_251_out : notOp_251_out;
	end
	// controller for andOp_254.andOp_254_in0
	// controller for andOp_254.andOp_254_in1
	// Insensitive connections
	always @(*) begin
		andOp_254_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_254_in1 = valid ? notOp_253_out : notOp_253_out;
	end
	// controller for andOp_256.andOp_256_in0
	// controller for andOp_256.andOp_256_in1
	// Insensitive connections
	always @(*) begin
		andOp_256_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_256_in1 = valid ? notOp_255_out : notOp_255_out;
	end
	// controller for andOp_258.andOp_258_in0
	// controller for andOp_258.andOp_258_in1
	// Insensitive connections
	always @(*) begin
		andOp_258_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_258_in1 = valid ? eq_257_out : eq_257_out;
	end
	// controller for andOp_260.andOp_260_in0
	// controller for andOp_260.andOp_260_in1
	// Insensitive connections
	always @(*) begin
		andOp_260_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_260_in1 = valid ? eq_259_out : eq_259_out;
	end
	// controller for andOp_262.andOp_262_in0
	// controller for andOp_262.andOp_262_in1
	// Insensitive connections
	always @(*) begin
		andOp_262_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_262_in1 = valid ? eq_261_out : eq_261_out;
	end
	// controller for andOp_264.andOp_264_in0
	// controller for andOp_264.andOp_264_in1
	// Insensitive connections
	always @(*) begin
		andOp_264_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_264_in1 = valid ? eq_263_out : eq_263_out;
	end
	// controller for andOp_266.andOp_266_in0
	// controller for andOp_266.andOp_266_in1
	// Insensitive connections
	always @(*) begin
		andOp_266_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_266_in1 = valid ? eq_265_out : eq_265_out;
	end
	// controller for andOp_267.andOp_267_in0
	// controller for andOp_267.andOp_267_in1
	// Insensitive connections
	always @(*) begin
		andOp_267_in0 = valid ? 1'd0 : 1'd0;
		andOp_267_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_269.andOp_269_in0
	// controller for andOp_269.andOp_269_in1
	// Insensitive connections
	always @(*) begin
		andOp_269_in0 = valid ? andOp_267_out : andOp_267_out;
		andOp_269_in1 = valid ? eq_268_out : eq_268_out;
	end
	// controller for andOp_271.andOp_271_in0
	// controller for andOp_271.andOp_271_in1
	// Insensitive connections
	always @(*) begin
		andOp_271_in0 = valid ? andOp_267_out : andOp_267_out;
		andOp_271_in1 = valid ? notOp_270_out : notOp_270_out;
	end
	// controller for andOp_273.andOp_273_in0
	// controller for andOp_273.andOp_273_in1
	// Insensitive connections
	always @(*) begin
		andOp_273_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_273_in1 = valid ? notOp_272_out : notOp_272_out;
	end
	// controller for andOp_275.andOp_275_in0
	// controller for andOp_275.andOp_275_in1
	// Insensitive connections
	always @(*) begin
		andOp_275_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_275_in1 = valid ? notOp_274_out : notOp_274_out;
	end
	// controller for andOp_276.andOp_276_in0
	// controller for andOp_276.andOp_276_in1
	// Insensitive connections
	always @(*) begin
		andOp_276_in0 = valid ? 1'd0 : 1'd0;
		andOp_276_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_278.andOp_278_in0
	// controller for andOp_278.andOp_278_in1
	// Insensitive connections
	always @(*) begin
		andOp_278_in0 = valid ? andOp_276_out : andOp_276_out;
		andOp_278_in1 = valid ? eq_277_out : eq_277_out;
	end
	// controller for andOp_280.andOp_280_in0
	// controller for andOp_280.andOp_280_in1
	// Insensitive connections
	always @(*) begin
		andOp_280_in0 = valid ? andOp_276_out : andOp_276_out;
		andOp_280_in1 = valid ? notOp_279_out : notOp_279_out;
	end
	// controller for andOp_282.andOp_282_in0
	// controller for andOp_282.andOp_282_in1
	// Insensitive connections
	always @(*) begin
		andOp_282_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_282_in1 = valid ? notOp_281_out : notOp_281_out;
	end
	// controller for andOp_284.andOp_284_in0
	// controller for andOp_284.andOp_284_in1
	// Insensitive connections
	always @(*) begin
		andOp_284_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_284_in1 = valid ? notOp_283_out : notOp_283_out;
	end
	// controller for andOp_285.andOp_285_in0
	// controller for andOp_285.andOp_285_in1
	// Insensitive connections
	always @(*) begin
		andOp_285_in0 = valid ? 1'd0 : 1'd0;
		andOp_285_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_287.andOp_287_in0
	// controller for andOp_287.andOp_287_in1
	// Insensitive connections
	always @(*) begin
		andOp_287_in0 = valid ? andOp_285_out : andOp_285_out;
		andOp_287_in1 = valid ? eq_286_out : eq_286_out;
	end
	// controller for andOp_289.andOp_289_in0
	// controller for andOp_289.andOp_289_in1
	// Insensitive connections
	always @(*) begin
		andOp_289_in0 = valid ? andOp_285_out : andOp_285_out;
		andOp_289_in1 = valid ? notOp_288_out : notOp_288_out;
	end
	// controller for andOp_291.andOp_291_in0
	// controller for andOp_291.andOp_291_in1
	// Insensitive connections
	always @(*) begin
		andOp_291_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_291_in1 = valid ? notOp_290_out : notOp_290_out;
	end
	// controller for andOp_293.andOp_293_in0
	// controller for andOp_293.andOp_293_in1
	// Insensitive connections
	always @(*) begin
		andOp_293_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_293_in1 = valid ? notOp_292_out : notOp_292_out;
	end
	// controller for andOp_295.andOp_295_in0
	// controller for andOp_295.andOp_295_in1
	// Insensitive connections
	always @(*) begin
		andOp_295_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_295_in1 = valid ? eq_294_out : eq_294_out;
	end
	// controller for andOp_297.andOp_297_in0
	// controller for andOp_297.andOp_297_in1
	// Insensitive connections
	always @(*) begin
		andOp_297_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_297_in1 = valid ? eq_296_out : eq_296_out;
	end
	// controller for andOp_299.andOp_299_in0
	// controller for andOp_299.andOp_299_in1
	// Insensitive connections
	always @(*) begin
		andOp_299_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_299_in1 = valid ? eq_298_out : eq_298_out;
	end
	// controller for andOp_30.andOp_30_in0
	// controller for andOp_30.andOp_30_in1
	// Insensitive connections
	always @(*) begin
		andOp_30_in0 = valid ? bb_0_active_in_state_1_out_data : bb_0_active_in_state_1_out_data;
		andOp_30_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_301.andOp_301_in0
	// controller for andOp_301.andOp_301_in1
	// Insensitive connections
	always @(*) begin
		andOp_301_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_301_in1 = valid ? eq_300_out : eq_300_out;
	end
	// controller for andOp_303.andOp_303_in0
	// controller for andOp_303.andOp_303_in1
	// Insensitive connections
	always @(*) begin
		andOp_303_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_303_in1 = valid ? eq_302_out : eq_302_out;
	end
	// controller for andOp_304.andOp_304_in0
	// controller for andOp_304.andOp_304_in1
	// Insensitive connections
	always @(*) begin
		andOp_304_in0 = valid ? 1'd0 : 1'd0;
		andOp_304_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_306.andOp_306_in0
	// controller for andOp_306.andOp_306_in1
	// Insensitive connections
	always @(*) begin
		andOp_306_in0 = valid ? andOp_304_out : andOp_304_out;
		andOp_306_in1 = valid ? eq_305_out : eq_305_out;
	end
	// controller for andOp_308.andOp_308_in0
	// controller for andOp_308.andOp_308_in1
	// Insensitive connections
	always @(*) begin
		andOp_308_in0 = valid ? andOp_304_out : andOp_304_out;
		andOp_308_in1 = valid ? notOp_307_out : notOp_307_out;
	end
	// controller for andOp_31.andOp_31_in0
	// controller for andOp_31.andOp_31_in1
	// Insensitive connections
	always @(*) begin
		andOp_31_in0 = valid ? andOp_30_out : andOp_30_out;
		andOp_31_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_310.andOp_310_in0
	// controller for andOp_310.andOp_310_in1
	// Insensitive connections
	always @(*) begin
		andOp_310_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_310_in1 = valid ? notOp_309_out : notOp_309_out;
	end
	// controller for andOp_312.andOp_312_in0
	// controller for andOp_312.andOp_312_in1
	// Insensitive connections
	always @(*) begin
		andOp_312_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_312_in1 = valid ? notOp_311_out : notOp_311_out;
	end
	// controller for andOp_313.andOp_313_in0
	// controller for andOp_313.andOp_313_in1
	// Insensitive connections
	always @(*) begin
		andOp_313_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_313_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_315.andOp_315_in0
	// controller for andOp_315.andOp_315_in1
	// Insensitive connections
	always @(*) begin
		andOp_315_in0 = valid ? andOp_313_out : andOp_313_out;
		andOp_315_in1 = valid ? eq_314_out : eq_314_out;
	end
	// controller for andOp_317.andOp_317_in0
	// controller for andOp_317.andOp_317_in1
	// Insensitive connections
	always @(*) begin
		andOp_317_in0 = valid ? andOp_313_out : andOp_313_out;
		andOp_317_in1 = valid ? notOp_316_out : notOp_316_out;
	end
	// controller for andOp_319.andOp_319_in0
	// controller for andOp_319.andOp_319_in1
	// Insensitive connections
	always @(*) begin
		andOp_319_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_319_in1 = valid ? notOp_318_out : notOp_318_out;
	end
	// controller for andOp_321.andOp_321_in0
	// controller for andOp_321.andOp_321_in1
	// Insensitive connections
	always @(*) begin
		andOp_321_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_321_in1 = valid ? notOp_320_out : notOp_320_out;
	end
	// controller for andOp_322.andOp_322_in0
	// controller for andOp_322.andOp_322_in1
	// Insensitive connections
	always @(*) begin
		andOp_322_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_322_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_324.andOp_324_in0
	// controller for andOp_324.andOp_324_in1
	// Insensitive connections
	always @(*) begin
		andOp_324_in0 = valid ? andOp_322_out : andOp_322_out;
		andOp_324_in1 = valid ? eq_323_out : eq_323_out;
	end
	// controller for andOp_326.andOp_326_in0
	// controller for andOp_326.andOp_326_in1
	// Insensitive connections
	always @(*) begin
		andOp_326_in0 = valid ? andOp_322_out : andOp_322_out;
		andOp_326_in1 = valid ? notOp_325_out : notOp_325_out;
	end
	// controller for andOp_328.andOp_328_in0
	// controller for andOp_328.andOp_328_in1
	// Insensitive connections
	always @(*) begin
		andOp_328_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_328_in1 = valid ? notOp_327_out : notOp_327_out;
	end
	// controller for andOp_33.andOp_33_in0
	// controller for andOp_33.andOp_33_in1
	// Insensitive connections
	always @(*) begin
		andOp_33_in0 = valid ? bb_0_active_in_state_1_out_data : bb_0_active_in_state_1_out_data;
		andOp_33_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_330.andOp_330_in0
	// controller for andOp_330.andOp_330_in1
	// Insensitive connections
	always @(*) begin
		andOp_330_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_330_in1 = valid ? notOp_329_out : notOp_329_out;
	end
	// controller for andOp_332.andOp_332_in0
	// controller for andOp_332.andOp_332_in1
	// Insensitive connections
	always @(*) begin
		andOp_332_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_332_in1 = valid ? eq_331_out : eq_331_out;
	end
	// controller for andOp_334.andOp_334_in0
	// controller for andOp_334.andOp_334_in1
	// Insensitive connections
	always @(*) begin
		andOp_334_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_334_in1 = valid ? eq_333_out : eq_333_out;
	end
	// controller for andOp_336.andOp_336_in0
	// controller for andOp_336.andOp_336_in1
	// Insensitive connections
	always @(*) begin
		andOp_336_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_336_in1 = valid ? eq_335_out : eq_335_out;
	end
	// controller for andOp_338.andOp_338_in0
	// controller for andOp_338.andOp_338_in1
	// Insensitive connections
	always @(*) begin
		andOp_338_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_338_in1 = valid ? eq_337_out : eq_337_out;
	end
	// controller for andOp_34.andOp_34_in0
	// controller for andOp_34.andOp_34_in1
	// Insensitive connections
	always @(*) begin
		andOp_34_in0 = valid ? andOp_33_out : andOp_33_out;
		andOp_34_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_340.andOp_340_in0
	// controller for andOp_340.andOp_340_in1
	// Insensitive connections
	always @(*) begin
		andOp_340_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_340_in1 = valid ? eq_339_out : eq_339_out;
	end
	// controller for andOp_341.andOp_341_in0
	// controller for andOp_341.andOp_341_in1
	// Insensitive connections
	always @(*) begin
		andOp_341_in0 = valid ? 1'd0 : 1'd0;
		andOp_341_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_343.andOp_343_in0
	// controller for andOp_343.andOp_343_in1
	// Insensitive connections
	always @(*) begin
		andOp_343_in0 = valid ? andOp_341_out : andOp_341_out;
		andOp_343_in1 = valid ? eq_342_out : eq_342_out;
	end
	// controller for andOp_345.andOp_345_in0
	// controller for andOp_345.andOp_345_in1
	// Insensitive connections
	always @(*) begin
		andOp_345_in0 = valid ? andOp_341_out : andOp_341_out;
		andOp_345_in1 = valid ? notOp_344_out : notOp_344_out;
	end
	// controller for andOp_347.andOp_347_in0
	// controller for andOp_347.andOp_347_in1
	// Insensitive connections
	always @(*) begin
		andOp_347_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_347_in1 = valid ? notOp_346_out : notOp_346_out;
	end
	// controller for andOp_349.andOp_349_in0
	// controller for andOp_349.andOp_349_in1
	// Insensitive connections
	always @(*) begin
		andOp_349_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_349_in1 = valid ? notOp_348_out : notOp_348_out;
	end
	// controller for andOp_350.andOp_350_in0
	// controller for andOp_350.andOp_350_in1
	// Insensitive connections
	always @(*) begin
		andOp_350_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_350_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_352.andOp_352_in0
	// controller for andOp_352.andOp_352_in1
	// Insensitive connections
	always @(*) begin
		andOp_352_in0 = valid ? andOp_350_out : andOp_350_out;
		andOp_352_in1 = valid ? eq_351_out : eq_351_out;
	end
	// controller for andOp_354.andOp_354_in0
	// controller for andOp_354.andOp_354_in1
	// Insensitive connections
	always @(*) begin
		andOp_354_in0 = valid ? andOp_350_out : andOp_350_out;
		andOp_354_in1 = valid ? notOp_353_out : notOp_353_out;
	end
	// controller for andOp_356.andOp_356_in0
	// controller for andOp_356.andOp_356_in1
	// Insensitive connections
	always @(*) begin
		andOp_356_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_356_in1 = valid ? notOp_355_out : notOp_355_out;
	end
	// controller for andOp_358.andOp_358_in0
	// controller for andOp_358.andOp_358_in1
	// Insensitive connections
	always @(*) begin
		andOp_358_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_358_in1 = valid ? notOp_357_out : notOp_357_out;
	end
	// controller for andOp_359.andOp_359_in0
	// controller for andOp_359.andOp_359_in1
	// Insensitive connections
	always @(*) begin
		andOp_359_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_359_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_36.andOp_36_in0
	// controller for andOp_36.andOp_36_in1
	// Insensitive connections
	always @(*) begin
		andOp_36_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_36_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_361.andOp_361_in0
	// controller for andOp_361.andOp_361_in1
	// Insensitive connections
	always @(*) begin
		andOp_361_in0 = valid ? andOp_359_out : andOp_359_out;
		andOp_361_in1 = valid ? eq_360_out : eq_360_out;
	end
	// controller for andOp_363.andOp_363_in0
	// controller for andOp_363.andOp_363_in1
	// Insensitive connections
	always @(*) begin
		andOp_363_in0 = valid ? andOp_359_out : andOp_359_out;
		andOp_363_in1 = valid ? notOp_362_out : notOp_362_out;
	end
	// controller for andOp_365.andOp_365_in0
	// controller for andOp_365.andOp_365_in1
	// Insensitive connections
	always @(*) begin
		andOp_365_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_365_in1 = valid ? notOp_364_out : notOp_364_out;
	end
	// controller for andOp_367.andOp_367_in0
	// controller for andOp_367.andOp_367_in1
	// Insensitive connections
	always @(*) begin
		andOp_367_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_367_in1 = valid ? notOp_366_out : notOp_366_out;
	end
	// controller for andOp_37.andOp_37_in0
	// controller for andOp_37.andOp_37_in1
	// Insensitive connections
	always @(*) begin
		andOp_37_in0 = valid ? andOp_36_out : andOp_36_out;
		andOp_37_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_39.andOp_39_in0
	// controller for andOp_39.andOp_39_in1
	// Insensitive connections
	always @(*) begin
		andOp_39_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
		andOp_39_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_40.andOp_40_in0
	// controller for andOp_40.andOp_40_in1
	// Insensitive connections
	always @(*) begin
		andOp_40_in0 = valid ? andOp_39_out : andOp_39_out;
		andOp_40_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_42.andOp_42_in0
	// controller for andOp_42.andOp_42_in1
	// Insensitive connections
	always @(*) begin
		andOp_42_in0 = valid ? andOp_40_out : andOp_40_out;
		andOp_42_in1 = valid ? in_read_ready : in_read_ready;
	end
	// controller for andOp_44.andOp_44_in0
	// controller for andOp_44.andOp_44_in1
	// Insensitive connections
	always @(*) begin
		andOp_44_in0 = valid ? andOp_40_out : andOp_40_out;
		andOp_44_in1 = valid ? notOp_43_out : notOp_43_out;
	end
	// controller for andOp_45.andOp_45_in0
	// controller for andOp_45.andOp_45_in1
	// Insensitive connections
	always @(*) begin
		andOp_45_in0 = valid ? bb_8_active_in_state_1_out_data : bb_8_active_in_state_1_out_data;
		andOp_45_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_46.andOp_46_in0
	// controller for andOp_46.andOp_46_in1
	// Insensitive connections
	always @(*) begin
		andOp_46_in0 = valid ? andOp_45_out : andOp_45_out;
		andOp_46_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_48.andOp_48_in0
	// controller for andOp_48.andOp_48_in1
	// Insensitive connections
	always @(*) begin
		andOp_48_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_48_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_49.andOp_49_in0
	// controller for andOp_49.andOp_49_in1
	// Insensitive connections
	always @(*) begin
		andOp_49_in0 = valid ? andOp_48_out : andOp_48_out;
		andOp_49_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_51.andOp_51_in0
	// controller for andOp_51.andOp_51_in1
	// Insensitive connections
	always @(*) begin
		andOp_51_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_51_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_52.andOp_52_in0
	// controller for andOp_52.andOp_52_in1
	// Insensitive connections
	always @(*) begin
		andOp_52_in0 = valid ? andOp_51_out : andOp_51_out;
		andOp_52_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_54.andOp_54_in0
	// controller for andOp_54.andOp_54_in1
	// Insensitive connections
	always @(*) begin
		andOp_54_in0 = valid ? andOp_52_out : andOp_52_out;
		andOp_54_in1 = valid ? data_in_4_29_out_data : data_in_4_29_out_data;
	end
	// controller for andOp_56.andOp_56_in0
	// controller for andOp_56.andOp_56_in1
	// Insensitive connections
	always @(*) begin
		andOp_56_in0 = valid ? andOp_52_out : andOp_52_out;
		andOp_56_in1 = valid ? notOp_55_out : notOp_55_out;
	end
	// controller for andOp_57.andOp_57_in0
	// controller for andOp_57.andOp_57_in1
	// Insensitive connections
	always @(*) begin
		andOp_57_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_57_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_58.andOp_58_in0
	// controller for andOp_58.andOp_58_in1
	// Insensitive connections
	always @(*) begin
		andOp_58_in0 = valid ? andOp_57_out : andOp_57_out;
		andOp_58_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_60.andOp_60_in0
	// controller for andOp_60.andOp_60_in1
	// Insensitive connections
	always @(*) begin
		andOp_60_in0 = valid ? bb_5_active_in_state_4_out_data : bb_5_active_in_state_4_out_data;
		andOp_60_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_61.andOp_61_in0
	// controller for andOp_61.andOp_61_in1
	// Insensitive connections
	always @(*) begin
		andOp_61_in0 = valid ? andOp_60_out : andOp_60_out;
		andOp_61_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_63.andOp_63_in0
	// controller for andOp_63.andOp_63_in1
	// Insensitive connections
	always @(*) begin
		andOp_63_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
		andOp_63_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_64.andOp_64_in0
	// controller for andOp_64.andOp_64_in1
	// Insensitive connections
	always @(*) begin
		andOp_64_in0 = valid ? andOp_63_out : andOp_63_out;
		andOp_64_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_66.andOp_66_in0
	// controller for andOp_66.andOp_66_in1
	// Insensitive connections
	always @(*) begin
		andOp_66_in0 = valid ? andOp_64_out : andOp_64_out;
		andOp_66_in1 = valid ? out_write_ready : out_write_ready;
	end
	// controller for andOp_68.andOp_68_in0
	// controller for andOp_68.andOp_68_in1
	// Insensitive connections
	always @(*) begin
		andOp_68_in0 = valid ? andOp_64_out : andOp_64_out;
		andOp_68_in1 = valid ? notOp_67_out : notOp_67_out;
	end
	// controller for andOp_69.andOp_69_in0
	// controller for andOp_69.andOp_69_in1
	// Insensitive connections
	always @(*) begin
		andOp_69_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_69_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_70.andOp_70_in0
	// controller for andOp_70.andOp_70_in1
	// Insensitive connections
	always @(*) begin
		andOp_70_in0 = valid ? andOp_69_out : andOp_69_out;
		andOp_70_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_72.andOp_72_in0
	// controller for andOp_72.andOp_72_in1
	// Insensitive connections
	always @(*) begin
		andOp_72_in0 = valid ? bb_1_active_in_state_4_out_data : bb_1_active_in_state_4_out_data;
		andOp_72_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_73.andOp_73_in0
	// controller for andOp_73.andOp_73_in1
	// Insensitive connections
	always @(*) begin
		andOp_73_in0 = valid ? andOp_72_out : andOp_72_out;
		andOp_73_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_75.andOp_75_in0
	// controller for andOp_75.andOp_75_in1
	// Insensitive connections
	always @(*) begin
		andOp_75_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_75_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_76.andOp_76_in0
	// controller for andOp_76.andOp_76_in1
	// Insensitive connections
	always @(*) begin
		andOp_76_in0 = valid ? andOp_75_out : andOp_75_out;
		andOp_76_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_78.andOp_78_in0
	// controller for andOp_78.andOp_78_in1
	// Insensitive connections
	always @(*) begin
		andOp_78_in0 = valid ? andOp_76_out : andOp_76_out;
		andOp_78_in1 = valid ? data_in_4_29_out_data : data_in_4_29_out_data;
	end
	// controller for andOp_80.andOp_80_in0
	// controller for andOp_80.andOp_80_in1
	// Insensitive connections
	always @(*) begin
		andOp_80_in0 = valid ? andOp_76_out : andOp_76_out;
		andOp_80_in1 = valid ? notOp_79_out : notOp_79_out;
	end
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_81_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_active_in_state_1.bb_0_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_1_in_data = eq_82_out;
		end else begin
			bb_0_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_104_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_1.bb_0_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_105_out) begin 
			bb_0_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_2.bb_10_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_2_in_data = eq_89_out;
		end else begin
			bb_10_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_3.bb_10_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_3_in_data = eq_92_out;
		end else begin
			bb_10_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_2.bb_10_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_115_out) begin 
			bb_10_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_3.bb_10_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_119_out) begin 
			bb_10_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_4.bb_1_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_4_in_data = orOp_102_out;
		end else begin
			bb_1_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_4.bb_1_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_134_out) begin 
			bb_1_predecessor_in_state_4_in_data = 32'd4;
		end else if (eq_132_out) begin 
			bb_1_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_4.bb_2_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_4_in_data = orOp_100_out;
		end else begin
			bb_2_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_4.bb_2_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_131_out) begin 
			bb_2_predecessor_in_state_4_in_data = 32'd7;
		end else if (eq_129_out) begin 
			bb_2_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_1.bb_3_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_1_in_data = orOp_84_out;
		end else begin
			bb_3_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_1.bb_3_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_108_out) begin 
			bb_3_predecessor_in_state_1_in_data = 32'd0;
		end else if (eq_106_out) begin 
			bb_3_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_3.bb_4_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_3_in_data = orOp_91_out;
		end else begin
			bb_4_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_4.bb_4_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_4_in_data = eq_103_out;
		end else begin
			bb_4_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_3.bb_4_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_118_out) begin 
			bb_4_predecessor_in_state_3_in_data = 32'd10;
		end else if (eq_116_out) begin 
			bb_4_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_4.bb_4_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_135_out) begin 
			bb_4_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_5_active_in_state_4.bb_5_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_5_active_in_state_4_in_data = orOp_94_out;
		end else begin
			bb_5_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_5_predecessor_in_state_4.bb_5_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_122_out) begin 
			bb_5_predecessor_in_state_4_in_data = 32'd1;
		end else if (eq_120_out) begin 
			bb_5_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_5_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_6_active_in_state_4.bb_6_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_6_active_in_state_4_in_data = orOp_96_out;
		end else begin
			bb_6_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_6_predecessor_in_state_4.bb_6_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_125_out) begin 
			bb_6_predecessor_in_state_4_in_data = 32'd5;
		end else if (eq_123_out) begin 
			bb_6_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_6_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_7_active_in_state_4.bb_7_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_7_active_in_state_4_in_data = orOp_98_out;
		end else begin
			bb_7_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_7_predecessor_in_state_4.bb_7_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_128_out) begin 
			bb_7_predecessor_in_state_4_in_data = 32'd6;
		end else if (eq_126_out) begin 
			bb_7_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_7_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_8_active_in_state_1.bb_8_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_state_1_in_data = orOp_88_out;
		end else begin
			bb_8_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_8_predecessor_in_state_1.bb_8_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_114_out) begin 
			bb_8_predecessor_in_state_1_in_data = 32'd3;
		end else if (eq_112_out) begin 
			bb_8_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_8_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_9_active_in_state_1.bb_9_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_9_active_in_state_1_in_data = orOp_86_out;
		end else begin
			bb_9_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_9_predecessor_in_state_1.bb_9_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_111_out) begin 
			bb_9_predecessor_in_state_1_in_data = 32'd8;
		end else if (eq_109_out) begin 
			bb_9_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_9_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_31_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_32_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_1.br_0_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_34_out) begin 
			br_0_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_35_out) begin 
			br_0_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_2.br_10_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_49_out) begin 
			br_10_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_50_out) begin 
			br_10_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_3.br_10_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_58_out) begin 
			br_10_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_59_out) begin 
			br_10_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_1_happened_in_state_4.br_1_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_73_out) begin 
			br_1_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_74_out) begin 
			br_1_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_1_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_1.br_3_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_37_out) begin 
			br_3_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_38_out) begin 
			br_3_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_3.br_4_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_52_out) begin 
			br_4_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_53_out) begin 
			br_4_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_4.br_4_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_76_out) begin 
			br_4_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_77_out) begin 
			br_4_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_5_happened_in_state_4.br_5_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_61_out) begin 
			br_5_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_62_out) begin 
			br_5_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_5_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_6_happened_in_state_4.br_6_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_64_out) begin 
			br_6_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_65_out) begin 
			br_6_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_6_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_7_happened_in_state_4.br_7_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_70_out) begin 
			br_7_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_71_out) begin 
			br_7_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_7_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_8_happened_in_state_1.br_8_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_46_out) begin 
			br_8_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_47_out) begin 
			br_8_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_8_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_9_happened_in_state_1.br_9_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_40_out) begin 
			br_9_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_41_out) begin 
			br_9_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_9_happened_in_state_1_in_data = 0;
		end
	end
	// controller for concat_147.concat_147_in0
	// controller for concat_147.concat_147_in1
	// Insensitive connections
	always @(*) begin
		concat_147_in0 = valid ? data_in_1_9_out_data : data_in_1_9_out_data;
		concat_147_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for concat_148.concat_148_in0
	// controller for concat_148.concat_148_in1
	// Insensitive connections
	always @(*) begin
		concat_148_in0 = valid ? 32'd4 : 32'd4;
		concat_148_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for data_in_0_1.data_in_0_1_in_data
	always @(*) begin
		if (andOp_184_out) begin 
			data_in_0_1_in_data = data_store_0_0;
		end else if (andOp_186_out) begin 
			data_in_0_1_in_data = data_store_1_6;
		end else if (andOp_188_out) begin 
			data_in_0_1_in_data = data_store_2_12;
		end else if (andOp_190_out) begin 
			data_in_0_1_in_data = data_store_3_18;
		end else if (andOp_192_out) begin 
			data_in_0_1_in_data = data_store_4_24;
		end else begin
			data_in_0_1_in_data = 0;
		end
	end
	// controller for data_in_0_3.data_in_0_3_in_data
	always @(*) begin
		if (andOp_184_out) begin 
			data_in_0_3_in_data = data_store_0_2;
		end else if (andOp_186_out) begin 
			data_in_0_3_in_data = data_store_1_8;
		end else if (andOp_188_out) begin 
			data_in_0_3_in_data = data_store_2_14;
		end else if (andOp_190_out) begin 
			data_in_0_3_in_data = data_store_3_20;
		end else if (andOp_192_out) begin 
			data_in_0_3_in_data = data_store_4_26;
		end else begin
			data_in_0_3_in_data = 0;
		end
	end
	// controller for data_in_0_5.data_in_0_5_in_data
	always @(*) begin
		if (andOp_184_out) begin 
			data_in_0_5_in_data = data_store_0_4;
		end else if (andOp_186_out) begin 
			data_in_0_5_in_data = data_store_1_10;
		end else if (andOp_188_out) begin 
			data_in_0_5_in_data = data_store_2_16;
		end else if (andOp_190_out) begin 
			data_in_0_5_in_data = data_store_3_22;
		end else if (andOp_192_out) begin 
			data_in_0_5_in_data = data_store_4_28;
		end else begin
			data_in_0_5_in_data = 0;
		end
	end
	// controller for data_in_1_11.data_in_1_11_in_data
	always @(*) begin
		if (andOp_221_out) begin 
			data_in_1_11_in_data = data_store_0_4;
		end else if (andOp_223_out) begin 
			data_in_1_11_in_data = data_store_1_10;
		end else if (andOp_225_out) begin 
			data_in_1_11_in_data = data_store_2_16;
		end else if (andOp_227_out) begin 
			data_in_1_11_in_data = data_store_3_22;
		end else if (andOp_229_out) begin 
			data_in_1_11_in_data = data_store_4_28;
		end else begin
			data_in_1_11_in_data = 0;
		end
	end
	// controller for data_in_1_7.data_in_1_7_in_data
	always @(*) begin
		if (andOp_221_out) begin 
			data_in_1_7_in_data = data_store_0_0;
		end else if (andOp_223_out) begin 
			data_in_1_7_in_data = data_store_1_6;
		end else if (andOp_225_out) begin 
			data_in_1_7_in_data = data_store_2_12;
		end else if (andOp_227_out) begin 
			data_in_1_7_in_data = data_store_3_18;
		end else if (andOp_229_out) begin 
			data_in_1_7_in_data = data_store_4_24;
		end else begin
			data_in_1_7_in_data = 0;
		end
	end
	// controller for data_in_1_9.data_in_1_9_in_data
	always @(*) begin
		if (andOp_221_out) begin 
			data_in_1_9_in_data = data_store_0_2;
		end else if (andOp_223_out) begin 
			data_in_1_9_in_data = data_store_1_8;
		end else if (andOp_225_out) begin 
			data_in_1_9_in_data = data_store_2_14;
		end else if (andOp_227_out) begin 
			data_in_1_9_in_data = data_store_3_20;
		end else if (andOp_229_out) begin 
			data_in_1_9_in_data = data_store_4_26;
		end else begin
			data_in_1_9_in_data = 0;
		end
	end
	// controller for data_in_2_13.data_in_2_13_in_data
	always @(*) begin
		if (andOp_258_out) begin 
			data_in_2_13_in_data = data_store_0_0;
		end else if (andOp_260_out) begin 
			data_in_2_13_in_data = data_store_1_6;
		end else if (andOp_262_out) begin 
			data_in_2_13_in_data = data_store_2_12;
		end else if (andOp_264_out) begin 
			data_in_2_13_in_data = data_store_3_18;
		end else if (andOp_266_out) begin 
			data_in_2_13_in_data = data_store_4_24;
		end else begin
			data_in_2_13_in_data = 0;
		end
	end
	// controller for data_in_2_15.data_in_2_15_in_data
	always @(*) begin
		if (andOp_258_out) begin 
			data_in_2_15_in_data = data_store_0_2;
		end else if (andOp_260_out) begin 
			data_in_2_15_in_data = data_store_1_8;
		end else if (andOp_262_out) begin 
			data_in_2_15_in_data = data_store_2_14;
		end else if (andOp_264_out) begin 
			data_in_2_15_in_data = data_store_3_20;
		end else if (andOp_266_out) begin 
			data_in_2_15_in_data = data_store_4_26;
		end else begin
			data_in_2_15_in_data = 0;
		end
	end
	// controller for data_in_2_17.data_in_2_17_in_data
	always @(*) begin
		if (andOp_258_out) begin 
			data_in_2_17_in_data = data_store_0_4;
		end else if (andOp_260_out) begin 
			data_in_2_17_in_data = data_store_1_10;
		end else if (andOp_262_out) begin 
			data_in_2_17_in_data = data_store_2_16;
		end else if (andOp_264_out) begin 
			data_in_2_17_in_data = data_store_3_22;
		end else if (andOp_266_out) begin 
			data_in_2_17_in_data = data_store_4_28;
		end else begin
			data_in_2_17_in_data = 0;
		end
	end
	// controller for data_in_3_19.data_in_3_19_in_data
	always @(*) begin
		if (andOp_295_out) begin 
			data_in_3_19_in_data = data_store_0_0;
		end else if (andOp_297_out) begin 
			data_in_3_19_in_data = data_store_1_6;
		end else if (andOp_299_out) begin 
			data_in_3_19_in_data = data_store_2_12;
		end else if (andOp_301_out) begin 
			data_in_3_19_in_data = data_store_3_18;
		end else if (andOp_303_out) begin 
			data_in_3_19_in_data = data_store_4_24;
		end else begin
			data_in_3_19_in_data = 0;
		end
	end
	// controller for data_in_3_21.data_in_3_21_in_data
	always @(*) begin
		if (andOp_295_out) begin 
			data_in_3_21_in_data = data_store_0_2;
		end else if (andOp_297_out) begin 
			data_in_3_21_in_data = data_store_1_8;
		end else if (andOp_299_out) begin 
			data_in_3_21_in_data = data_store_2_14;
		end else if (andOp_301_out) begin 
			data_in_3_21_in_data = data_store_3_20;
		end else if (andOp_303_out) begin 
			data_in_3_21_in_data = data_store_4_26;
		end else begin
			data_in_3_21_in_data = 0;
		end
	end
	// controller for data_in_3_23.data_in_3_23_in_data
	always @(*) begin
		if (andOp_295_out) begin 
			data_in_3_23_in_data = data_store_0_4;
		end else if (andOp_297_out) begin 
			data_in_3_23_in_data = data_store_1_10;
		end else if (andOp_299_out) begin 
			data_in_3_23_in_data = data_store_2_16;
		end else if (andOp_301_out) begin 
			data_in_3_23_in_data = data_store_3_22;
		end else if (andOp_303_out) begin 
			data_in_3_23_in_data = data_store_4_28;
		end else begin
			data_in_3_23_in_data = 0;
		end
	end
	// controller for data_in_4_25.data_in_4_25_in_data
	always @(*) begin
		if (andOp_332_out) begin 
			data_in_4_25_in_data = data_store_0_0;
		end else if (andOp_334_out) begin 
			data_in_4_25_in_data = data_store_1_6;
		end else if (andOp_336_out) begin 
			data_in_4_25_in_data = data_store_2_12;
		end else if (andOp_338_out) begin 
			data_in_4_25_in_data = data_store_3_18;
		end else if (andOp_340_out) begin 
			data_in_4_25_in_data = data_store_4_24;
		end else begin
			data_in_4_25_in_data = 0;
		end
	end
	// controller for data_in_4_27.data_in_4_27_in_data
	always @(*) begin
		if (andOp_332_out) begin 
			data_in_4_27_in_data = data_store_0_2;
		end else if (andOp_334_out) begin 
			data_in_4_27_in_data = data_store_1_8;
		end else if (andOp_336_out) begin 
			data_in_4_27_in_data = data_store_2_14;
		end else if (andOp_338_out) begin 
			data_in_4_27_in_data = data_store_3_20;
		end else if (andOp_340_out) begin 
			data_in_4_27_in_data = data_store_4_26;
		end else begin
			data_in_4_27_in_data = 0;
		end
	end
	// controller for data_in_4_29.data_in_4_29_in_data
	always @(*) begin
		if (andOp_332_out) begin 
			data_in_4_29_in_data = data_store_0_4;
		end else if (andOp_334_out) begin 
			data_in_4_29_in_data = data_store_1_10;
		end else if (andOp_336_out) begin 
			data_in_4_29_in_data = data_store_2_16;
		end else if (andOp_338_out) begin 
			data_in_4_29_in_data = data_store_3_22;
		end else if (andOp_340_out) begin 
			data_in_4_29_in_data = data_store_4_28;
		end else begin
			data_in_4_29_in_data = 0;
		end
	end
	// controller for eq_101.eq_101_in0
	// controller for eq_101.eq_101_in1
	// Insensitive connections
	always @(*) begin
		eq_101_in0 = valid ? 32'd1 : 32'd1;
		eq_101_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_103.eq_103_in0
	// controller for eq_103.eq_103_in1
	// Insensitive connections
	always @(*) begin
		eq_103_in0 = valid ? 32'd4 : 32'd4;
		eq_103_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_104.eq_104_in0
	// controller for eq_104.eq_104_in1
	// Insensitive connections
	always @(*) begin
		eq_104_in0 = valid ? 32'd0 : 32'd0;
		eq_104_in1 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
	end
	// controller for eq_105.eq_105_in0
	// controller for eq_105.eq_105_in1
	// Insensitive connections
	always @(*) begin
		eq_105_in0 = valid ? 32'd0 : 32'd0;
		eq_105_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_106.eq_106_in0
	// controller for eq_106.eq_106_in1
	// Insensitive connections
	always @(*) begin
		eq_106_in0 = valid ? 32'd3 : 32'd3;
		eq_106_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_109.eq_109_in0
	// controller for eq_109.eq_109_in1
	// Insensitive connections
	always @(*) begin
		eq_109_in0 = valid ? 32'd9 : 32'd9;
		eq_109_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_112.eq_112_in0
	// controller for eq_112.eq_112_in1
	// Insensitive connections
	always @(*) begin
		eq_112_in0 = valid ? 32'd8 : 32'd8;
		eq_112_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_115.eq_115_in0
	// controller for eq_115.eq_115_in1
	// Insensitive connections
	always @(*) begin
		eq_115_in0 = valid ? 32'd10 : 32'd10;
		eq_115_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_116.eq_116_in0
	// controller for eq_116.eq_116_in1
	// Insensitive connections
	always @(*) begin
		eq_116_in0 = valid ? 32'd4 : 32'd4;
		eq_116_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_119.eq_119_in0
	// controller for eq_119.eq_119_in1
	// Insensitive connections
	always @(*) begin
		eq_119_in0 = valid ? 32'd10 : 32'd10;
		eq_119_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_120.eq_120_in0
	// controller for eq_120.eq_120_in1
	// Insensitive connections
	always @(*) begin
		eq_120_in0 = valid ? 32'd5 : 32'd5;
		eq_120_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_123.eq_123_in0
	// controller for eq_123.eq_123_in1
	// Insensitive connections
	always @(*) begin
		eq_123_in0 = valid ? 32'd6 : 32'd6;
		eq_123_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_126.eq_126_in0
	// controller for eq_126.eq_126_in1
	// Insensitive connections
	always @(*) begin
		eq_126_in0 = valid ? 32'd7 : 32'd7;
		eq_126_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_129.eq_129_in0
	// controller for eq_129.eq_129_in1
	// Insensitive connections
	always @(*) begin
		eq_129_in0 = valid ? 32'd2 : 32'd2;
		eq_129_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_132.eq_132_in0
	// controller for eq_132.eq_132_in1
	// Insensitive connections
	always @(*) begin
		eq_132_in0 = valid ? 32'd1 : 32'd1;
		eq_132_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_135.eq_135_in0
	// controller for eq_135.eq_135_in1
	// Insensitive connections
	always @(*) begin
		eq_135_in0 = valid ? 32'd4 : 32'd4;
		eq_135_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_151.eq_151_in0
	// controller for eq_151.eq_151_in1
	// Insensitive connections
	always @(*) begin
		eq_151_in0 = valid ? 32'd10 : 32'd10;
		eq_151_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_183.eq_183_in0
	// controller for eq_183.eq_183_in1
	// Insensitive connections
	always @(*) begin
		eq_183_in0 = valid ? 32'd0 : 32'd0;
		eq_183_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_185.eq_185_in0
	// controller for eq_185.eq_185_in1
	// Insensitive connections
	always @(*) begin
		eq_185_in0 = valid ? 32'd1 : 32'd1;
		eq_185_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_187.eq_187_in0
	// controller for eq_187.eq_187_in1
	// Insensitive connections
	always @(*) begin
		eq_187_in0 = valid ? 32'd2 : 32'd2;
		eq_187_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_189.eq_189_in0
	// controller for eq_189.eq_189_in1
	// Insensitive connections
	always @(*) begin
		eq_189_in0 = valid ? 32'd3 : 32'd3;
		eq_189_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_191.eq_191_in0
	// controller for eq_191.eq_191_in1
	// Insensitive connections
	always @(*) begin
		eq_191_in0 = valid ? 32'd4 : 32'd4;
		eq_191_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_194.eq_194_in0
	// controller for eq_194.eq_194_in1
	// Insensitive connections
	always @(*) begin
		eq_194_in0 = valid ? 32'd1 : 32'd1;
		eq_194_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_203.eq_203_in0
	// controller for eq_203.eq_203_in1
	// Insensitive connections
	always @(*) begin
		eq_203_in0 = valid ? 32'd3 : 32'd3;
		eq_203_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_212.eq_212_in0
	// controller for eq_212.eq_212_in1
	// Insensitive connections
	always @(*) begin
		eq_212_in0 = valid ? 32'd3 : 32'd3;
		eq_212_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_220.eq_220_in0
	// controller for eq_220.eq_220_in1
	// Insensitive connections
	always @(*) begin
		eq_220_in0 = valid ? 32'd0 : 32'd0;
		eq_220_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_222.eq_222_in0
	// controller for eq_222.eq_222_in1
	// Insensitive connections
	always @(*) begin
		eq_222_in0 = valid ? 32'd1 : 32'd1;
		eq_222_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_224.eq_224_in0
	// controller for eq_224.eq_224_in1
	// Insensitive connections
	always @(*) begin
		eq_224_in0 = valid ? 32'd2 : 32'd2;
		eq_224_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_226.eq_226_in0
	// controller for eq_226.eq_226_in1
	// Insensitive connections
	always @(*) begin
		eq_226_in0 = valid ? 32'd3 : 32'd3;
		eq_226_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_228.eq_228_in0
	// controller for eq_228.eq_228_in1
	// Insensitive connections
	always @(*) begin
		eq_228_in0 = valid ? 32'd4 : 32'd4;
		eq_228_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_231.eq_231_in0
	// controller for eq_231.eq_231_in1
	// Insensitive connections
	always @(*) begin
		eq_231_in0 = valid ? 32'd1 : 32'd1;
		eq_231_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_240.eq_240_in0
	// controller for eq_240.eq_240_in1
	// Insensitive connections
	always @(*) begin
		eq_240_in0 = valid ? 32'd3 : 32'd3;
		eq_240_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_249.eq_249_in0
	// controller for eq_249.eq_249_in1
	// Insensitive connections
	always @(*) begin
		eq_249_in0 = valid ? 32'd3 : 32'd3;
		eq_249_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_257.eq_257_in0
	// controller for eq_257.eq_257_in1
	// Insensitive connections
	always @(*) begin
		eq_257_in0 = valid ? 32'd0 : 32'd0;
		eq_257_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_259.eq_259_in0
	// controller for eq_259.eq_259_in1
	// Insensitive connections
	always @(*) begin
		eq_259_in0 = valid ? 32'd1 : 32'd1;
		eq_259_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_261.eq_261_in0
	// controller for eq_261.eq_261_in1
	// Insensitive connections
	always @(*) begin
		eq_261_in0 = valid ? 32'd2 : 32'd2;
		eq_261_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_263.eq_263_in0
	// controller for eq_263.eq_263_in1
	// Insensitive connections
	always @(*) begin
		eq_263_in0 = valid ? 32'd3 : 32'd3;
		eq_263_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_265.eq_265_in0
	// controller for eq_265.eq_265_in1
	// Insensitive connections
	always @(*) begin
		eq_265_in0 = valid ? 32'd4 : 32'd4;
		eq_265_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_268.eq_268_in0
	// controller for eq_268.eq_268_in1
	// Insensitive connections
	always @(*) begin
		eq_268_in0 = valid ? 32'd1 : 32'd1;
		eq_268_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_277.eq_277_in0
	// controller for eq_277.eq_277_in1
	// Insensitive connections
	always @(*) begin
		eq_277_in0 = valid ? 32'd3 : 32'd3;
		eq_277_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_286.eq_286_in0
	// controller for eq_286.eq_286_in1
	// Insensitive connections
	always @(*) begin
		eq_286_in0 = valid ? 32'd3 : 32'd3;
		eq_286_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_294.eq_294_in0
	// controller for eq_294.eq_294_in1
	// Insensitive connections
	always @(*) begin
		eq_294_in0 = valid ? 32'd0 : 32'd0;
		eq_294_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_296.eq_296_in0
	// controller for eq_296.eq_296_in1
	// Insensitive connections
	always @(*) begin
		eq_296_in0 = valid ? 32'd1 : 32'd1;
		eq_296_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_298.eq_298_in0
	// controller for eq_298.eq_298_in1
	// Insensitive connections
	always @(*) begin
		eq_298_in0 = valid ? 32'd2 : 32'd2;
		eq_298_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_300.eq_300_in0
	// controller for eq_300.eq_300_in1
	// Insensitive connections
	always @(*) begin
		eq_300_in0 = valid ? 32'd3 : 32'd3;
		eq_300_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_302.eq_302_in0
	// controller for eq_302.eq_302_in1
	// Insensitive connections
	always @(*) begin
		eq_302_in0 = valid ? 32'd4 : 32'd4;
		eq_302_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_305.eq_305_in0
	// controller for eq_305.eq_305_in1
	// Insensitive connections
	always @(*) begin
		eq_305_in0 = valid ? 32'd1 : 32'd1;
		eq_305_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_314.eq_314_in0
	// controller for eq_314.eq_314_in1
	// Insensitive connections
	always @(*) begin
		eq_314_in0 = valid ? 32'd3 : 32'd3;
		eq_314_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_323.eq_323_in0
	// controller for eq_323.eq_323_in1
	// Insensitive connections
	always @(*) begin
		eq_323_in0 = valid ? 32'd3 : 32'd3;
		eq_323_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_331.eq_331_in0
	// controller for eq_331.eq_331_in1
	// Insensitive connections
	always @(*) begin
		eq_331_in0 = valid ? 32'd0 : 32'd0;
		eq_331_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_333.eq_333_in0
	// controller for eq_333.eq_333_in1
	// Insensitive connections
	always @(*) begin
		eq_333_in0 = valid ? 32'd1 : 32'd1;
		eq_333_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_335.eq_335_in0
	// controller for eq_335.eq_335_in1
	// Insensitive connections
	always @(*) begin
		eq_335_in0 = valid ? 32'd2 : 32'd2;
		eq_335_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_337.eq_337_in0
	// controller for eq_337.eq_337_in1
	// Insensitive connections
	always @(*) begin
		eq_337_in0 = valid ? 32'd3 : 32'd3;
		eq_337_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_339.eq_339_in0
	// controller for eq_339.eq_339_in1
	// Insensitive connections
	always @(*) begin
		eq_339_in0 = valid ? 32'd4 : 32'd4;
		eq_339_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_342.eq_342_in0
	// controller for eq_342.eq_342_in1
	// Insensitive connections
	always @(*) begin
		eq_342_in0 = valid ? 32'd1 : 32'd1;
		eq_342_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_351.eq_351_in0
	// controller for eq_351.eq_351_in1
	// Insensitive connections
	always @(*) begin
		eq_351_in0 = valid ? 32'd3 : 32'd3;
		eq_351_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_360.eq_360_in0
	// controller for eq_360.eq_360_in1
	// Insensitive connections
	always @(*) begin
		eq_360_in0 = valid ? 32'd3 : 32'd3;
		eq_360_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_81.eq_81_in0
	// controller for eq_81.eq_81_in1
	// Insensitive connections
	always @(*) begin
		eq_81_in0 = valid ? 32'd0 : 32'd0;
		eq_81_in1 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
	end
	// controller for eq_82.eq_82_in0
	// controller for eq_82.eq_82_in1
	// Insensitive connections
	always @(*) begin
		eq_82_in0 = valid ? 32'd0 : 32'd0;
		eq_82_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_83.eq_83_in0
	// controller for eq_83.eq_83_in1
	// Insensitive connections
	always @(*) begin
		eq_83_in0 = valid ? 32'd3 : 32'd3;
		eq_83_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_85.eq_85_in0
	// controller for eq_85.eq_85_in1
	// Insensitive connections
	always @(*) begin
		eq_85_in0 = valid ? 32'd9 : 32'd9;
		eq_85_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_87.eq_87_in0
	// controller for eq_87.eq_87_in1
	// Insensitive connections
	always @(*) begin
		eq_87_in0 = valid ? 32'd8 : 32'd8;
		eq_87_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_89.eq_89_in0
	// controller for eq_89.eq_89_in1
	// Insensitive connections
	always @(*) begin
		eq_89_in0 = valid ? 32'd10 : 32'd10;
		eq_89_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_90.eq_90_in0
	// controller for eq_90.eq_90_in1
	// Insensitive connections
	always @(*) begin
		eq_90_in0 = valid ? 32'd4 : 32'd4;
		eq_90_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_92.eq_92_in0
	// controller for eq_92.eq_92_in1
	// Insensitive connections
	always @(*) begin
		eq_92_in0 = valid ? 32'd10 : 32'd10;
		eq_92_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_93.eq_93_in0
	// controller for eq_93.eq_93_in1
	// Insensitive connections
	always @(*) begin
		eq_93_in0 = valid ? 32'd5 : 32'd5;
		eq_93_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_95.eq_95_in0
	// controller for eq_95.eq_95_in1
	// Insensitive connections
	always @(*) begin
		eq_95_in0 = valid ? 32'd6 : 32'd6;
		eq_95_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_97.eq_97_in0
	// controller for eq_97.eq_97_in1
	// Insensitive connections
	always @(*) begin
		eq_97_in0 = valid ? 32'd7 : 32'd7;
		eq_97_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_99.eq_99_in0
	// controller for eq_99.eq_99_in1
	// Insensitive connections
	always @(*) begin
		eq_99_in0 = valid ? 32'd2 : 32'd2;
		eq_99_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for icmp_17.cmp_in0_icmp_17
	// controller for icmp_17.cmp_in1_icmp_17
	// Insensitive connections
	always @(*) begin
		cmp_in0_icmp_17 = valid ? add_out_add_16 : add_out_add_16;
		cmp_in1_icmp_17 = valid ? 32'd4 : 32'd4;
	end
	// controller for in.in_read_valid_reg
	always @(*) begin
		if (andOp_144_out) begin 
			in_read_valid_reg = -(1'd1);
		end else begin
			in_read_valid_reg = 0;
		end
	end
	// controller for notOp_107.notOp_107_in0
	// Insensitive connections
	always @(*) begin
		notOp_107_in0 = valid ? eq_106_out : eq_106_out;
	end
	// controller for notOp_110.notOp_110_in0
	// Insensitive connections
	always @(*) begin
		notOp_110_in0 = valid ? eq_109_out : eq_109_out;
	end
	// controller for notOp_113.notOp_113_in0
	// Insensitive connections
	always @(*) begin
		notOp_113_in0 = valid ? eq_112_out : eq_112_out;
	end
	// controller for notOp_117.notOp_117_in0
	// Insensitive connections
	always @(*) begin
		notOp_117_in0 = valid ? eq_116_out : eq_116_out;
	end
	// controller for notOp_121.notOp_121_in0
	// Insensitive connections
	always @(*) begin
		notOp_121_in0 = valid ? eq_120_out : eq_120_out;
	end
	// controller for notOp_124.notOp_124_in0
	// Insensitive connections
	always @(*) begin
		notOp_124_in0 = valid ? eq_123_out : eq_123_out;
	end
	// controller for notOp_127.notOp_127_in0
	// Insensitive connections
	always @(*) begin
		notOp_127_in0 = valid ? eq_126_out : eq_126_out;
	end
	// controller for notOp_130.notOp_130_in0
	// Insensitive connections
	always @(*) begin
		notOp_130_in0 = valid ? eq_129_out : eq_129_out;
	end
	// controller for notOp_133.notOp_133_in0
	// Insensitive connections
	always @(*) begin
		notOp_133_in0 = valid ? eq_132_out : eq_132_out;
	end
	// controller for notOp_163.notOp_163_in0
	// Insensitive connections
	always @(*) begin
		notOp_163_in0 = valid ? andOp_159_out : andOp_159_out;
	end
	// controller for notOp_165.notOp_165_in0
	// Insensitive connections
	always @(*) begin
		notOp_165_in0 = valid ? andOp_44_out : andOp_44_out;
	end
	// controller for notOp_167.notOp_167_in0
	// Insensitive connections
	always @(*) begin
		notOp_167_in0 = valid ? andOp_56_out : andOp_56_out;
	end
	// controller for notOp_169.notOp_169_in0
	// Insensitive connections
	always @(*) begin
		notOp_169_in0 = valid ? andOp_42_out : andOp_42_out;
	end
	// controller for notOp_171.notOp_171_in0
	// Insensitive connections
	always @(*) begin
		notOp_171_in0 = valid ? andOp_160_out : andOp_160_out;
	end
	// controller for notOp_173.notOp_173_in0
	// Insensitive connections
	always @(*) begin
		notOp_173_in0 = valid ? andOp_161_out : andOp_161_out;
	end
	// controller for notOp_175.notOp_175_in0
	// Insensitive connections
	always @(*) begin
		notOp_175_in0 = valid ? andOp_162_out : andOp_162_out;
	end
	// controller for notOp_177.notOp_177_in0
	// Insensitive connections
	always @(*) begin
		notOp_177_in0 = valid ? andOp_68_out : andOp_68_out;
	end
	// controller for notOp_196.notOp_196_in0
	// Insensitive connections
	always @(*) begin
		notOp_196_in0 = valid ? eq_194_out : eq_194_out;
	end
	// controller for notOp_198.notOp_198_in0
	// Insensitive connections
	always @(*) begin
		notOp_198_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_200.notOp_200_in0
	// Insensitive connections
	always @(*) begin
		notOp_200_in0 = valid ? andOp_195_out : andOp_195_out;
	end
	// controller for notOp_205.notOp_205_in0
	// Insensitive connections
	always @(*) begin
		notOp_205_in0 = valid ? eq_203_out : eq_203_out;
	end
	// controller for notOp_207.notOp_207_in0
	// Insensitive connections
	always @(*) begin
		notOp_207_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_209.notOp_209_in0
	// Insensitive connections
	always @(*) begin
		notOp_209_in0 = valid ? andOp_204_out : andOp_204_out;
	end
	// controller for notOp_214.notOp_214_in0
	// Insensitive connections
	always @(*) begin
		notOp_214_in0 = valid ? eq_212_out : eq_212_out;
	end
	// controller for notOp_216.notOp_216_in0
	// Insensitive connections
	always @(*) begin
		notOp_216_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_218.notOp_218_in0
	// Insensitive connections
	always @(*) begin
		notOp_218_in0 = valid ? andOp_213_out : andOp_213_out;
	end
	// controller for notOp_233.notOp_233_in0
	// Insensitive connections
	always @(*) begin
		notOp_233_in0 = valid ? eq_231_out : eq_231_out;
	end
	// controller for notOp_235.notOp_235_in0
	// Insensitive connections
	always @(*) begin
		notOp_235_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
	end
	// controller for notOp_237.notOp_237_in0
	// Insensitive connections
	always @(*) begin
		notOp_237_in0 = valid ? andOp_232_out : andOp_232_out;
	end
	// controller for notOp_242.notOp_242_in0
	// Insensitive connections
	always @(*) begin
		notOp_242_in0 = valid ? eq_240_out : eq_240_out;
	end
	// controller for notOp_244.notOp_244_in0
	// Insensitive connections
	always @(*) begin
		notOp_244_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_246.notOp_246_in0
	// Insensitive connections
	always @(*) begin
		notOp_246_in0 = valid ? andOp_241_out : andOp_241_out;
	end
	// controller for notOp_251.notOp_251_in0
	// Insensitive connections
	always @(*) begin
		notOp_251_in0 = valid ? eq_249_out : eq_249_out;
	end
	// controller for notOp_253.notOp_253_in0
	// Insensitive connections
	always @(*) begin
		notOp_253_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_255.notOp_255_in0
	// Insensitive connections
	always @(*) begin
		notOp_255_in0 = valid ? andOp_250_out : andOp_250_out;
	end
	// controller for notOp_270.notOp_270_in0
	// Insensitive connections
	always @(*) begin
		notOp_270_in0 = valid ? eq_268_out : eq_268_out;
	end
	// controller for notOp_272.notOp_272_in0
	// Insensitive connections
	always @(*) begin
		notOp_272_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_274.notOp_274_in0
	// Insensitive connections
	always @(*) begin
		notOp_274_in0 = valid ? andOp_269_out : andOp_269_out;
	end
	// controller for notOp_279.notOp_279_in0
	// Insensitive connections
	always @(*) begin
		notOp_279_in0 = valid ? eq_277_out : eq_277_out;
	end
	// controller for notOp_281.notOp_281_in0
	// Insensitive connections
	always @(*) begin
		notOp_281_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_283.notOp_283_in0
	// Insensitive connections
	always @(*) begin
		notOp_283_in0 = valid ? andOp_278_out : andOp_278_out;
	end
	// controller for notOp_288.notOp_288_in0
	// Insensitive connections
	always @(*) begin
		notOp_288_in0 = valid ? eq_286_out : eq_286_out;
	end
	// controller for notOp_290.notOp_290_in0
	// Insensitive connections
	always @(*) begin
		notOp_290_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_292.notOp_292_in0
	// Insensitive connections
	always @(*) begin
		notOp_292_in0 = valid ? andOp_287_out : andOp_287_out;
	end
	// controller for notOp_307.notOp_307_in0
	// Insensitive connections
	always @(*) begin
		notOp_307_in0 = valid ? eq_305_out : eq_305_out;
	end
	// controller for notOp_309.notOp_309_in0
	// Insensitive connections
	always @(*) begin
		notOp_309_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_311.notOp_311_in0
	// Insensitive connections
	always @(*) begin
		notOp_311_in0 = valid ? andOp_306_out : andOp_306_out;
	end
	// controller for notOp_316.notOp_316_in0
	// Insensitive connections
	always @(*) begin
		notOp_316_in0 = valid ? eq_314_out : eq_314_out;
	end
	// controller for notOp_318.notOp_318_in0
	// Insensitive connections
	always @(*) begin
		notOp_318_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
	end
	// controller for notOp_32.notOp_32_in0
	// Insensitive connections
	always @(*) begin
		notOp_32_in0 = valid ? andOp_31_out : andOp_31_out;
	end
	// controller for notOp_320.notOp_320_in0
	// Insensitive connections
	always @(*) begin
		notOp_320_in0 = valid ? andOp_315_out : andOp_315_out;
	end
	// controller for notOp_325.notOp_325_in0
	// Insensitive connections
	always @(*) begin
		notOp_325_in0 = valid ? eq_323_out : eq_323_out;
	end
	// controller for notOp_327.notOp_327_in0
	// Insensitive connections
	always @(*) begin
		notOp_327_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
	end
	// controller for notOp_329.notOp_329_in0
	// Insensitive connections
	always @(*) begin
		notOp_329_in0 = valid ? andOp_324_out : andOp_324_out;
	end
	// controller for notOp_344.notOp_344_in0
	// Insensitive connections
	always @(*) begin
		notOp_344_in0 = valid ? eq_342_out : eq_342_out;
	end
	// controller for notOp_346.notOp_346_in0
	// Insensitive connections
	always @(*) begin
		notOp_346_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_348.notOp_348_in0
	// Insensitive connections
	always @(*) begin
		notOp_348_in0 = valid ? andOp_343_out : andOp_343_out;
	end
	// controller for notOp_35.notOp_35_in0
	// Insensitive connections
	always @(*) begin
		notOp_35_in0 = valid ? andOp_34_out : andOp_34_out;
	end
	// controller for notOp_353.notOp_353_in0
	// Insensitive connections
	always @(*) begin
		notOp_353_in0 = valid ? eq_351_out : eq_351_out;
	end
	// controller for notOp_355.notOp_355_in0
	// Insensitive connections
	always @(*) begin
		notOp_355_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
	end
	// controller for notOp_357.notOp_357_in0
	// Insensitive connections
	always @(*) begin
		notOp_357_in0 = valid ? andOp_352_out : andOp_352_out;
	end
	// controller for notOp_362.notOp_362_in0
	// Insensitive connections
	always @(*) begin
		notOp_362_in0 = valid ? eq_360_out : eq_360_out;
	end
	// controller for notOp_364.notOp_364_in0
	// Insensitive connections
	always @(*) begin
		notOp_364_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
	end
	// controller for notOp_366.notOp_366_in0
	// Insensitive connections
	always @(*) begin
		notOp_366_in0 = valid ? andOp_361_out : andOp_361_out;
	end
	// controller for notOp_38.notOp_38_in0
	// Insensitive connections
	always @(*) begin
		notOp_38_in0 = valid ? andOp_37_out : andOp_37_out;
	end
	// controller for notOp_41.notOp_41_in0
	// Insensitive connections
	always @(*) begin
		notOp_41_in0 = valid ? andOp_40_out : andOp_40_out;
	end
	// controller for notOp_43.notOp_43_in0
	// Insensitive connections
	always @(*) begin
		notOp_43_in0 = valid ? in_read_ready : in_read_ready;
	end
	// controller for notOp_47.notOp_47_in0
	// Insensitive connections
	always @(*) begin
		notOp_47_in0 = valid ? andOp_46_out : andOp_46_out;
	end
	// controller for notOp_50.notOp_50_in0
	// Insensitive connections
	always @(*) begin
		notOp_50_in0 = valid ? andOp_49_out : andOp_49_out;
	end
	// controller for notOp_53.notOp_53_in0
	// Insensitive connections
	always @(*) begin
		notOp_53_in0 = valid ? andOp_52_out : andOp_52_out;
	end
	// controller for notOp_55.notOp_55_in0
	// Insensitive connections
	always @(*) begin
		notOp_55_in0 = valid ? data_in_4_29_out_data : data_in_4_29_out_data;
	end
	// controller for notOp_59.notOp_59_in0
	// Insensitive connections
	always @(*) begin
		notOp_59_in0 = valid ? andOp_58_out : andOp_58_out;
	end
	// controller for notOp_62.notOp_62_in0
	// Insensitive connections
	always @(*) begin
		notOp_62_in0 = valid ? andOp_61_out : andOp_61_out;
	end
	// controller for notOp_65.notOp_65_in0
	// Insensitive connections
	always @(*) begin
		notOp_65_in0 = valid ? andOp_64_out : andOp_64_out;
	end
	// controller for notOp_67.notOp_67_in0
	// Insensitive connections
	always @(*) begin
		notOp_67_in0 = valid ? out_write_ready : out_write_ready;
	end
	// controller for notOp_71.notOp_71_in0
	// Insensitive connections
	always @(*) begin
		notOp_71_in0 = valid ? andOp_70_out : andOp_70_out;
	end
	// controller for notOp_74.notOp_74_in0
	// Insensitive connections
	always @(*) begin
		notOp_74_in0 = valid ? andOp_73_out : andOp_73_out;
	end
	// controller for notOp_77.notOp_77_in0
	// Insensitive connections
	always @(*) begin
		notOp_77_in0 = valid ? andOp_76_out : andOp_76_out;
	end
	// controller for notOp_79.notOp_79_in0
	// Insensitive connections
	always @(*) begin
		notOp_79_in0 = valid ? data_in_4_29_out_data : data_in_4_29_out_data;
	end
	// controller for orOp_100.orOp_100_in0
	// controller for orOp_100.orOp_100_in1
	// Insensitive connections
	always @(*) begin
		orOp_100_in0 = valid ? eq_99_out : eq_99_out;
		orOp_100_in1 = valid ? andOp_70_out : andOp_70_out;
	end
	// controller for orOp_102.orOp_102_in0
	// controller for orOp_102.orOp_102_in1
	// Insensitive connections
	always @(*) begin
		orOp_102_in0 = valid ? eq_101_out : eq_101_out;
		orOp_102_in1 = valid ? andOp_54_out : andOp_54_out;
	end
	// controller for orOp_84.orOp_84_in0
	// controller for orOp_84.orOp_84_in1
	// Insensitive connections
	always @(*) begin
		orOp_84_in0 = valid ? eq_83_out : eq_83_out;
		orOp_84_in1 = valid ? andOp_31_out : andOp_31_out;
	end
	// controller for orOp_86.orOp_86_in0
	// controller for orOp_86.orOp_86_in1
	// Insensitive connections
	always @(*) begin
		orOp_86_in0 = valid ? eq_85_out : eq_85_out;
		orOp_86_in1 = valid ? andOp_46_out : andOp_46_out;
	end
	// controller for orOp_88.orOp_88_in0
	// controller for orOp_88.orOp_88_in1
	// Insensitive connections
	always @(*) begin
		orOp_88_in0 = valid ? eq_87_out : eq_87_out;
		orOp_88_in1 = valid ? andOp_37_out : andOp_37_out;
	end
	// controller for orOp_91.orOp_91_in0
	// controller for orOp_91.orOp_91_in1
	// Insensitive connections
	always @(*) begin
		orOp_91_in0 = valid ? eq_90_out : eq_90_out;
		orOp_91_in1 = valid ? andOp_49_out : andOp_49_out;
	end
	// controller for orOp_94.orOp_94_in0
	// controller for orOp_94.orOp_94_in1
	// Insensitive connections
	always @(*) begin
		orOp_94_in0 = valid ? eq_93_out : eq_93_out;
		orOp_94_in1 = valid ? andOp_73_out : andOp_73_out;
	end
	// controller for orOp_96.orOp_96_in0
	// controller for orOp_96.orOp_96_in1
	// Insensitive connections
	always @(*) begin
		orOp_96_in0 = valid ? eq_95_out : eq_95_out;
		orOp_96_in1 = valid ? andOp_61_out : andOp_61_out;
	end
	// controller for orOp_98.orOp_98_in0
	// controller for orOp_98.orOp_98_in1
	// Insensitive connections
	always @(*) begin
		orOp_98_in0 = valid ? eq_97_out : eq_97_out;
		orOp_98_in1 = valid ? andOp_66_out : andOp_66_out;
	end
	// controller for out.out_in_data_reg
	always @(*) begin
		if (andOp_155_out) begin 
			out_in_data_reg = rdata_ram_0;
		end else begin
			out_in_data_reg = 0;
		end
	end
	// controller for out.out_write_valid_reg
	always @(*) begin
		if (andOp_154_out) begin 
			out_write_valid_reg = -(1'd1);
		end else begin
			out_write_valid_reg = 0;
		end
	end
	// controller for phi_8.phi_in_phi_8
	// controller for phi_8.phi_last_block_phi_8
	// controller for phi_8.phi_s_phi_8
	// Insensitive connections
	always @(*) begin
		phi_in_phi_8 = valid ? concat_147_out : concat_147_out;
		phi_last_block_phi_8 = valid ? bb_3_predecessor_in_state_1_out_data : bb_3_predecessor_in_state_1_out_data;
		phi_s_phi_8 = valid ? concat_148_out : concat_148_out;
	end
	// controller for ram_0.raddr_ram_0_reg
	always @(*) begin
		if (andOp_140_out) begin 
			raddr_ram_0_reg = 32'd0;
		end else if (andOp_142_out) begin 
			raddr_ram_0_reg = 32'd0;
		end else begin
			raddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.waddr_ram_0_reg
	always @(*) begin
		if (andOp_139_out) begin 
			waddr_ram_0_reg = 32'd0;
		end else if (andOp_141_out) begin 
			waddr_ram_0_reg = 32'd0;
		end else begin
			waddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wdata_ram_0_reg
	always @(*) begin
		if (andOp_139_out) begin 
			wdata_ram_0_reg = 32'd0;
		end else if (andOp_141_out) begin 
			wdata_ram_0_reg = add_out_add_14;
		end else begin
			wdata_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wen_ram_0_reg
	always @(*) begin
		if (andOp_139_out) begin 
			wen_ram_0_reg = 1'd1;
		end else if (andOp_141_out) begin 
			wen_ram_0_reg = 1'd1;
		end else begin
			wen_ram_0_reg = 0;
		end
	end
	// controller for ret_21.valid_reg
	always @(*) begin
		if (andOp_158_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// controller for tmp_output_150.tmp_output_150_in_data
	always @(*) begin
		if (eq_151_out) begin 
			tmp_output_150_in_data = in_out_data;
		end else begin
			tmp_output_150_in_data = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			add_tmp_5 <= 0;
		end else begin
			if (andOp_181_out) begin
				add_tmp_5 <= add_out_add_16;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			call_tmp_2 <= 0;
		end else begin
			if (andOp_180_out) begin
				call_tmp_2 <= in_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_0 <= 0;
		end else begin
			if (andOp_195_out) begin
				data_store_0_0 <= phi_out_phi_8;
			end
			if (andOp_201_out) begin
				data_store_0_0 <= data_in_0_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_2 <= 0;
		end else begin
			if (andOp_204_out) begin
				data_store_0_2 <= add_out_add_16;
			end
			if (andOp_210_out) begin
				data_store_0_2 <= data_in_0_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_4 <= 0;
		end else begin
			if (andOp_213_out) begin
				data_store_0_4 <= cmp_out_icmp_17;
			end
			if (andOp_219_out) begin
				data_store_0_4 <= data_in_0_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_10 <= 0;
		end else begin
			if (andOp_250_out) begin
				data_store_1_10 <= cmp_out_icmp_17;
			end
			if (andOp_256_out) begin
				data_store_1_10 <= data_in_1_11_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_6 <= 0;
		end else begin
			if (andOp_232_out) begin
				data_store_1_6 <= phi_out_phi_8;
			end
			if (andOp_238_out) begin
				data_store_1_6 <= data_in_1_7_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_8 <= 0;
		end else begin
			if (andOp_241_out) begin
				data_store_1_8 <= add_out_add_16;
			end
			if (andOp_247_out) begin
				data_store_1_8 <= data_in_1_9_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_12 <= 0;
		end else begin
			if (andOp_269_out) begin
				data_store_2_12 <= phi_out_phi_8;
			end
			if (andOp_275_out) begin
				data_store_2_12 <= data_in_2_13_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_14 <= 0;
		end else begin
			if (andOp_278_out) begin
				data_store_2_14 <= add_out_add_16;
			end
			if (andOp_284_out) begin
				data_store_2_14 <= data_in_2_15_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_16 <= 0;
		end else begin
			if (andOp_287_out) begin
				data_store_2_16 <= cmp_out_icmp_17;
			end
			if (andOp_293_out) begin
				data_store_2_16 <= data_in_2_17_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_18 <= 0;
		end else begin
			if (andOp_306_out) begin
				data_store_3_18 <= phi_out_phi_8;
			end
			if (andOp_312_out) begin
				data_store_3_18 <= data_in_3_19_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_20 <= 0;
		end else begin
			if (andOp_315_out) begin
				data_store_3_20 <= add_out_add_16;
			end
			if (andOp_321_out) begin
				data_store_3_20 <= data_in_3_21_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_22 <= 0;
		end else begin
			if (andOp_324_out) begin
				data_store_3_22 <= cmp_out_icmp_17;
			end
			if (andOp_330_out) begin
				data_store_3_22 <= data_in_3_23_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_24 <= 0;
		end else begin
			if (andOp_343_out) begin
				data_store_4_24 <= phi_out_phi_8;
			end
			if (andOp_349_out) begin
				data_store_4_24 <= data_in_4_25_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_26 <= 0;
		end else begin
			if (andOp_352_out) begin
				data_store_4_26 <= add_out_add_16;
			end
			if (andOp_358_out) begin
				data_store_4_26 <= data_in_4_27_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_28 <= 0;
		end else begin
			if (andOp_361_out) begin
				data_store_4_28 <= cmp_out_icmp_17;
			end
			if (andOp_367_out) begin
				data_store_4_28 <= data_in_4_29_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_159_out) begin
				global_state <= 32'd1;
			end
			if (andOp_160_out) begin
				global_state <= 32'd3;
			end
			if (andOp_161_out) begin
				global_state <= 32'd4;
			end
			if (andOp_162_out) begin
				global_state <= 32'd4;
			end
			if (andOp_42_out) begin
				global_state <= 32'd2;
			end
			if (andOp_44_out) begin
				global_state <= 32'd1;
			end
			if (andOp_56_out) begin
				global_state <= 32'd1;
			end
			if (andOp_68_out) begin
				global_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			icmp_tmp_6 <= 0;
		end else begin
			if (andOp_182_out) begin
				icmp_tmp_6 <= cmp_out_icmp_17;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			phi_tmp_1 <= 0;
		end else begin
			if (andOp_179_out) begin
				phi_tmp_1 <= phi_out_phi_8;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (1'd1) begin
				state_0_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_159_out) begin
				state_1_entry_BB_reg <= 32'd0;
			end
			if (andOp_44_out) begin
				state_1_entry_BB_reg <= 32'd9;
			end
			if (andOp_56_out) begin
				state_1_entry_BB_reg <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_159_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_168_out) begin
				state_1_is_active <= 1'd0;
			end
			if (andOp_44_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_56_out) begin
				state_1_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_159_out) begin
				state_1_last_BB_reg <= bb_0_predecessor_in_state_0_out_data;
			end
			if (andOp_44_out) begin
				state_1_last_BB_reg <= 32'd9;
			end
			if (andOp_56_out) begin
				state_1_last_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_159_out) begin
				state_1_last_state <= 32'd0;
			end
			if (andOp_44_out) begin
				state_1_last_state <= 32'd1;
			end
			if (andOp_56_out) begin
				state_1_last_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_42_out) begin
				state_2_entry_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_170_out) begin
				state_2_is_active <= 1'd0;
			end
			if (andOp_42_out) begin
				state_2_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_42_out) begin
				state_2_last_BB_reg <= 32'd9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_42_out) begin
				state_2_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_160_out) begin
				state_3_entry_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_160_out) begin
				state_3_is_active <= 1'd1;
			end
			if (andOp_172_out) begin
				state_3_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_160_out) begin
				state_3_last_BB_reg <= bb_10_predecessor_in_state_2_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_state <= 0;
		end else begin
			if (andOp_160_out) begin
				state_3_last_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_161_out) begin
				state_4_entry_BB_reg <= 32'd4;
			end
			if (andOp_162_out) begin
				state_4_entry_BB_reg <= 32'd2;
			end
			if (andOp_68_out) begin
				state_4_entry_BB_reg <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_161_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_162_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_178_out) begin
				state_4_is_active <= 1'd0;
			end
			if (andOp_68_out) begin
				state_4_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_161_out) begin
				state_4_last_BB_reg <= bb_4_predecessor_in_state_3_out_data;
			end
			if (andOp_162_out) begin
				state_4_last_BB_reg <= bb_2_predecessor_in_state_4_out_data;
			end
			if (andOp_68_out) begin
				state_4_last_BB_reg <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_state <= 0;
		end else begin
			if (andOp_161_out) begin
				state_4_last_state <= 32'd3;
			end
			if (andOp_162_out) begin
				state_4_last_state <= 32'd4;
			end
			if (andOp_68_out) begin
				state_4_last_state <= 32'd4;
			end
		end
	end

endmodule

