module channel_reduce_4(input [0:0] clk, input [0:0] rst, output [0:0] valid, output [31:0] out_in_data, output [0:0] out_read_valid, output [0:0] out_rst, output [0:0] out_write_valid, input [31:0] out_out_data, input [0:0] out_read_ready, input [0:0] out_write_ready, output [31:0] in_in_data, output [0:0] in_read_valid, output [0:0] in_rst, output [0:0] in_write_valid, input [31:0] in_out_data, input [0:0] in_read_ready, input [0:0] in_write_ready);

	reg [0:0] valid_reg;
	reg [31:0] out_in_data_reg;
	reg [0:0] out_read_valid_reg;
	reg [0:0] out_rst_reg;
	reg [0:0] out_write_valid_reg;
	reg [31:0] in_in_data_reg;
	reg [0:0] in_read_valid_reg;
	reg [0:0] in_rst_reg;
	reg [0:0] in_write_valid_reg;

	assign valid = valid_reg;
	assign out_in_data = out_in_data_reg;
	assign out_read_valid = out_read_valid_reg;
	assign out_rst = out_rst_reg;
	assign out_write_valid = out_write_valid_reg;
	assign in_in_data = in_in_data_reg;
	assign in_read_valid = in_read_valid_reg;
	assign in_rst = in_rst_reg;
	assign in_write_valid = in_write_valid_reg;

	// Start debug wires and ports

	initial begin
	end





	// End debug wires and ports

	// Start Functional Units
	add alloca_0();

	add bitcast_1();

	add call_2();

	reg [31:0] raddr_ram_0_reg;
	reg [31:0] waddr_ram_0_reg;
	reg [31:0] wdata_ram_0_reg;
	reg [0:0] wen_ram_0_reg;
	wire [31:0] rdata_ram_0;
	register #(.WIDTH(32)) ram_0(.clk(clk), .raddr(raddr_ram_0_reg), .rdata(rdata_ram_0), .rst(rst), .waddr(waddr_ram_0_reg), .wdata(wdata_ram_0_reg), .wen(wen_ram_0_reg));

	br_dummy br_unit();

	add call_27();

	reg [63:0] phi_in_phi_5;
	reg [31:0] phi_last_block_phi_5;
	reg [63:0] phi_s_phi_5;
	wire [31:0] phi_out_phi_5;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_5(.in(phi_in_phi_5), .last_block(phi_last_block_phi_5), .out(phi_out_phi_5), .s(phi_s_phi_5));

	reg [31:0] add_in0_add_14;
	reg [31:0] add_in1_add_14;
	wire [31:0] add_out_add_14;
	add #(.WIDTH(32)) add_add_14(.in0(add_in0_add_14), .in1(add_in1_add_14), .out(add_out_add_14));

	reg [31:0] add_in0_add_16;
	reg [31:0] add_in1_add_16;
	wire [31:0] add_out_add_16;
	add #(.WIDTH(32)) add_add_16(.in0(add_in0_add_16), .in1(add_in1_add_16), .out(add_out_add_16));

	reg [31:0] cmp_in0_icmp_17;
	reg [31:0] cmp_in1_icmp_17;
	wire [0:0] cmp_out_icmp_17;
	eq #(.WIDTH(32)) icmp_17(.in0(cmp_in0_icmp_17), .in1(cmp_in1_icmp_17), .out(cmp_out_icmp_17));

	reg [0:0] bb_0_active_in_data;
	wire [0:0] bb_0_active_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active(.in_data(bb_0_active_in_data), .out_data(bb_0_active_out_data));

	reg [31:0] eq_0_in0;
	reg [31:0] eq_0_in1;
	wire [0:0] eq_0_out;
	eq #(.WIDTH(32)) eq_0(.in0(eq_0_in0), .in1(eq_0_in1), .out(eq_0_out));

	reg [0:0] andOp_1_in0;
	reg [0:0] andOp_1_in1;
	wire [0:0] andOp_1_out;
	andOp #(.WIDTH(1)) andOp_1(.in0(andOp_1_in0), .in1(andOp_1_in1), .out(andOp_1_out));

	reg [0:0] andOp_2_in0;
	reg [0:0] andOp_2_in1;
	wire [0:0] andOp_2_out;
	andOp #(.WIDTH(1)) andOp_2(.in0(andOp_2_in0), .in1(andOp_2_in1), .out(andOp_2_out));

	reg [0:0] br_0_happened_in_data;
	wire [0:0] br_0_happened_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened(.in_data(br_0_happened_in_data), .out_data(br_0_happened_out_data));

	reg [0:0] notOp_3_in0;
	wire [0:0] notOp_3_out;
	notOp #(.WIDTH(1)) notOp_3(.in(notOp_3_in0), .out(notOp_3_out));

	reg [0:0] bb_1_active_in_data;
	wire [0:0] bb_1_active_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active(.in_data(bb_1_active_in_data), .out_data(bb_1_active_out_data));

	reg [31:0] eq_4_in0;
	reg [31:0] eq_4_in1;
	wire [0:0] eq_4_out;
	eq #(.WIDTH(32)) eq_4(.in0(eq_4_in0), .in1(eq_4_in1), .out(eq_4_out));

	reg [0:0] andOp_5_in0;
	reg [0:0] andOp_5_in1;
	wire [0:0] andOp_5_out;
	andOp #(.WIDTH(1)) andOp_5(.in0(andOp_5_in0), .in1(andOp_5_in1), .out(andOp_5_out));

	reg [0:0] andOp_6_in0;
	reg [0:0] andOp_6_in1;
	wire [0:0] andOp_6_out;
	andOp #(.WIDTH(1)) andOp_6(.in0(andOp_6_in0), .in1(andOp_6_in1), .out(andOp_6_out));

	reg [0:0] br_1_happened_in_data;
	wire [0:0] br_1_happened_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened(.in_data(br_1_happened_in_data), .out_data(br_1_happened_out_data));

	reg [0:0] notOp_7_in0;
	wire [0:0] notOp_7_out;
	notOp #(.WIDTH(1)) notOp_7(.in(notOp_7_in0), .out(notOp_7_out));

	reg [0:0] bb_2_active_in_data;
	wire [0:0] bb_2_active_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active(.in_data(bb_2_active_in_data), .out_data(bb_2_active_out_data));

	reg [0:0] bb_3_active_in_data;
	wire [0:0] bb_3_active_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active(.in_data(bb_3_active_in_data), .out_data(bb_3_active_out_data));

	reg [31:0] eq_8_in0;
	reg [31:0] eq_8_in1;
	wire [0:0] eq_8_out;
	eq #(.WIDTH(32)) eq_8(.in0(eq_8_in0), .in1(eq_8_in1), .out(eq_8_out));

	reg [0:0] andOp_9_in0;
	reg [0:0] andOp_9_in1;
	wire [0:0] andOp_9_out;
	andOp #(.WIDTH(1)) andOp_9(.in0(andOp_9_in0), .in1(andOp_9_in1), .out(andOp_9_out));

	reg [0:0] andOp_10_in0;
	reg [0:0] andOp_10_in1;
	wire [0:0] andOp_10_out;
	andOp #(.WIDTH(1)) andOp_10(.in0(andOp_10_in0), .in1(andOp_10_in1), .out(andOp_10_out));

	reg [0:0] br_3_happened_in_data;
	wire [0:0] br_3_happened_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened(.in_data(br_3_happened_in_data), .out_data(br_3_happened_out_data));

	reg [0:0] notOp_11_in0;
	wire [0:0] notOp_11_out;
	notOp #(.WIDTH(1)) notOp_11(.in(notOp_11_in0), .out(notOp_11_out));

	reg [0:0] bb_4_active_in_data;
	wire [0:0] bb_4_active_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active(.in_data(bb_4_active_in_data), .out_data(bb_4_active_out_data));

	reg [31:0] eq_12_in0;
	reg [31:0] eq_12_in1;
	wire [0:0] eq_12_out;
	eq #(.WIDTH(32)) eq_12(.in0(eq_12_in0), .in1(eq_12_in1), .out(eq_12_out));

	reg [0:0] andOp_13_in0;
	reg [0:0] andOp_13_in1;
	wire [0:0] andOp_13_out;
	andOp #(.WIDTH(1)) andOp_13(.in0(andOp_13_in0), .in1(andOp_13_in1), .out(andOp_13_out));

	reg [0:0] andOp_14_in0;
	reg [0:0] andOp_14_in1;
	wire [0:0] andOp_14_out;
	andOp #(.WIDTH(1)) andOp_14(.in0(andOp_14_in0), .in1(andOp_14_in1), .out(andOp_14_out));

	reg [0:0] br_4_happened_in_data;
	wire [0:0] br_4_happened_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened(.in_data(br_4_happened_in_data), .out_data(br_4_happened_out_data));

	reg [0:0] notOp_15_in0;
	wire [0:0] notOp_15_out;
	notOp #(.WIDTH(1)) notOp_15(.in(notOp_15_in0), .out(notOp_15_out));

	reg [0:0] andOp_16_in0;
	reg [0:0] andOp_16_in1;
	wire [0:0] andOp_16_out;
	andOp #(.WIDTH(1)) andOp_16(.in0(andOp_16_in0), .in1(andOp_16_in1), .out(andOp_16_out));

	reg [0:0] notOp_17_in0;
	wire [0:0] notOp_17_out;
	notOp #(.WIDTH(1)) notOp_17(.in(notOp_17_in0), .out(notOp_17_out));

	reg [0:0] andOp_18_in0;
	reg [0:0] andOp_18_in1;
	wire [0:0] andOp_18_out;
	andOp #(.WIDTH(1)) andOp_18(.in0(andOp_18_in0), .in1(andOp_18_in1), .out(andOp_18_out));

	reg [0:0] bb_5_active_in_data;
	wire [0:0] bb_5_active_out_data;
	hls_wire #(.WIDTH(1)) bb_5_active(.in_data(bb_5_active_in_data), .out_data(bb_5_active_out_data));

	reg [31:0] eq_19_in0;
	reg [31:0] eq_19_in1;
	wire [0:0] eq_19_out;
	eq #(.WIDTH(32)) eq_19(.in0(eq_19_in0), .in1(eq_19_in1), .out(eq_19_out));

	reg [0:0] andOp_20_in0;
	reg [0:0] andOp_20_in1;
	wire [0:0] andOp_20_out;
	andOp #(.WIDTH(1)) andOp_20(.in0(andOp_20_in0), .in1(andOp_20_in1), .out(andOp_20_out));

	reg [0:0] andOp_21_in0;
	reg [0:0] andOp_21_in1;
	wire [0:0] andOp_21_out;
	andOp #(.WIDTH(1)) andOp_21(.in0(andOp_21_in0), .in1(andOp_21_in1), .out(andOp_21_out));

	reg [0:0] br_5_happened_in_data;
	wire [0:0] br_5_happened_out_data;
	hls_wire #(.WIDTH(1)) br_5_happened(.in_data(br_5_happened_in_data), .out_data(br_5_happened_out_data));

	reg [0:0] notOp_22_in0;
	wire [0:0] notOp_22_out;
	notOp #(.WIDTH(1)) notOp_22(.in(notOp_22_in0), .out(notOp_22_out));

	reg [0:0] bb_6_active_in_data;
	wire [0:0] bb_6_active_out_data;
	hls_wire #(.WIDTH(1)) bb_6_active(.in_data(bb_6_active_in_data), .out_data(bb_6_active_out_data));

	reg [31:0] eq_23_in0;
	reg [31:0] eq_23_in1;
	wire [0:0] eq_23_out;
	eq #(.WIDTH(32)) eq_23(.in0(eq_23_in0), .in1(eq_23_in1), .out(eq_23_out));

	reg [0:0] andOp_24_in0;
	reg [0:0] andOp_24_in1;
	wire [0:0] andOp_24_out;
	andOp #(.WIDTH(1)) andOp_24(.in0(andOp_24_in0), .in1(andOp_24_in1), .out(andOp_24_out));

	reg [0:0] andOp_25_in0;
	reg [0:0] andOp_25_in1;
	wire [0:0] andOp_25_out;
	andOp #(.WIDTH(1)) andOp_25(.in0(andOp_25_in0), .in1(andOp_25_in1), .out(andOp_25_out));

	reg [0:0] br_6_happened_in_data;
	wire [0:0] br_6_happened_out_data;
	hls_wire #(.WIDTH(1)) br_6_happened(.in_data(br_6_happened_in_data), .out_data(br_6_happened_out_data));

	reg [0:0] notOp_26_in0;
	wire [0:0] notOp_26_out;
	notOp #(.WIDTH(1)) notOp_26(.in(notOp_26_in0), .out(notOp_26_out));

	reg [0:0] andOp_27_in0;
	reg [0:0] andOp_27_in1;
	wire [0:0] andOp_27_out;
	andOp #(.WIDTH(1)) andOp_27(.in0(andOp_27_in0), .in1(andOp_27_in1), .out(andOp_27_out));

	reg [0:0] notOp_28_in0;
	wire [0:0] notOp_28_out;
	notOp #(.WIDTH(1)) notOp_28(.in(notOp_28_in0), .out(notOp_28_out));

	reg [0:0] andOp_29_in0;
	reg [0:0] andOp_29_in1;
	wire [0:0] andOp_29_out;
	andOp #(.WIDTH(1)) andOp_29(.in0(andOp_29_in0), .in1(andOp_29_in1), .out(andOp_29_out));

	reg [0:0] bb_7_active_in_data;
	wire [0:0] bb_7_active_out_data;
	hls_wire #(.WIDTH(1)) bb_7_active(.in_data(bb_7_active_in_data), .out_data(bb_7_active_out_data));

	reg [31:0] eq_30_in0;
	reg [31:0] eq_30_in1;
	wire [0:0] eq_30_out;
	eq #(.WIDTH(32)) eq_30(.in0(eq_30_in0), .in1(eq_30_in1), .out(eq_30_out));

	reg [0:0] andOp_31_in0;
	reg [0:0] andOp_31_in1;
	wire [0:0] andOp_31_out;
	andOp #(.WIDTH(1)) andOp_31(.in0(andOp_31_in0), .in1(andOp_31_in1), .out(andOp_31_out));

	reg [0:0] andOp_32_in0;
	reg [0:0] andOp_32_in1;
	wire [0:0] andOp_32_out;
	andOp #(.WIDTH(1)) andOp_32(.in0(andOp_32_in0), .in1(andOp_32_in1), .out(andOp_32_out));

	reg [0:0] br_7_happened_in_data;
	wire [0:0] br_7_happened_out_data;
	hls_wire #(.WIDTH(1)) br_7_happened(.in_data(br_7_happened_in_data), .out_data(br_7_happened_out_data));

	reg [0:0] notOp_33_in0;
	wire [0:0] notOp_33_out;
	notOp #(.WIDTH(1)) notOp_33(.in(notOp_33_in0), .out(notOp_33_out));

	reg [0:0] bb_8_active_in_data;
	wire [0:0] bb_8_active_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active(.in_data(bb_8_active_in_data), .out_data(bb_8_active_out_data));

	reg [31:0] eq_34_in0;
	reg [31:0] eq_34_in1;
	wire [0:0] eq_34_out;
	eq #(.WIDTH(32)) eq_34(.in0(eq_34_in0), .in1(eq_34_in1), .out(eq_34_out));

	reg [0:0] andOp_35_in0;
	reg [0:0] andOp_35_in1;
	wire [0:0] andOp_35_out;
	andOp #(.WIDTH(1)) andOp_35(.in0(andOp_35_in0), .in1(andOp_35_in1), .out(andOp_35_out));

	reg [0:0] andOp_36_in0;
	reg [0:0] andOp_36_in1;
	wire [0:0] andOp_36_out;
	andOp #(.WIDTH(1)) andOp_36(.in0(andOp_36_in0), .in1(andOp_36_in1), .out(andOp_36_out));

	reg [0:0] br_8_happened_in_data;
	wire [0:0] br_8_happened_out_data;
	hls_wire #(.WIDTH(1)) br_8_happened(.in_data(br_8_happened_in_data), .out_data(br_8_happened_out_data));

	reg [0:0] notOp_37_in0;
	wire [0:0] notOp_37_out;
	notOp #(.WIDTH(1)) notOp_37(.in(notOp_37_in0), .out(notOp_37_out));

	reg [0:0] bb_9_active_in_data;
	wire [0:0] bb_9_active_out_data;
	hls_wire #(.WIDTH(1)) bb_9_active(.in_data(bb_9_active_in_data), .out_data(bb_9_active_out_data));

	reg [31:0] eq_38_in0;
	reg [31:0] eq_38_in1;
	wire [0:0] eq_38_out;
	eq #(.WIDTH(32)) eq_38(.in0(eq_38_in0), .in1(eq_38_in1), .out(eq_38_out));

	reg [0:0] andOp_39_in0;
	reg [0:0] andOp_39_in1;
	wire [0:0] andOp_39_out;
	andOp #(.WIDTH(1)) andOp_39(.in0(andOp_39_in0), .in1(andOp_39_in1), .out(andOp_39_out));

	reg [0:0] andOp_40_in0;
	reg [0:0] andOp_40_in1;
	wire [0:0] andOp_40_out;
	andOp #(.WIDTH(1)) andOp_40(.in0(andOp_40_in0), .in1(andOp_40_in1), .out(andOp_40_out));

	reg [0:0] br_9_happened_in_data;
	wire [0:0] br_9_happened_out_data;
	hls_wire #(.WIDTH(1)) br_9_happened(.in_data(br_9_happened_in_data), .out_data(br_9_happened_out_data));

	reg [0:0] notOp_41_in0;
	wire [0:0] notOp_41_out;
	notOp #(.WIDTH(1)) notOp_41(.in(notOp_41_in0), .out(notOp_41_out));

	reg [0:0] andOp_42_in0;
	reg [0:0] andOp_42_in1;
	wire [0:0] andOp_42_out;
	andOp #(.WIDTH(1)) andOp_42(.in0(andOp_42_in0), .in1(andOp_42_in1), .out(andOp_42_out));

	reg [0:0] notOp_43_in0;
	wire [0:0] notOp_43_out;
	notOp #(.WIDTH(1)) notOp_43(.in(notOp_43_in0), .out(notOp_43_out));

	reg [0:0] andOp_44_in0;
	reg [0:0] andOp_44_in1;
	wire [0:0] andOp_44_out;
	andOp #(.WIDTH(1)) andOp_44(.in0(andOp_44_in0), .in1(andOp_44_in1), .out(andOp_44_out));

	reg [0:0] bb_10_active_in_data;
	wire [0:0] bb_10_active_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active(.in_data(bb_10_active_in_data), .out_data(bb_10_active_out_data));

	reg [31:0] eq_45_in0;
	reg [31:0] eq_45_in1;
	wire [0:0] eq_45_out;
	eq #(.WIDTH(32)) eq_45(.in0(eq_45_in0), .in1(eq_45_in1), .out(eq_45_out));

	reg [0:0] andOp_46_in0;
	reg [0:0] andOp_46_in1;
	wire [0:0] andOp_46_out;
	andOp #(.WIDTH(1)) andOp_46(.in0(andOp_46_in0), .in1(andOp_46_in1), .out(andOp_46_out));

	reg [0:0] andOp_47_in0;
	reg [0:0] andOp_47_in1;
	wire [0:0] andOp_47_out;
	andOp #(.WIDTH(1)) andOp_47(.in0(andOp_47_in0), .in1(andOp_47_in1), .out(andOp_47_out));

	reg [0:0] br_10_happened_in_data;
	wire [0:0] br_10_happened_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened(.in_data(br_10_happened_in_data), .out_data(br_10_happened_out_data));

	reg [0:0] notOp_48_in0;
	wire [0:0] notOp_48_out;
	notOp #(.WIDTH(1)) notOp_48(.in(notOp_48_in0), .out(notOp_48_out));

	reg [31:0] eq_49_in0;
	reg [31:0] eq_49_in1;
	wire [0:0] eq_49_out;
	eq #(.WIDTH(32)) eq_49(.in0(eq_49_in0), .in1(eq_49_in1), .out(eq_49_out));

	reg [31:0] eq_50_in0;
	reg [31:0] eq_50_in1;
	wire [0:0] eq_50_out;
	eq #(.WIDTH(32)) eq_50(.in0(eq_50_in0), .in1(eq_50_in1), .out(eq_50_out));

	reg [0:0] orOp_51_in0;
	reg [0:0] orOp_51_in1;
	wire [0:0] orOp_51_out;
	orOp #(.WIDTH(1)) orOp_51(.in0(orOp_51_in0), .in1(orOp_51_in1), .out(orOp_51_out));

	reg [31:0] eq_52_in0;
	reg [31:0] eq_52_in1;
	wire [0:0] eq_52_out;
	eq #(.WIDTH(32)) eq_52(.in0(eq_52_in0), .in1(eq_52_in1), .out(eq_52_out));

	reg [31:0] eq_53_in0;
	reg [31:0] eq_53_in1;
	wire [0:0] eq_53_out;
	eq #(.WIDTH(32)) eq_53(.in0(eq_53_in0), .in1(eq_53_in1), .out(eq_53_out));

	reg [0:0] orOp_54_in0;
	reg [0:0] orOp_54_in1;
	wire [0:0] orOp_54_out;
	orOp #(.WIDTH(1)) orOp_54(.in0(orOp_54_in0), .in1(orOp_54_in1), .out(orOp_54_out));

	reg [31:0] eq_55_in0;
	reg [31:0] eq_55_in1;
	wire [0:0] eq_55_out;
	eq #(.WIDTH(32)) eq_55(.in0(eq_55_in0), .in1(eq_55_in1), .out(eq_55_out));

	reg [31:0] eq_56_in0;
	reg [31:0] eq_56_in1;
	wire [0:0] eq_56_out;
	eq #(.WIDTH(32)) eq_56(.in0(eq_56_in0), .in1(eq_56_in1), .out(eq_56_out));

	reg [0:0] orOp_57_in0;
	reg [0:0] orOp_57_in1;
	wire [0:0] orOp_57_out;
	orOp #(.WIDTH(1)) orOp_57(.in0(orOp_57_in0), .in1(orOp_57_in1), .out(orOp_57_out));

	reg [31:0] eq_58_in0;
	reg [31:0] eq_58_in1;
	wire [0:0] eq_58_out;
	eq #(.WIDTH(32)) eq_58(.in0(eq_58_in0), .in1(eq_58_in1), .out(eq_58_out));

	reg [31:0] eq_59_in0;
	reg [31:0] eq_59_in1;
	wire [0:0] eq_59_out;
	eq #(.WIDTH(32)) eq_59(.in0(eq_59_in0), .in1(eq_59_in1), .out(eq_59_out));

	reg [31:0] eq_60_in0;
	reg [31:0] eq_60_in1;
	wire [0:0] eq_60_out;
	eq #(.WIDTH(32)) eq_60(.in0(eq_60_in0), .in1(eq_60_in1), .out(eq_60_out));

	reg [0:0] orOp_61_in0;
	reg [0:0] orOp_61_in1;
	wire [0:0] orOp_61_out;
	orOp #(.WIDTH(1)) orOp_61(.in0(orOp_61_in0), .in1(orOp_61_in1), .out(orOp_61_out));

	reg [31:0] eq_62_in0;
	reg [31:0] eq_62_in1;
	wire [0:0] eq_62_out;
	eq #(.WIDTH(32)) eq_62(.in0(eq_62_in0), .in1(eq_62_in1), .out(eq_62_out));

	reg [31:0] eq_63_in0;
	reg [31:0] eq_63_in1;
	wire [0:0] eq_63_out;
	eq #(.WIDTH(32)) eq_63(.in0(eq_63_in0), .in1(eq_63_in1), .out(eq_63_out));

	reg [31:0] eq_64_in0;
	reg [31:0] eq_64_in1;
	wire [0:0] eq_64_out;
	eq #(.WIDTH(32)) eq_64(.in0(eq_64_in0), .in1(eq_64_in1), .out(eq_64_out));

	reg [0:0] andOp_65_in0;
	reg [0:0] andOp_65_in1;
	wire [0:0] andOp_65_out;
	andOp #(.WIDTH(1)) andOp_65(.in0(andOp_65_in0), .in1(andOp_65_in1), .out(andOp_65_out));

	reg [31:0] eq_66_in0;
	reg [31:0] eq_66_in1;
	wire [0:0] eq_66_out;
	eq #(.WIDTH(32)) eq_66(.in0(eq_66_in0), .in1(eq_66_in1), .out(eq_66_out));

	reg [0:0] andOp_67_in0;
	reg [0:0] andOp_67_in1;
	wire [0:0] andOp_67_out;
	andOp #(.WIDTH(1)) andOp_67(.in0(andOp_67_in0), .in1(andOp_67_in1), .out(andOp_67_out));

	reg [31:0] eq_68_in0;
	reg [31:0] eq_68_in1;
	wire [0:0] eq_68_out;
	eq #(.WIDTH(32)) eq_68(.in0(eq_68_in0), .in1(eq_68_in1), .out(eq_68_out));

	reg [0:0] andOp_69_in0;
	reg [0:0] andOp_69_in1;
	wire [0:0] andOp_69_out;
	andOp #(.WIDTH(1)) andOp_69(.in0(andOp_69_in0), .in1(andOp_69_in1), .out(andOp_69_out));

	reg [31:0] eq_70_in0;
	reg [31:0] eq_70_in1;
	wire [0:0] eq_70_out;
	eq #(.WIDTH(32)) eq_70(.in0(eq_70_in0), .in1(eq_70_in1), .out(eq_70_out));

	reg [0:0] andOp_71_in0;
	reg [0:0] andOp_71_in1;
	wire [0:0] andOp_71_out;
	andOp #(.WIDTH(1)) andOp_71(.in0(andOp_71_in0), .in1(andOp_71_in1), .out(andOp_71_out));

	reg [31:0] bb_0_predecessor_in_data;
	wire [31:0] bb_0_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor(.in_data(bb_0_predecessor_in_data), .out_data(bb_0_predecessor_out_data));

	reg [31:0] eq_72_in0;
	reg [31:0] eq_72_in1;
	wire [0:0] eq_72_out;
	eq #(.WIDTH(32)) eq_72(.in0(eq_72_in0), .in1(eq_72_in1), .out(eq_72_out));

	reg [31:0] bb_1_predecessor_in_data;
	wire [31:0] bb_1_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor(.in_data(bb_1_predecessor_in_data), .out_data(bb_1_predecessor_out_data));

	reg [31:0] eq_73_in0;
	reg [31:0] eq_73_in1;
	wire [0:0] eq_73_out;
	eq #(.WIDTH(32)) eq_73(.in0(eq_73_in0), .in1(eq_73_in1), .out(eq_73_out));

	reg [0:0] notOp_74_in0;
	wire [0:0] notOp_74_out;
	notOp #(.WIDTH(1)) notOp_74(.in(notOp_74_in0), .out(notOp_74_out));

	reg [0:0] andOp_75_in0;
	reg [0:0] andOp_75_in1;
	wire [0:0] andOp_75_out;
	andOp #(.WIDTH(1)) andOp_75(.in0(andOp_75_in0), .in1(andOp_75_in1), .out(andOp_75_out));

	reg [31:0] bb_2_predecessor_in_data;
	wire [31:0] bb_2_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor(.in_data(bb_2_predecessor_in_data), .out_data(bb_2_predecessor_out_data));

	reg [31:0] eq_76_in0;
	reg [31:0] eq_76_in1;
	wire [0:0] eq_76_out;
	eq #(.WIDTH(32)) eq_76(.in0(eq_76_in0), .in1(eq_76_in1), .out(eq_76_out));

	reg [31:0] bb_3_predecessor_in_data;
	wire [31:0] bb_3_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor(.in_data(bb_3_predecessor_in_data), .out_data(bb_3_predecessor_out_data));

	reg [31:0] eq_77_in0;
	reg [31:0] eq_77_in1;
	wire [0:0] eq_77_out;
	eq #(.WIDTH(32)) eq_77(.in0(eq_77_in0), .in1(eq_77_in1), .out(eq_77_out));

	reg [0:0] notOp_78_in0;
	wire [0:0] notOp_78_out;
	notOp #(.WIDTH(1)) notOp_78(.in(notOp_78_in0), .out(notOp_78_out));

	reg [0:0] andOp_79_in0;
	reg [0:0] andOp_79_in1;
	wire [0:0] andOp_79_out;
	andOp #(.WIDTH(1)) andOp_79(.in0(andOp_79_in0), .in1(andOp_79_in1), .out(andOp_79_out));

	reg [31:0] bb_4_predecessor_in_data;
	wire [31:0] bb_4_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor(.in_data(bb_4_predecessor_in_data), .out_data(bb_4_predecessor_out_data));

	reg [31:0] eq_80_in0;
	reg [31:0] eq_80_in1;
	wire [0:0] eq_80_out;
	eq #(.WIDTH(32)) eq_80(.in0(eq_80_in0), .in1(eq_80_in1), .out(eq_80_out));

	reg [31:0] bb_5_predecessor_in_data;
	wire [31:0] bb_5_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_5_predecessor(.in_data(bb_5_predecessor_in_data), .out_data(bb_5_predecessor_out_data));

	reg [31:0] eq_81_in0;
	reg [31:0] eq_81_in1;
	wire [0:0] eq_81_out;
	eq #(.WIDTH(32)) eq_81(.in0(eq_81_in0), .in1(eq_81_in1), .out(eq_81_out));

	reg [0:0] notOp_82_in0;
	wire [0:0] notOp_82_out;
	notOp #(.WIDTH(1)) notOp_82(.in(notOp_82_in0), .out(notOp_82_out));

	reg [0:0] andOp_83_in0;
	reg [0:0] andOp_83_in1;
	wire [0:0] andOp_83_out;
	andOp #(.WIDTH(1)) andOp_83(.in0(andOp_83_in0), .in1(andOp_83_in1), .out(andOp_83_out));

	reg [31:0] bb_6_predecessor_in_data;
	wire [31:0] bb_6_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_6_predecessor(.in_data(bb_6_predecessor_in_data), .out_data(bb_6_predecessor_out_data));

	reg [31:0] eq_84_in0;
	reg [31:0] eq_84_in1;
	wire [0:0] eq_84_out;
	eq #(.WIDTH(32)) eq_84(.in0(eq_84_in0), .in1(eq_84_in1), .out(eq_84_out));

	reg [31:0] bb_7_predecessor_in_data;
	wire [31:0] bb_7_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_7_predecessor(.in_data(bb_7_predecessor_in_data), .out_data(bb_7_predecessor_out_data));

	reg [31:0] eq_85_in0;
	reg [31:0] eq_85_in1;
	wire [0:0] eq_85_out;
	eq #(.WIDTH(32)) eq_85(.in0(eq_85_in0), .in1(eq_85_in1), .out(eq_85_out));

	reg [31:0] bb_8_predecessor_in_data;
	wire [31:0] bb_8_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor(.in_data(bb_8_predecessor_in_data), .out_data(bb_8_predecessor_out_data));

	reg [31:0] eq_86_in0;
	reg [31:0] eq_86_in1;
	wire [0:0] eq_86_out;
	eq #(.WIDTH(32)) eq_86(.in0(eq_86_in0), .in1(eq_86_in1), .out(eq_86_out));

	reg [0:0] notOp_87_in0;
	wire [0:0] notOp_87_out;
	notOp #(.WIDTH(1)) notOp_87(.in(notOp_87_in0), .out(notOp_87_out));

	reg [0:0] andOp_88_in0;
	reg [0:0] andOp_88_in1;
	wire [0:0] andOp_88_out;
	andOp #(.WIDTH(1)) andOp_88(.in0(andOp_88_in0), .in1(andOp_88_in1), .out(andOp_88_out));

	reg [31:0] bb_9_predecessor_in_data;
	wire [31:0] bb_9_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_9_predecessor(.in_data(bb_9_predecessor_in_data), .out_data(bb_9_predecessor_out_data));

	reg [31:0] eq_89_in0;
	reg [31:0] eq_89_in1;
	wire [0:0] eq_89_out;
	eq #(.WIDTH(32)) eq_89(.in0(eq_89_in0), .in1(eq_89_in1), .out(eq_89_out));

	reg [31:0] bb_10_predecessor_in_data;
	wire [31:0] bb_10_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor(.in_data(bb_10_predecessor_in_data), .out_data(bb_10_predecessor_out_data));

	reg [31:0] eq_90_in0;
	reg [31:0] eq_90_in1;
	wire [0:0] eq_90_out;
	eq #(.WIDTH(32)) eq_90(.in0(eq_90_in0), .in1(eq_90_in1), .out(eq_90_out));

	reg [31:0] eq_91_in0;
	reg [31:0] eq_91_in1;
	wire [0:0] eq_91_out;
	eq #(.WIDTH(32)) eq_91(.in0(eq_91_in0), .in1(eq_91_in1), .out(eq_91_out));

	reg [0:0] andOp_92_in0;
	reg [0:0] andOp_92_in1;
	wire [0:0] andOp_92_out;
	andOp #(.WIDTH(1)) andOp_92(.in0(andOp_92_in0), .in1(andOp_92_in1), .out(andOp_92_out));

	reg [31:0] eq_93_in0;
	reg [31:0] eq_93_in1;
	wire [0:0] eq_93_out;
	eq #(.WIDTH(32)) eq_93(.in0(eq_93_in0), .in1(eq_93_in1), .out(eq_93_out));

	reg [0:0] andOp_94_in0;
	reg [0:0] andOp_94_in1;
	wire [0:0] andOp_94_out;
	andOp #(.WIDTH(1)) andOp_94(.in0(andOp_94_in0), .in1(andOp_94_in1), .out(andOp_94_out));

	reg [31:0] eq_95_in0;
	reg [31:0] eq_95_in1;
	wire [0:0] eq_95_out;
	eq #(.WIDTH(32)) eq_95(.in0(eq_95_in0), .in1(eq_95_in1), .out(eq_95_out));

	reg [0:0] andOp_96_in0;
	reg [0:0] andOp_96_in1;
	wire [0:0] andOp_96_out;
	andOp #(.WIDTH(1)) andOp_96(.in0(andOp_96_in0), .in1(andOp_96_in1), .out(andOp_96_out));

	reg [31:0] eq_97_in0;
	reg [31:0] eq_97_in1;
	wire [0:0] eq_97_out;
	eq #(.WIDTH(32)) eq_97(.in0(eq_97_in0), .in1(eq_97_in1), .out(eq_97_out));

	reg [0:0] andOp_98_in0;
	reg [0:0] andOp_98_in1;
	wire [0:0] andOp_98_out;
	andOp #(.WIDTH(1)) andOp_98(.in0(andOp_98_in0), .in1(andOp_98_in1), .out(andOp_98_out));

	reg [31:0] eq_99_in0;
	reg [31:0] eq_99_in1;
	wire [0:0] eq_99_out;
	eq #(.WIDTH(32)) eq_99(.in0(eq_99_in0), .in1(eq_99_in1), .out(eq_99_out));

	reg [0:0] andOp_100_in0;
	reg [0:0] andOp_100_in1;
	wire [0:0] andOp_100_out;
	andOp #(.WIDTH(1)) andOp_100(.in0(andOp_100_in0), .in1(andOp_100_in1), .out(andOp_100_out));

	reg [31:0] eq_101_in0;
	reg [31:0] eq_101_in1;
	wire [0:0] eq_101_out;
	eq #(.WIDTH(32)) eq_101(.in0(eq_101_in0), .in1(eq_101_in1), .out(eq_101_out));

	reg [0:0] andOp_102_in0;
	reg [0:0] andOp_102_in1;
	wire [0:0] andOp_102_out;
	andOp #(.WIDTH(1)) andOp_102(.in0(andOp_102_in0), .in1(andOp_102_in1), .out(andOp_102_out));

	reg [31:0] eq_103_in0;
	reg [31:0] eq_103_in1;
	wire [0:0] eq_103_out;
	eq #(.WIDTH(32)) eq_103(.in0(eq_103_in0), .in1(eq_103_in1), .out(eq_103_out));

	reg [0:0] andOp_104_in0;
	reg [0:0] andOp_104_in1;
	wire [0:0] andOp_104_out;
	andOp #(.WIDTH(1)) andOp_104(.in0(andOp_104_in0), .in1(andOp_104_in1), .out(andOp_104_out));

	reg [31:0] eq_105_in0;
	reg [31:0] eq_105_in1;
	wire [0:0] eq_105_out;
	eq #(.WIDTH(32)) eq_105(.in0(eq_105_in0), .in1(eq_105_in1), .out(eq_105_out));

	reg [0:0] andOp_106_in0;
	reg [0:0] andOp_106_in1;
	wire [0:0] andOp_106_out;
	andOp #(.WIDTH(1)) andOp_106(.in0(andOp_106_in0), .in1(andOp_106_in1), .out(andOp_106_out));

	reg [31:0] eq_107_in0;
	reg [31:0] eq_107_in1;
	wire [0:0] eq_107_out;
	eq #(.WIDTH(32)) eq_107(.in0(eq_107_in0), .in1(eq_107_in1), .out(eq_107_out));

	reg [0:0] andOp_108_in0;
	reg [0:0] andOp_108_in1;
	wire [0:0] andOp_108_out;
	andOp #(.WIDTH(1)) andOp_108(.in0(andOp_108_in0), .in1(andOp_108_in1), .out(andOp_108_out));

	reg [31:0] eq_109_in0;
	reg [31:0] eq_109_in1;
	wire [0:0] eq_109_out;
	eq #(.WIDTH(32)) eq_109(.in0(eq_109_in0), .in1(eq_109_in1), .out(eq_109_out));

	reg [0:0] andOp_110_in0;
	reg [0:0] andOp_110_in1;
	wire [0:0] andOp_110_out;
	andOp #(.WIDTH(1)) andOp_110(.in0(andOp_110_in0), .in1(andOp_110_in1), .out(andOp_110_out));

	reg [31:0] eq_111_in0;
	reg [31:0] eq_111_in1;
	wire [0:0] eq_111_out;
	eq #(.WIDTH(32)) eq_111(.in0(eq_111_in0), .in1(eq_111_in1), .out(eq_111_out));

	reg [0:0] andOp_112_in0;
	reg [0:0] andOp_112_in1;
	wire [0:0] andOp_112_out;
	andOp #(.WIDTH(1)) andOp_112(.in0(andOp_112_in0), .in1(andOp_112_in1), .out(andOp_112_out));

	reg [31:0] eq_113_in0;
	reg [31:0] eq_113_in1;
	wire [0:0] eq_113_out;
	eq #(.WIDTH(32)) eq_113(.in0(eq_113_in0), .in1(eq_113_in1), .out(eq_113_out));

	reg [0:0] andOp_114_in0;
	reg [0:0] andOp_114_in1;
	wire [0:0] andOp_114_out;
	andOp #(.WIDTH(1)) andOp_114(.in0(andOp_114_in0), .in1(andOp_114_in1), .out(andOp_114_out));

	reg [31:0] eq_115_in0;
	reg [31:0] eq_115_in1;
	wire [0:0] eq_115_out;
	eq #(.WIDTH(32)) eq_115(.in0(eq_115_in0), .in1(eq_115_in1), .out(eq_115_out));

	reg [0:0] andOp_116_in0;
	reg [0:0] andOp_116_in1;
	wire [0:0] andOp_116_out;
	andOp #(.WIDTH(1)) andOp_116(.in0(andOp_116_in0), .in1(andOp_116_in1), .out(andOp_116_out));

	reg [31:0] eq_117_in0;
	reg [31:0] eq_117_in1;
	wire [0:0] eq_117_out;
	eq #(.WIDTH(32)) eq_117(.in0(eq_117_in0), .in1(eq_117_in1), .out(eq_117_out));

	reg [0:0] andOp_118_in0;
	reg [0:0] andOp_118_in1;
	wire [0:0] andOp_118_out;
	andOp #(.WIDTH(1)) andOp_118(.in0(andOp_118_in0), .in1(andOp_118_in1), .out(andOp_118_out));

	reg [31:0] eq_119_in0;
	reg [31:0] eq_119_in1;
	wire [0:0] eq_119_out;
	eq #(.WIDTH(32)) eq_119(.in0(eq_119_in0), .in1(eq_119_in1), .out(eq_119_out));

	reg [0:0] andOp_120_in0;
	reg [0:0] andOp_120_in1;
	wire [0:0] andOp_120_out;
	andOp #(.WIDTH(1)) andOp_120(.in0(andOp_120_in0), .in1(andOp_120_in1), .out(andOp_120_out));

	reg [31:0] eq_121_in0;
	reg [31:0] eq_121_in1;
	wire [0:0] eq_121_out;
	eq #(.WIDTH(32)) eq_121(.in0(eq_121_in0), .in1(eq_121_in1), .out(eq_121_out));

	reg [0:0] andOp_122_in0;
	reg [0:0] andOp_122_in1;
	wire [0:0] andOp_122_out;
	andOp #(.WIDTH(1)) andOp_122(.in0(andOp_122_in0), .in1(andOp_122_in1), .out(andOp_122_out));

	reg [31:0] eq_123_in0;
	reg [31:0] eq_123_in1;
	wire [0:0] eq_123_out;
	eq #(.WIDTH(32)) eq_123(.in0(eq_123_in0), .in1(eq_123_in1), .out(eq_123_out));

	reg [0:0] andOp_124_in0;
	reg [0:0] andOp_124_in1;
	wire [0:0] andOp_124_out;
	andOp #(.WIDTH(1)) andOp_124(.in0(andOp_124_in0), .in1(andOp_124_in1), .out(andOp_124_out));

	reg [31:0] eq_125_in0;
	reg [31:0] eq_125_in1;
	wire [0:0] eq_125_out;
	eq #(.WIDTH(32)) eq_125(.in0(eq_125_in0), .in1(eq_125_in1), .out(eq_125_out));

	reg [0:0] andOp_126_in0;
	reg [0:0] andOp_126_in1;
	wire [0:0] andOp_126_out;
	andOp #(.WIDTH(1)) andOp_126(.in0(andOp_126_in0), .in1(andOp_126_in1), .out(andOp_126_out));

	reg [31:0] eq_127_in0;
	reg [31:0] eq_127_in1;
	wire [0:0] eq_127_out;
	eq #(.WIDTH(32)) eq_127(.in0(eq_127_in0), .in1(eq_127_in1), .out(eq_127_out));

	reg [0:0] andOp_128_in0;
	reg [0:0] andOp_128_in1;
	wire [0:0] andOp_128_out;
	andOp #(.WIDTH(1)) andOp_128(.in0(andOp_128_in0), .in1(andOp_128_in1), .out(andOp_128_out));

	reg [31:0] eq_129_in0;
	reg [31:0] eq_129_in1;
	wire [0:0] eq_129_out;
	eq #(.WIDTH(32)) eq_129(.in0(eq_129_in0), .in1(eq_129_in1), .out(eq_129_out));

	reg [0:0] andOp_130_in0;
	reg [0:0] andOp_130_in1;
	wire [0:0] andOp_130_out;
	andOp #(.WIDTH(1)) andOp_130(.in0(andOp_130_in0), .in1(andOp_130_in1), .out(andOp_130_out));

	reg [31:0] eq_131_in0;
	reg [31:0] eq_131_in1;
	wire [0:0] eq_131_out;
	eq #(.WIDTH(32)) eq_131(.in0(eq_131_in0), .in1(eq_131_in1), .out(eq_131_out));

	reg [0:0] andOp_132_in0;
	reg [0:0] andOp_132_in1;
	wire [0:0] andOp_132_out;
	andOp #(.WIDTH(1)) andOp_132(.in0(andOp_132_in0), .in1(andOp_132_in1), .out(andOp_132_out));

	reg [0:0] notOp_133_in0;
	wire [0:0] notOp_133_out;
	notOp #(.WIDTH(1)) notOp_133(.in(notOp_133_in0), .out(notOp_133_out));

	reg [0:0] andOp_134_in0;
	reg [0:0] andOp_134_in1;
	wire [0:0] andOp_134_out;
	andOp #(.WIDTH(1)) andOp_134(.in0(andOp_134_in0), .in1(andOp_134_in1), .out(andOp_134_out));

	reg [31:0] eq_135_in0;
	reg [31:0] eq_135_in1;
	wire [0:0] eq_135_out;
	eq #(.WIDTH(32)) eq_135(.in0(eq_135_in0), .in1(eq_135_in1), .out(eq_135_out));

	reg [0:0] andOp_136_in0;
	reg [0:0] andOp_136_in1;
	wire [0:0] andOp_136_out;
	andOp #(.WIDTH(1)) andOp_136(.in0(andOp_136_in0), .in1(andOp_136_in1), .out(andOp_136_out));

	reg [31:0] eq_137_in0;
	reg [31:0] eq_137_in1;
	wire [0:0] eq_137_out;
	eq #(.WIDTH(32)) eq_137(.in0(eq_137_in0), .in1(eq_137_in1), .out(eq_137_out));

	reg [0:0] andOp_138_in0;
	reg [0:0] andOp_138_in1;
	wire [0:0] andOp_138_out;
	andOp #(.WIDTH(1)) andOp_138(.in0(andOp_138_in0), .in1(andOp_138_in1), .out(andOp_138_out));

	reg [0:0] notOp_139_in0;
	wire [0:0] notOp_139_out;
	notOp #(.WIDTH(1)) notOp_139(.in(notOp_139_in0), .out(notOp_139_out));

	reg [0:0] andOp_140_in0;
	reg [0:0] andOp_140_in1;
	wire [0:0] andOp_140_out;
	andOp #(.WIDTH(1)) andOp_140(.in0(andOp_140_in0), .in1(andOp_140_in1), .out(andOp_140_out));

	reg [31:0] eq_141_in0;
	reg [31:0] eq_141_in1;
	wire [0:0] eq_141_out;
	eq #(.WIDTH(32)) eq_141(.in0(eq_141_in0), .in1(eq_141_in1), .out(eq_141_out));

	reg [0:0] andOp_142_in0;
	reg [0:0] andOp_142_in1;
	wire [0:0] andOp_142_out;
	andOp #(.WIDTH(1)) andOp_142(.in0(andOp_142_in0), .in1(andOp_142_in1), .out(andOp_142_out));

	reg [31:0] eq_143_in0;
	reg [31:0] eq_143_in1;
	wire [0:0] eq_143_out;
	eq #(.WIDTH(32)) eq_143(.in0(eq_143_in0), .in1(eq_143_in1), .out(eq_143_out));

	reg [0:0] andOp_144_in0;
	reg [0:0] andOp_144_in1;
	wire [0:0] andOp_144_out;
	andOp #(.WIDTH(1)) andOp_144(.in0(andOp_144_in0), .in1(andOp_144_in1), .out(andOp_144_out));

	reg [0:0] notOp_145_in0;
	wire [0:0] notOp_145_out;
	notOp #(.WIDTH(1)) notOp_145(.in(notOp_145_in0), .out(notOp_145_out));

	reg [0:0] andOp_146_in0;
	reg [0:0] andOp_146_in1;
	wire [0:0] andOp_146_out;
	andOp #(.WIDTH(1)) andOp_146(.in0(andOp_146_in0), .in1(andOp_146_in1), .out(andOp_146_out));

	reg [31:0] eq_147_in0;
	reg [31:0] eq_147_in1;
	wire [0:0] eq_147_out;
	eq #(.WIDTH(32)) eq_147(.in0(eq_147_in0), .in1(eq_147_in1), .out(eq_147_out));

	reg [0:0] andOp_148_in0;
	reg [0:0] andOp_148_in1;
	wire [0:0] andOp_148_out;
	andOp #(.WIDTH(1)) andOp_148(.in0(andOp_148_in0), .in1(andOp_148_in1), .out(andOp_148_out));

	reg [31:0] eq_149_in0;
	reg [31:0] eq_149_in1;
	wire [0:0] eq_149_out;
	eq #(.WIDTH(32)) eq_149(.in0(eq_149_in0), .in1(eq_149_in1), .out(eq_149_out));

	reg [0:0] andOp_150_in0;
	reg [0:0] andOp_150_in1;
	wire [0:0] andOp_150_out;
	andOp #(.WIDTH(1)) andOp_150(.in0(andOp_150_in0), .in1(andOp_150_in1), .out(andOp_150_out));

	reg [0:0] notOp_151_in0;
	wire [0:0] notOp_151_out;
	notOp #(.WIDTH(1)) notOp_151(.in(notOp_151_in0), .out(notOp_151_out));

	reg [0:0] andOp_152_in0;
	reg [0:0] andOp_152_in1;
	wire [0:0] andOp_152_out;
	andOp #(.WIDTH(1)) andOp_152(.in0(andOp_152_in0), .in1(andOp_152_in1), .out(andOp_152_out));

	reg [31:0] eq_153_in0;
	reg [31:0] eq_153_in1;
	wire [0:0] eq_153_out;
	eq #(.WIDTH(32)) eq_153(.in0(eq_153_in0), .in1(eq_153_in1), .out(eq_153_out));

	reg [0:0] andOp_154_in0;
	reg [0:0] andOp_154_in1;
	wire [0:0] andOp_154_out;
	andOp #(.WIDTH(1)) andOp_154(.in0(andOp_154_in0), .in1(andOp_154_in1), .out(andOp_154_out));

	reg [31:0] eq_155_in0;
	reg [31:0] eq_155_in1;
	wire [0:0] eq_155_out;
	eq #(.WIDTH(32)) eq_155(.in0(eq_155_in0), .in1(eq_155_in1), .out(eq_155_out));

	reg [0:0] andOp_156_in0;
	reg [0:0] andOp_156_in1;
	wire [0:0] andOp_156_out;
	andOp #(.WIDTH(1)) andOp_156(.in0(andOp_156_in0), .in1(andOp_156_in1), .out(andOp_156_out));

	reg [0:0] notOp_157_in0;
	wire [0:0] notOp_157_out;
	notOp #(.WIDTH(1)) notOp_157(.in(notOp_157_in0), .out(notOp_157_out));

	reg [0:0] andOp_158_in0;
	reg [0:0] andOp_158_in1;
	wire [0:0] andOp_158_out;
	andOp #(.WIDTH(1)) andOp_158(.in0(andOp_158_in0), .in1(andOp_158_in1), .out(andOp_158_out));

	reg [31:0] eq_159_in0;
	reg [31:0] eq_159_in1;
	wire [0:0] eq_159_out;
	eq #(.WIDTH(32)) eq_159(.in0(eq_159_in0), .in1(eq_159_in1), .out(eq_159_out));

	reg [0:0] andOp_160_in0;
	reg [0:0] andOp_160_in1;
	wire [0:0] andOp_160_out;
	andOp #(.WIDTH(1)) andOp_160(.in0(andOp_160_in0), .in1(andOp_160_in1), .out(andOp_160_out));

	reg [31:0] eq_161_in0;
	reg [31:0] eq_161_in1;
	wire [0:0] eq_161_out;
	eq #(.WIDTH(32)) eq_161(.in0(eq_161_in0), .in1(eq_161_in1), .out(eq_161_out));

	reg [0:0] andOp_162_in0;
	reg [0:0] andOp_162_in1;
	wire [0:0] andOp_162_out;
	andOp #(.WIDTH(1)) andOp_162(.in0(andOp_162_in0), .in1(andOp_162_in1), .out(andOp_162_out));

	reg [0:0] notOp_163_in0;
	wire [0:0] notOp_163_out;
	notOp #(.WIDTH(1)) notOp_163(.in(notOp_163_in0), .out(notOp_163_out));

	reg [0:0] andOp_164_in0;
	reg [0:0] andOp_164_in1;
	wire [0:0] andOp_164_out;
	andOp #(.WIDTH(1)) andOp_164(.in0(andOp_164_in0), .in1(andOp_164_in1), .out(andOp_164_out));

	reg [31:0] eq_165_in0;
	reg [31:0] eq_165_in1;
	wire [0:0] eq_165_out;
	eq #(.WIDTH(32)) eq_165(.in0(eq_165_in0), .in1(eq_165_in1), .out(eq_165_out));

	reg [0:0] andOp_166_in0;
	reg [0:0] andOp_166_in1;
	wire [0:0] andOp_166_out;
	andOp #(.WIDTH(1)) andOp_166(.in0(andOp_166_in0), .in1(andOp_166_in1), .out(andOp_166_out));

	reg [0:0] notOp_167_in0;
	wire [0:0] notOp_167_out;
	notOp #(.WIDTH(1)) notOp_167(.in(notOp_167_in0), .out(notOp_167_out));

	reg [0:0] andOp_168_in0;
	reg [0:0] andOp_168_in1;
	wire [0:0] andOp_168_out;
	andOp #(.WIDTH(1)) andOp_168(.in0(andOp_168_in0), .in1(andOp_168_in1), .out(andOp_168_out));

	reg [31:0] eq_169_in0;
	reg [31:0] eq_169_in1;
	wire [0:0] eq_169_out;
	eq #(.WIDTH(32)) eq_169(.in0(eq_169_in0), .in1(eq_169_in1), .out(eq_169_out));

	reg [0:0] andOp_170_in0;
	reg [0:0] andOp_170_in1;
	wire [0:0] andOp_170_out;
	andOp #(.WIDTH(1)) andOp_170(.in0(andOp_170_in0), .in1(andOp_170_in1), .out(andOp_170_out));

	reg [31:0] eq_171_in0;
	reg [31:0] eq_171_in1;
	wire [0:0] eq_171_out;
	eq #(.WIDTH(32)) eq_171(.in0(eq_171_in0), .in1(eq_171_in1), .out(eq_171_out));

	reg [0:0] andOp_172_in0;
	reg [0:0] andOp_172_in1;
	wire [0:0] andOp_172_out;
	andOp #(.WIDTH(1)) andOp_172(.in0(andOp_172_in0), .in1(andOp_172_in1), .out(andOp_172_out));

	reg [0:0] notOp_173_in0;
	wire [0:0] notOp_173_out;
	notOp #(.WIDTH(1)) notOp_173(.in(notOp_173_in0), .out(notOp_173_out));

	reg [0:0] andOp_174_in0;
	reg [0:0] andOp_174_in1;
	wire [0:0] andOp_174_out;
	andOp #(.WIDTH(1)) andOp_174(.in0(andOp_174_in0), .in1(andOp_174_in1), .out(andOp_174_out));

	reg [31:0] eq_175_in0;
	reg [31:0] eq_175_in1;
	wire [0:0] eq_175_out;
	eq #(.WIDTH(32)) eq_175(.in0(eq_175_in0), .in1(eq_175_in1), .out(eq_175_out));

	reg [0:0] andOp_176_in0;
	reg [0:0] andOp_176_in1;
	wire [0:0] andOp_176_out;
	andOp #(.WIDTH(1)) andOp_176(.in0(andOp_176_in0), .in1(andOp_176_in1), .out(andOp_176_out));

	reg [31:0] eq_177_in0;
	reg [31:0] eq_177_in1;
	wire [0:0] eq_177_out;
	eq #(.WIDTH(32)) eq_177(.in0(eq_177_in0), .in1(eq_177_in1), .out(eq_177_out));

	reg [0:0] andOp_178_in0;
	reg [0:0] andOp_178_in1;
	wire [0:0] andOp_178_out;
	andOp #(.WIDTH(1)) andOp_178(.in0(andOp_178_in0), .in1(andOp_178_in1), .out(andOp_178_out));

	reg [0:0] notOp_179_in0;
	wire [0:0] notOp_179_out;
	notOp #(.WIDTH(1)) notOp_179(.in(notOp_179_in0), .out(notOp_179_out));

	reg [0:0] andOp_180_in0;
	reg [0:0] andOp_180_in1;
	wire [0:0] andOp_180_out;
	andOp #(.WIDTH(1)) andOp_180(.in0(andOp_180_in0), .in1(andOp_180_in1), .out(andOp_180_out));

	reg [31:0] eq_181_in0;
	reg [31:0] eq_181_in1;
	wire [0:0] eq_181_out;
	eq #(.WIDTH(32)) eq_181(.in0(eq_181_in0), .in1(eq_181_in1), .out(eq_181_out));

	reg [0:0] andOp_182_in0;
	reg [0:0] andOp_182_in1;
	wire [0:0] andOp_182_out;
	andOp #(.WIDTH(1)) andOp_182(.in0(andOp_182_in0), .in1(andOp_182_in1), .out(andOp_182_out));

	reg [31:0] eq_183_in0;
	reg [31:0] eq_183_in1;
	wire [0:0] eq_183_out;
	eq #(.WIDTH(32)) eq_183(.in0(eq_183_in0), .in1(eq_183_in1), .out(eq_183_out));

	reg [0:0] andOp_184_in0;
	reg [0:0] andOp_184_in1;
	wire [0:0] andOp_184_out;
	andOp #(.WIDTH(1)) andOp_184(.in0(andOp_184_in0), .in1(andOp_184_in1), .out(andOp_184_out));

	reg [0:0] notOp_185_in0;
	wire [0:0] notOp_185_out;
	notOp #(.WIDTH(1)) notOp_185(.in(notOp_185_in0), .out(notOp_185_out));

	reg [0:0] andOp_186_in0;
	reg [0:0] andOp_186_in1;
	wire [0:0] andOp_186_out;
	andOp #(.WIDTH(1)) andOp_186(.in0(andOp_186_in0), .in1(andOp_186_in1), .out(andOp_186_out));

	reg [31:0] eq_187_in0;
	reg [31:0] eq_187_in1;
	wire [0:0] eq_187_out;
	eq #(.WIDTH(32)) eq_187(.in0(eq_187_in0), .in1(eq_187_in1), .out(eq_187_out));

	reg [0:0] andOp_188_in0;
	reg [0:0] andOp_188_in1;
	wire [0:0] andOp_188_out;
	andOp #(.WIDTH(1)) andOp_188(.in0(andOp_188_in0), .in1(andOp_188_in1), .out(andOp_188_out));

	reg [31:0] eq_189_in0;
	reg [31:0] eq_189_in1;
	wire [0:0] eq_189_out;
	eq #(.WIDTH(32)) eq_189(.in0(eq_189_in0), .in1(eq_189_in1), .out(eq_189_out));

	reg [0:0] andOp_190_in0;
	reg [0:0] andOp_190_in1;
	wire [0:0] andOp_190_out;
	andOp #(.WIDTH(1)) andOp_190(.in0(andOp_190_in0), .in1(andOp_190_in1), .out(andOp_190_out));

	reg [0:0] notOp_191_in0;
	wire [0:0] notOp_191_out;
	notOp #(.WIDTH(1)) notOp_191(.in(notOp_191_in0), .out(notOp_191_out));

	reg [0:0] andOp_192_in0;
	reg [0:0] andOp_192_in1;
	wire [0:0] andOp_192_out;
	andOp #(.WIDTH(1)) andOp_192(.in0(andOp_192_in0), .in1(andOp_192_in1), .out(andOp_192_out));

	reg [31:0] eq_193_in0;
	reg [31:0] eq_193_in1;
	wire [0:0] eq_193_out;
	eq #(.WIDTH(32)) eq_193(.in0(eq_193_in0), .in1(eq_193_in1), .out(eq_193_out));

	reg [0:0] andOp_194_in0;
	reg [0:0] andOp_194_in1;
	wire [0:0] andOp_194_out;
	andOp #(.WIDTH(1)) andOp_194(.in0(andOp_194_in0), .in1(andOp_194_in1), .out(andOp_194_out));

	reg [31:0] eq_195_in0;
	reg [31:0] eq_195_in1;
	wire [0:0] eq_195_out;
	eq #(.WIDTH(32)) eq_195(.in0(eq_195_in0), .in1(eq_195_in1), .out(eq_195_out));

	reg [0:0] andOp_196_in0;
	reg [0:0] andOp_196_in1;
	wire [0:0] andOp_196_out;
	andOp #(.WIDTH(1)) andOp_196(.in0(andOp_196_in0), .in1(andOp_196_in1), .out(andOp_196_out));

	reg [0:0] andOp_197_in0;
	reg [0:0] andOp_197_in1;
	wire [0:0] andOp_197_out;
	andOp #(.WIDTH(1)) andOp_197(.in0(andOp_197_in0), .in1(andOp_197_in1), .out(andOp_197_out));

	reg [31:0] eq_198_in0;
	reg [31:0] eq_198_in1;
	wire [0:0] eq_198_out;
	eq #(.WIDTH(32)) eq_198(.in0(eq_198_in0), .in1(eq_198_in1), .out(eq_198_out));

	reg [31:0] andOp_199_in0;
	reg [31:0] andOp_199_in1;
	wire [31:0] andOp_199_out;
	andOp #(.WIDTH(32)) andOp_199(.in0(andOp_199_in0), .in1(andOp_199_in1), .out(andOp_199_out));

	reg [31:0] eq_200_in0;
	reg [31:0] eq_200_in1;
	wire [0:0] eq_200_out;
	eq #(.WIDTH(32)) eq_200(.in0(eq_200_in0), .in1(eq_200_in1), .out(eq_200_out));

	reg [0:0] andOp_201_in0;
	reg [0:0] andOp_201_in1;
	wire [0:0] andOp_201_out;
	andOp #(.WIDTH(1)) andOp_201(.in0(andOp_201_in0), .in1(andOp_201_in1), .out(andOp_201_out));

	reg [0:0] andOp_202_in0;
	reg [0:0] andOp_202_in1;
	wire [0:0] andOp_202_out;
	andOp #(.WIDTH(1)) andOp_202(.in0(andOp_202_in0), .in1(andOp_202_in1), .out(andOp_202_out));

	reg [31:0] eq_203_in0;
	reg [31:0] eq_203_in1;
	wire [0:0] eq_203_out;
	eq #(.WIDTH(32)) eq_203(.in0(eq_203_in0), .in1(eq_203_in1), .out(eq_203_out));

	reg [31:0] andOp_204_in0;
	reg [31:0] andOp_204_in1;
	wire [31:0] andOp_204_out;
	andOp #(.WIDTH(32)) andOp_204(.in0(andOp_204_in0), .in1(andOp_204_in1), .out(andOp_204_out));

	reg [31:0] eq_205_in0;
	reg [31:0] eq_205_in1;
	wire [0:0] eq_205_out;
	eq #(.WIDTH(32)) eq_205(.in0(eq_205_in0), .in1(eq_205_in1), .out(eq_205_out));

	reg [0:0] andOp_206_in0;
	reg [0:0] andOp_206_in1;
	wire [0:0] andOp_206_out;
	andOp #(.WIDTH(1)) andOp_206(.in0(andOp_206_in0), .in1(andOp_206_in1), .out(andOp_206_out));

	reg [0:0] andOp_207_in0;
	reg [0:0] andOp_207_in1;
	wire [0:0] andOp_207_out;
	andOp #(.WIDTH(1)) andOp_207(.in0(andOp_207_in0), .in1(andOp_207_in1), .out(andOp_207_out));

	reg [31:0] eq_208_in0;
	reg [31:0] eq_208_in1;
	wire [0:0] eq_208_out;
	eq #(.WIDTH(32)) eq_208(.in0(eq_208_in0), .in1(eq_208_in1), .out(eq_208_out));

	reg [31:0] andOp_209_in0;
	reg [31:0] andOp_209_in1;
	wire [31:0] andOp_209_out;
	andOp #(.WIDTH(32)) andOp_209(.in0(andOp_209_in0), .in1(andOp_209_in1), .out(andOp_209_out));

	reg [0:0] notOp_210_in0;
	wire [0:0] notOp_210_out;
	notOp #(.WIDTH(1)) notOp_210(.in(notOp_210_in0), .out(notOp_210_out));

	reg [31:0] eq_211_in0;
	reg [31:0] eq_211_in1;
	wire [0:0] eq_211_out;
	eq #(.WIDTH(32)) eq_211(.in0(eq_211_in0), .in1(eq_211_in1), .out(eq_211_out));

	reg [0:0] andOp_212_in0;
	reg [0:0] andOp_212_in1;
	wire [0:0] andOp_212_out;
	andOp #(.WIDTH(1)) andOp_212(.in0(andOp_212_in0), .in1(andOp_212_in1), .out(andOp_212_out));

	reg [0:0] andOp_213_in0;
	reg [0:0] andOp_213_in1;
	wire [0:0] andOp_213_out;
	andOp #(.WIDTH(1)) andOp_213(.in0(andOp_213_in0), .in1(andOp_213_in1), .out(andOp_213_out));

	reg [31:0] eq_214_in0;
	reg [31:0] eq_214_in1;
	wire [0:0] eq_214_out;
	eq #(.WIDTH(32)) eq_214(.in0(eq_214_in0), .in1(eq_214_in1), .out(eq_214_out));

	reg [31:0] andOp_215_in0;
	reg [31:0] andOp_215_in1;
	wire [31:0] andOp_215_out;
	andOp #(.WIDTH(32)) andOp_215(.in0(andOp_215_in0), .in1(andOp_215_in1), .out(andOp_215_out));

	reg [31:0] eq_216_in0;
	reg [31:0] eq_216_in1;
	wire [0:0] eq_216_out;
	eq #(.WIDTH(32)) eq_216(.in0(eq_216_in0), .in1(eq_216_in1), .out(eq_216_out));

	reg [0:0] andOp_217_in0;
	reg [0:0] andOp_217_in1;
	wire [0:0] andOp_217_out;
	andOp #(.WIDTH(1)) andOp_217(.in0(andOp_217_in0), .in1(andOp_217_in1), .out(andOp_217_out));

	reg [0:0] andOp_218_in0;
	reg [0:0] andOp_218_in1;
	wire [0:0] andOp_218_out;
	andOp #(.WIDTH(1)) andOp_218(.in0(andOp_218_in0), .in1(andOp_218_in1), .out(andOp_218_out));

	reg [31:0] eq_219_in0;
	reg [31:0] eq_219_in1;
	wire [0:0] eq_219_out;
	eq #(.WIDTH(32)) eq_219(.in0(eq_219_in0), .in1(eq_219_in1), .out(eq_219_out));

	reg [31:0] andOp_220_in0;
	reg [31:0] andOp_220_in1;
	wire [31:0] andOp_220_out;
	andOp #(.WIDTH(32)) andOp_220(.in0(andOp_220_in0), .in1(andOp_220_in1), .out(andOp_220_out));

	reg [31:0] eq_221_in0;
	reg [31:0] eq_221_in1;
	wire [0:0] eq_221_out;
	eq #(.WIDTH(32)) eq_221(.in0(eq_221_in0), .in1(eq_221_in1), .out(eq_221_out));

	reg [0:0] andOp_222_in0;
	reg [0:0] andOp_222_in1;
	wire [0:0] andOp_222_out;
	andOp #(.WIDTH(1)) andOp_222(.in0(andOp_222_in0), .in1(andOp_222_in1), .out(andOp_222_out));

	reg [0:0] andOp_223_in0;
	reg [0:0] andOp_223_in1;
	wire [0:0] andOp_223_out;
	andOp #(.WIDTH(1)) andOp_223(.in0(andOp_223_in0), .in1(andOp_223_in1), .out(andOp_223_out));

	reg [31:0] eq_224_in0;
	reg [31:0] eq_224_in1;
	wire [0:0] eq_224_out;
	eq #(.WIDTH(32)) eq_224(.in0(eq_224_in0), .in1(eq_224_in1), .out(eq_224_out));

	reg [31:0] andOp_225_in0;
	reg [31:0] andOp_225_in1;
	wire [31:0] andOp_225_out;
	andOp #(.WIDTH(32)) andOp_225(.in0(andOp_225_in0), .in1(andOp_225_in1), .out(andOp_225_out));

	reg [31:0] eq_226_in0;
	reg [31:0] eq_226_in1;
	wire [0:0] eq_226_out;
	eq #(.WIDTH(32)) eq_226(.in0(eq_226_in0), .in1(eq_226_in1), .out(eq_226_out));

	reg [0:0] andOp_227_in0;
	reg [0:0] andOp_227_in1;
	wire [0:0] andOp_227_out;
	andOp #(.WIDTH(1)) andOp_227(.in0(andOp_227_in0), .in1(andOp_227_in1), .out(andOp_227_out));

	reg [0:0] andOp_228_in0;
	reg [0:0] andOp_228_in1;
	wire [0:0] andOp_228_out;
	andOp #(.WIDTH(1)) andOp_228(.in0(andOp_228_in0), .in1(andOp_228_in1), .out(andOp_228_out));

	reg [31:0] eq_229_in0;
	reg [31:0] eq_229_in1;
	wire [0:0] eq_229_out;
	eq #(.WIDTH(32)) eq_229(.in0(eq_229_in0), .in1(eq_229_in1), .out(eq_229_out));

	reg [31:0] andOp_230_in0;
	reg [31:0] andOp_230_in1;
	wire [31:0] andOp_230_out;
	andOp #(.WIDTH(32)) andOp_230(.in0(andOp_230_in0), .in1(andOp_230_in1), .out(andOp_230_out));

	reg [0:0] notOp_231_in0;
	wire [0:0] notOp_231_out;
	notOp #(.WIDTH(1)) notOp_231(.in(notOp_231_in0), .out(notOp_231_out));

	reg [31:0] eq_232_in0;
	reg [31:0] eq_232_in1;
	wire [0:0] eq_232_out;
	eq #(.WIDTH(32)) eq_232(.in0(eq_232_in0), .in1(eq_232_in1), .out(eq_232_out));

	reg [0:0] andOp_233_in0;
	reg [0:0] andOp_233_in1;
	wire [0:0] andOp_233_out;
	andOp #(.WIDTH(1)) andOp_233(.in0(andOp_233_in0), .in1(andOp_233_in1), .out(andOp_233_out));

	reg [0:0] andOp_234_in0;
	reg [0:0] andOp_234_in1;
	wire [0:0] andOp_234_out;
	andOp #(.WIDTH(1)) andOp_234(.in0(andOp_234_in0), .in1(andOp_234_in1), .out(andOp_234_out));

	reg [31:0] eq_235_in0;
	reg [31:0] eq_235_in1;
	wire [0:0] eq_235_out;
	eq #(.WIDTH(32)) eq_235(.in0(eq_235_in0), .in1(eq_235_in1), .out(eq_235_out));

	reg [31:0] andOp_236_in0;
	reg [31:0] andOp_236_in1;
	wire [31:0] andOp_236_out;
	andOp #(.WIDTH(32)) andOp_236(.in0(andOp_236_in0), .in1(andOp_236_in1), .out(andOp_236_out));

	reg [31:0] eq_237_in0;
	reg [31:0] eq_237_in1;
	wire [0:0] eq_237_out;
	eq #(.WIDTH(32)) eq_237(.in0(eq_237_in0), .in1(eq_237_in1), .out(eq_237_out));

	reg [0:0] andOp_238_in0;
	reg [0:0] andOp_238_in1;
	wire [0:0] andOp_238_out;
	andOp #(.WIDTH(1)) andOp_238(.in0(andOp_238_in0), .in1(andOp_238_in1), .out(andOp_238_out));

	reg [0:0] andOp_239_in0;
	reg [0:0] andOp_239_in1;
	wire [0:0] andOp_239_out;
	andOp #(.WIDTH(1)) andOp_239(.in0(andOp_239_in0), .in1(andOp_239_in1), .out(andOp_239_out));

	reg [31:0] eq_240_in0;
	reg [31:0] eq_240_in1;
	wire [0:0] eq_240_out;
	eq #(.WIDTH(32)) eq_240(.in0(eq_240_in0), .in1(eq_240_in1), .out(eq_240_out));

	reg [31:0] andOp_241_in0;
	reg [31:0] andOp_241_in1;
	wire [31:0] andOp_241_out;
	andOp #(.WIDTH(32)) andOp_241(.in0(andOp_241_in0), .in1(andOp_241_in1), .out(andOp_241_out));

	reg [31:0] eq_242_in0;
	reg [31:0] eq_242_in1;
	wire [0:0] eq_242_out;
	eq #(.WIDTH(32)) eq_242(.in0(eq_242_in0), .in1(eq_242_in1), .out(eq_242_out));

	reg [0:0] andOp_243_in0;
	reg [0:0] andOp_243_in1;
	wire [0:0] andOp_243_out;
	andOp #(.WIDTH(1)) andOp_243(.in0(andOp_243_in0), .in1(andOp_243_in1), .out(andOp_243_out));

	reg [0:0] andOp_244_in0;
	reg [0:0] andOp_244_in1;
	wire [0:0] andOp_244_out;
	andOp #(.WIDTH(1)) andOp_244(.in0(andOp_244_in0), .in1(andOp_244_in1), .out(andOp_244_out));

	reg [31:0] eq_245_in0;
	reg [31:0] eq_245_in1;
	wire [0:0] eq_245_out;
	eq #(.WIDTH(32)) eq_245(.in0(eq_245_in0), .in1(eq_245_in1), .out(eq_245_out));

	reg [31:0] andOp_246_in0;
	reg [31:0] andOp_246_in1;
	wire [31:0] andOp_246_out;
	andOp #(.WIDTH(32)) andOp_246(.in0(andOp_246_in0), .in1(andOp_246_in1), .out(andOp_246_out));

	reg [0:0] notOp_247_in0;
	wire [0:0] notOp_247_out;
	notOp #(.WIDTH(1)) notOp_247(.in(notOp_247_in0), .out(notOp_247_out));

	reg [31:0] eq_248_in0;
	reg [31:0] eq_248_in1;
	wire [0:0] eq_248_out;
	eq #(.WIDTH(32)) eq_248(.in0(eq_248_in0), .in1(eq_248_in1), .out(eq_248_out));

	reg [0:0] andOp_249_in0;
	reg [0:0] andOp_249_in1;
	wire [0:0] andOp_249_out;
	andOp #(.WIDTH(1)) andOp_249(.in0(andOp_249_in0), .in1(andOp_249_in1), .out(andOp_249_out));

	reg [0:0] andOp_250_in0;
	reg [0:0] andOp_250_in1;
	wire [0:0] andOp_250_out;
	andOp #(.WIDTH(1)) andOp_250(.in0(andOp_250_in0), .in1(andOp_250_in1), .out(andOp_250_out));

	reg [31:0] eq_251_in0;
	reg [31:0] eq_251_in1;
	wire [0:0] eq_251_out;
	eq #(.WIDTH(32)) eq_251(.in0(eq_251_in0), .in1(eq_251_in1), .out(eq_251_out));

	reg [31:0] andOp_252_in0;
	reg [31:0] andOp_252_in1;
	wire [31:0] andOp_252_out;
	andOp #(.WIDTH(32)) andOp_252(.in0(andOp_252_in0), .in1(andOp_252_in1), .out(andOp_252_out));

	reg [31:0] eq_253_in0;
	reg [31:0] eq_253_in1;
	wire [0:0] eq_253_out;
	eq #(.WIDTH(32)) eq_253(.in0(eq_253_in0), .in1(eq_253_in1), .out(eq_253_out));

	reg [0:0] andOp_254_in0;
	reg [0:0] andOp_254_in1;
	wire [0:0] andOp_254_out;
	andOp #(.WIDTH(1)) andOp_254(.in0(andOp_254_in0), .in1(andOp_254_in1), .out(andOp_254_out));

	reg [0:0] andOp_255_in0;
	reg [0:0] andOp_255_in1;
	wire [0:0] andOp_255_out;
	andOp #(.WIDTH(1)) andOp_255(.in0(andOp_255_in0), .in1(andOp_255_in1), .out(andOp_255_out));

	reg [31:0] eq_256_in0;
	reg [31:0] eq_256_in1;
	wire [0:0] eq_256_out;
	eq #(.WIDTH(32)) eq_256(.in0(eq_256_in0), .in1(eq_256_in1), .out(eq_256_out));

	reg [31:0] andOp_257_in0;
	reg [31:0] andOp_257_in1;
	wire [31:0] andOp_257_out;
	andOp #(.WIDTH(32)) andOp_257(.in0(andOp_257_in0), .in1(andOp_257_in1), .out(andOp_257_out));

	reg [31:0] eq_258_in0;
	reg [31:0] eq_258_in1;
	wire [0:0] eq_258_out;
	eq #(.WIDTH(32)) eq_258(.in0(eq_258_in0), .in1(eq_258_in1), .out(eq_258_out));

	reg [0:0] andOp_259_in0;
	reg [0:0] andOp_259_in1;
	wire [0:0] andOp_259_out;
	andOp #(.WIDTH(1)) andOp_259(.in0(andOp_259_in0), .in1(andOp_259_in1), .out(andOp_259_out));

	reg [0:0] andOp_260_in0;
	reg [0:0] andOp_260_in1;
	wire [0:0] andOp_260_out;
	andOp #(.WIDTH(1)) andOp_260(.in0(andOp_260_in0), .in1(andOp_260_in1), .out(andOp_260_out));

	reg [31:0] eq_261_in0;
	reg [31:0] eq_261_in1;
	wire [0:0] eq_261_out;
	eq #(.WIDTH(32)) eq_261(.in0(eq_261_in0), .in1(eq_261_in1), .out(eq_261_out));

	reg [31:0] andOp_262_in0;
	reg [31:0] andOp_262_in1;
	wire [31:0] andOp_262_out;
	andOp #(.WIDTH(32)) andOp_262(.in0(andOp_262_in0), .in1(andOp_262_in1), .out(andOp_262_out));

	reg [31:0] eq_263_in0;
	reg [31:0] eq_263_in1;
	wire [0:0] eq_263_out;
	eq #(.WIDTH(32)) eq_263(.in0(eq_263_in0), .in1(eq_263_in1), .out(eq_263_out));

	reg [0:0] andOp_264_in0;
	reg [0:0] andOp_264_in1;
	wire [0:0] andOp_264_out;
	andOp #(.WIDTH(1)) andOp_264(.in0(andOp_264_in0), .in1(andOp_264_in1), .out(andOp_264_out));

	reg [31:0] eq_265_in0;
	reg [31:0] eq_265_in1;
	wire [0:0] eq_265_out;
	eq #(.WIDTH(32)) eq_265(.in0(eq_265_in0), .in1(eq_265_in1), .out(eq_265_out));

	reg [0:0] andOp_266_in0;
	reg [0:0] andOp_266_in1;
	wire [0:0] andOp_266_out;
	andOp #(.WIDTH(1)) andOp_266(.in0(andOp_266_in0), .in1(andOp_266_in1), .out(andOp_266_out));

	reg [31:0] eq_267_in0;
	reg [31:0] eq_267_in1;
	wire [0:0] eq_267_out;
	eq #(.WIDTH(32)) eq_267(.in0(eq_267_in0), .in1(eq_267_in1), .out(eq_267_out));

	reg [0:0] andOp_268_in0;
	reg [0:0] andOp_268_in1;
	wire [0:0] andOp_268_out;
	andOp #(.WIDTH(1)) andOp_268(.in0(andOp_268_in0), .in1(andOp_268_in1), .out(andOp_268_out));

	reg [31:0] eq_269_in0;
	reg [31:0] eq_269_in1;
	wire [0:0] eq_269_out;
	eq #(.WIDTH(32)) eq_269(.in0(eq_269_in0), .in1(eq_269_in1), .out(eq_269_out));

	reg [0:0] andOp_270_in0;
	reg [0:0] andOp_270_in1;
	wire [0:0] andOp_270_out;
	andOp #(.WIDTH(1)) andOp_270(.in0(andOp_270_in0), .in1(andOp_270_in1), .out(andOp_270_out));

	reg [31:0] eq_271_in0;
	reg [31:0] eq_271_in1;
	wire [0:0] eq_271_out;
	eq #(.WIDTH(32)) eq_271(.in0(eq_271_in0), .in1(eq_271_in1), .out(eq_271_out));

	reg [0:0] andOp_272_in0;
	reg [0:0] andOp_272_in1;
	wire [0:0] andOp_272_out;
	andOp #(.WIDTH(1)) andOp_272(.in0(andOp_272_in0), .in1(andOp_272_in1), .out(andOp_272_out));

	reg [31:0] eq_273_in0;
	reg [31:0] eq_273_in1;
	wire [0:0] eq_273_out;
	eq #(.WIDTH(32)) eq_273(.in0(eq_273_in0), .in1(eq_273_in1), .out(eq_273_out));

	reg [0:0] andOp_274_in0;
	reg [0:0] andOp_274_in1;
	wire [0:0] andOp_274_out;
	andOp #(.WIDTH(1)) andOp_274(.in0(andOp_274_in0), .in1(andOp_274_in1), .out(andOp_274_out));

	reg [31:0] eq_275_in0;
	reg [31:0] eq_275_in1;
	wire [0:0] eq_275_out;
	eq #(.WIDTH(32)) eq_275(.in0(eq_275_in0), .in1(eq_275_in1), .out(eq_275_out));

	reg [0:0] andOp_276_in0;
	reg [0:0] andOp_276_in1;
	wire [0:0] andOp_276_out;
	andOp #(.WIDTH(1)) andOp_276(.in0(andOp_276_in0), .in1(andOp_276_in1), .out(andOp_276_out));

	reg [31:0] andOp_277_in0;
	reg [31:0] andOp_277_in1;
	wire [31:0] andOp_277_out;
	andOp #(.WIDTH(32)) andOp_277(.in0(andOp_277_in0), .in1(andOp_277_in1), .out(andOp_277_out));

	reg [31:0] eq_278_in0;
	reg [31:0] eq_278_in1;
	wire [0:0] eq_278_out;
	eq #(.WIDTH(32)) eq_278(.in0(eq_278_in0), .in1(eq_278_in1), .out(eq_278_out));

	reg [0:0] andOp_279_in0;
	reg [0:0] andOp_279_in1;
	wire [0:0] andOp_279_out;
	andOp #(.WIDTH(1)) andOp_279(.in0(andOp_279_in0), .in1(andOp_279_in1), .out(andOp_279_out));

	reg [31:0] eq_280_in0;
	reg [31:0] eq_280_in1;
	wire [0:0] eq_280_out;
	eq #(.WIDTH(32)) eq_280(.in0(eq_280_in0), .in1(eq_280_in1), .out(eq_280_out));

	reg [0:0] andOp_281_in0;
	reg [0:0] andOp_281_in1;
	wire [0:0] andOp_281_out;
	andOp #(.WIDTH(1)) andOp_281(.in0(andOp_281_in0), .in1(andOp_281_in1), .out(andOp_281_out));

	reg [31:0] eq_282_in0;
	reg [31:0] eq_282_in1;
	wire [0:0] eq_282_out;
	eq #(.WIDTH(32)) eq_282(.in0(eq_282_in0), .in1(eq_282_in1), .out(eq_282_out));

	reg [0:0] andOp_283_in0;
	reg [0:0] andOp_283_in1;
	wire [0:0] andOp_283_out;
	andOp #(.WIDTH(1)) andOp_283(.in0(andOp_283_in0), .in1(andOp_283_in1), .out(andOp_283_out));

	reg [31:0] eq_284_in0;
	reg [31:0] eq_284_in1;
	wire [0:0] eq_284_out;
	eq #(.WIDTH(32)) eq_284(.in0(eq_284_in0), .in1(eq_284_in1), .out(eq_284_out));

	reg [0:0] andOp_285_in0;
	reg [0:0] andOp_285_in1;
	wire [0:0] andOp_285_out;
	andOp #(.WIDTH(1)) andOp_285(.in0(andOp_285_in0), .in1(andOp_285_in1), .out(andOp_285_out));

	reg [31:0] eq_286_in0;
	reg [31:0] eq_286_in1;
	wire [0:0] eq_286_out;
	eq #(.WIDTH(32)) eq_286(.in0(eq_286_in0), .in1(eq_286_in1), .out(eq_286_out));

	reg [0:0] andOp_287_in0;
	reg [0:0] andOp_287_in1;
	wire [0:0] andOp_287_out;
	andOp #(.WIDTH(1)) andOp_287(.in0(andOp_287_in0), .in1(andOp_287_in1), .out(andOp_287_out));

	reg [31:0] eq_288_in0;
	reg [31:0] eq_288_in1;
	wire [0:0] eq_288_out;
	eq #(.WIDTH(32)) eq_288(.in0(eq_288_in0), .in1(eq_288_in1), .out(eq_288_out));

	reg [0:0] andOp_289_in0;
	reg [0:0] andOp_289_in1;
	wire [0:0] andOp_289_out;
	andOp #(.WIDTH(1)) andOp_289(.in0(andOp_289_in0), .in1(andOp_289_in1), .out(andOp_289_out));

	reg [31:0] eq_290_in0;
	reg [31:0] eq_290_in1;
	wire [0:0] eq_290_out;
	eq #(.WIDTH(32)) eq_290(.in0(eq_290_in0), .in1(eq_290_in1), .out(eq_290_out));

	reg [0:0] andOp_291_in0;
	reg [0:0] andOp_291_in1;
	wire [0:0] andOp_291_out;
	andOp #(.WIDTH(1)) andOp_291(.in0(andOp_291_in0), .in1(andOp_291_in1), .out(andOp_291_out));

	reg [31:0] eq_292_in0;
	reg [31:0] eq_292_in1;
	wire [0:0] eq_292_out;
	eq #(.WIDTH(32)) eq_292(.in0(eq_292_in0), .in1(eq_292_in1), .out(eq_292_out));

	reg [0:0] andOp_293_in0;
	reg [0:0] andOp_293_in1;
	wire [0:0] andOp_293_out;
	andOp #(.WIDTH(1)) andOp_293(.in0(andOp_293_in0), .in1(andOp_293_in1), .out(andOp_293_out));

	reg [31:0] andOp_294_in0;
	reg [31:0] andOp_294_in1;
	wire [31:0] andOp_294_out;
	andOp #(.WIDTH(32)) andOp_294(.in0(andOp_294_in0), .in1(andOp_294_in1), .out(andOp_294_out));

	reg [31:0] eq_295_in0;
	reg [31:0] eq_295_in1;
	wire [0:0] eq_295_out;
	eq #(.WIDTH(32)) eq_295(.in0(eq_295_in0), .in1(eq_295_in1), .out(eq_295_out));

	reg [0:0] andOp_296_in0;
	reg [0:0] andOp_296_in1;
	wire [0:0] andOp_296_out;
	andOp #(.WIDTH(1)) andOp_296(.in0(andOp_296_in0), .in1(andOp_296_in1), .out(andOp_296_out));

	reg [31:0] eq_297_in0;
	reg [31:0] eq_297_in1;
	wire [0:0] eq_297_out;
	eq #(.WIDTH(32)) eq_297(.in0(eq_297_in0), .in1(eq_297_in1), .out(eq_297_out));

	reg [0:0] andOp_298_in0;
	reg [0:0] andOp_298_in1;
	wire [0:0] andOp_298_out;
	andOp #(.WIDTH(1)) andOp_298(.in0(andOp_298_in0), .in1(andOp_298_in1), .out(andOp_298_out));

	reg [31:0] eq_299_in0;
	reg [31:0] eq_299_in1;
	wire [0:0] eq_299_out;
	eq #(.WIDTH(32)) eq_299(.in0(eq_299_in0), .in1(eq_299_in1), .out(eq_299_out));

	reg [0:0] andOp_300_in0;
	reg [0:0] andOp_300_in1;
	wire [0:0] andOp_300_out;
	andOp #(.WIDTH(1)) andOp_300(.in0(andOp_300_in0), .in1(andOp_300_in1), .out(andOp_300_out));

	reg [31:0] eq_301_in0;
	reg [31:0] eq_301_in1;
	wire [0:0] eq_301_out;
	eq #(.WIDTH(32)) eq_301(.in0(eq_301_in0), .in1(eq_301_in1), .out(eq_301_out));

	reg [0:0] andOp_302_in0;
	reg [0:0] andOp_302_in1;
	wire [0:0] andOp_302_out;
	andOp #(.WIDTH(1)) andOp_302(.in0(andOp_302_in0), .in1(andOp_302_in1), .out(andOp_302_out));

	reg [31:0] andOp_303_in0;
	reg [31:0] andOp_303_in1;
	wire [31:0] andOp_303_out;
	andOp #(.WIDTH(32)) andOp_303(.in0(andOp_303_in0), .in1(andOp_303_in1), .out(andOp_303_out));

	reg [31:0] eq_304_in0;
	reg [31:0] eq_304_in1;
	wire [0:0] eq_304_out;
	eq #(.WIDTH(32)) eq_304(.in0(eq_304_in0), .in1(eq_304_in1), .out(eq_304_out));

	reg [0:0] andOp_305_in0;
	reg [0:0] andOp_305_in1;
	wire [0:0] andOp_305_out;
	andOp #(.WIDTH(1)) andOp_305(.in0(andOp_305_in0), .in1(andOp_305_in1), .out(andOp_305_out));

	reg [31:0] eq_306_in0;
	reg [31:0] eq_306_in1;
	wire [0:0] eq_306_out;
	eq #(.WIDTH(32)) eq_306(.in0(eq_306_in0), .in1(eq_306_in1), .out(eq_306_out));

	reg [0:0] andOp_307_in0;
	reg [0:0] andOp_307_in1;
	wire [0:0] andOp_307_out;
	andOp #(.WIDTH(1)) andOp_307(.in0(andOp_307_in0), .in1(andOp_307_in1), .out(andOp_307_out));

	reg [31:0] andOp_308_in0;
	reg [31:0] andOp_308_in1;
	wire [31:0] andOp_308_out;
	andOp #(.WIDTH(32)) andOp_308(.in0(andOp_308_in0), .in1(andOp_308_in1), .out(andOp_308_out));

	reg [31:0] eq_309_in0;
	reg [31:0] eq_309_in1;
	wire [0:0] eq_309_out;
	eq #(.WIDTH(32)) eq_309(.in0(eq_309_in0), .in1(eq_309_in1), .out(eq_309_out));

	reg [0:0] andOp_310_in0;
	reg [0:0] andOp_310_in1;
	wire [0:0] andOp_310_out;
	andOp #(.WIDTH(1)) andOp_310(.in0(andOp_310_in0), .in1(andOp_310_in1), .out(andOp_310_out));

	reg [31:0] eq_311_in0;
	reg [31:0] eq_311_in1;
	wire [0:0] eq_311_out;
	eq #(.WIDTH(32)) eq_311(.in0(eq_311_in0), .in1(eq_311_in1), .out(eq_311_out));

	reg [0:0] andOp_312_in0;
	reg [0:0] andOp_312_in1;
	wire [0:0] andOp_312_out;
	andOp #(.WIDTH(1)) andOp_312(.in0(andOp_312_in0), .in1(andOp_312_in1), .out(andOp_312_out));

	reg [31:0] eq_313_in0;
	reg [31:0] eq_313_in1;
	wire [0:0] eq_313_out;
	eq #(.WIDTH(32)) eq_313(.in0(eq_313_in0), .in1(eq_313_in1), .out(eq_313_out));

	reg [0:0] andOp_314_in0;
	reg [0:0] andOp_314_in1;
	wire [0:0] andOp_314_out;
	andOp #(.WIDTH(1)) andOp_314(.in0(andOp_314_in0), .in1(andOp_314_in1), .out(andOp_314_out));

	reg [31:0] eq_315_in0;
	reg [31:0] eq_315_in1;
	wire [0:0] eq_315_out;
	eq #(.WIDTH(32)) eq_315(.in0(eq_315_in0), .in1(eq_315_in1), .out(eq_315_out));

	reg [0:0] andOp_316_in0;
	reg [0:0] andOp_316_in1;
	wire [0:0] andOp_316_out;
	andOp #(.WIDTH(1)) andOp_316(.in0(andOp_316_in0), .in1(andOp_316_in1), .out(andOp_316_out));

	reg [31:0] eq_317_in0;
	reg [31:0] eq_317_in1;
	wire [0:0] eq_317_out;
	eq #(.WIDTH(32)) eq_317(.in0(eq_317_in0), .in1(eq_317_in1), .out(eq_317_out));

	reg [0:0] andOp_318_in0;
	reg [0:0] andOp_318_in1;
	wire [0:0] andOp_318_out;
	andOp #(.WIDTH(1)) andOp_318(.in0(andOp_318_in0), .in1(andOp_318_in1), .out(andOp_318_out));

	reg [31:0] eq_319_in0;
	reg [31:0] eq_319_in1;
	wire [0:0] eq_319_out;
	eq #(.WIDTH(32)) eq_319(.in0(eq_319_in0), .in1(eq_319_in1), .out(eq_319_out));

	reg [0:0] andOp_320_in0;
	reg [0:0] andOp_320_in1;
	wire [0:0] andOp_320_out;
	andOp #(.WIDTH(1)) andOp_320(.in0(andOp_320_in0), .in1(andOp_320_in1), .out(andOp_320_out));

	reg [31:0] eq_321_in0;
	reg [31:0] eq_321_in1;
	wire [0:0] eq_321_out;
	eq #(.WIDTH(32)) eq_321(.in0(eq_321_in0), .in1(eq_321_in1), .out(eq_321_out));

	reg [0:0] andOp_322_in0;
	reg [0:0] andOp_322_in1;
	wire [0:0] andOp_322_out;
	andOp #(.WIDTH(1)) andOp_322(.in0(andOp_322_in0), .in1(andOp_322_in1), .out(andOp_322_out));

	reg [31:0] eq_323_in0;
	reg [31:0] eq_323_in1;
	wire [0:0] eq_323_out;
	eq #(.WIDTH(32)) eq_323(.in0(eq_323_in0), .in1(eq_323_in1), .out(eq_323_out));

	reg [0:0] andOp_324_in0;
	reg [0:0] andOp_324_in1;
	wire [0:0] andOp_324_out;
	andOp #(.WIDTH(1)) andOp_324(.in0(andOp_324_in0), .in1(andOp_324_in1), .out(andOp_324_out));

	reg [31:0] eq_325_in0;
	reg [31:0] eq_325_in1;
	wire [0:0] eq_325_out;
	eq #(.WIDTH(32)) eq_325(.in0(eq_325_in0), .in1(eq_325_in1), .out(eq_325_out));

	reg [0:0] andOp_326_in0;
	reg [0:0] andOp_326_in1;
	wire [0:0] andOp_326_out;
	andOp #(.WIDTH(1)) andOp_326(.in0(andOp_326_in0), .in1(andOp_326_in1), .out(andOp_326_out));

	reg [31:0] eq_327_in0;
	reg [31:0] eq_327_in1;
	wire [0:0] eq_327_out;
	eq #(.WIDTH(32)) eq_327(.in0(eq_327_in0), .in1(eq_327_in1), .out(eq_327_out));

	reg [0:0] andOp_328_in0;
	reg [0:0] andOp_328_in1;
	wire [0:0] andOp_328_out;
	andOp #(.WIDTH(1)) andOp_328(.in0(andOp_328_in0), .in1(andOp_328_in1), .out(andOp_328_out));

	reg [31:0] eq_329_in0;
	reg [31:0] eq_329_in1;
	wire [0:0] eq_329_out;
	eq #(.WIDTH(32)) eq_329(.in0(eq_329_in0), .in1(eq_329_in1), .out(eq_329_out));

	reg [0:0] andOp_330_in0;
	reg [0:0] andOp_330_in1;
	wire [0:0] andOp_330_out;
	andOp #(.WIDTH(1)) andOp_330(.in0(andOp_330_in0), .in1(andOp_330_in1), .out(andOp_330_out));

	reg [31:0] eq_331_in0;
	reg [31:0] eq_331_in1;
	wire [0:0] eq_331_out;
	eq #(.WIDTH(32)) eq_331(.in0(eq_331_in0), .in1(eq_331_in1), .out(eq_331_out));

	reg [0:0] andOp_332_in0;
	reg [0:0] andOp_332_in1;
	wire [0:0] andOp_332_out;
	andOp #(.WIDTH(1)) andOp_332(.in0(andOp_332_in0), .in1(andOp_332_in1), .out(andOp_332_out));

	// End Functional Units

	reg [31:0] add_tmp_5;
	reg [31:0] call_tmp_2;
	reg [31:0] global_next_block;
	reg [31:0] global_state;
	reg [0:0] icmp_tmp_6;
	reg [31:0] last_BB_reg;
	reg [31:0] phi_tmp_0;

	// controller for add_add_14.add_in0_add_14
	// controller for add_add_14.add_in1_add_14
	// Insensitive connections
	always @(*) begin
		add_in0_add_14 = valid ? rdata_ram_0 : rdata_ram_0;
		add_in1_add_14 = valid ? call_tmp_2 : call_tmp_2;
	end
	// controller for add_add_16.add_in0_add_16
	// controller for add_add_16.add_in1_add_16
	// Insensitive connections
	always @(*) begin
		add_in0_add_16 = valid ? phi_tmp_0 : phi_tmp_0;
		add_in1_add_16 = valid ? (32'd1) : (32'd1);
	end
	// controller for andOp_1.andOp_1_in0
	// controller for andOp_1.andOp_1_in1
	// Insensitive connections
	always @(*) begin
		andOp_1_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_1_in1 = valid ? eq_0_out : eq_0_out;
	end
	// controller for andOp_10.andOp_10_in0
	// controller for andOp_10.andOp_10_in1
	// Insensitive connections
	always @(*) begin
		andOp_10_in0 = valid ? andOp_9_out : andOp_9_out;
		andOp_10_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_100.andOp_100_in0
	// controller for andOp_100.andOp_100_in1
	// Insensitive connections
	always @(*) begin
		andOp_100_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_100_in1 = valid ? eq_99_out : eq_99_out;
	end
	// controller for andOp_102.andOp_102_in0
	// controller for andOp_102.andOp_102_in1
	// Insensitive connections
	always @(*) begin
		andOp_102_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_102_in1 = valid ? eq_101_out : eq_101_out;
	end
	// controller for andOp_104.andOp_104_in0
	// controller for andOp_104.andOp_104_in1
	// Insensitive connections
	always @(*) begin
		andOp_104_in0 = valid ? bb_7_active_out_data : bb_7_active_out_data;
		andOp_104_in1 = valid ? eq_103_out : eq_103_out;
	end
	// controller for andOp_106.andOp_106_in0
	// controller for andOp_106.andOp_106_in1
	// Insensitive connections
	always @(*) begin
		andOp_106_in0 = valid ? bb_3_active_out_data : bb_3_active_out_data;
		andOp_106_in1 = valid ? eq_105_out : eq_105_out;
	end
	// controller for andOp_108.andOp_108_in0
	// controller for andOp_108.andOp_108_in1
	// Insensitive connections
	always @(*) begin
		andOp_108_in0 = valid ? bb_9_active_out_data : bb_9_active_out_data;
		andOp_108_in1 = valid ? eq_107_out : eq_107_out;
	end
	// controller for andOp_110.andOp_110_in0
	// controller for andOp_110.andOp_110_in1
	// Insensitive connections
	always @(*) begin
		andOp_110_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_110_in1 = valid ? eq_109_out : eq_109_out;
	end
	// controller for andOp_112.andOp_112_in0
	// controller for andOp_112.andOp_112_in1
	// Insensitive connections
	always @(*) begin
		andOp_112_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_112_in1 = valid ? eq_111_out : eq_111_out;
	end
	// controller for andOp_114.andOp_114_in0
	// controller for andOp_114.andOp_114_in1
	// Insensitive connections
	always @(*) begin
		andOp_114_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_114_in1 = valid ? eq_113_out : eq_113_out;
	end
	// controller for andOp_116.andOp_116_in0
	// controller for andOp_116.andOp_116_in1
	// Insensitive connections
	always @(*) begin
		andOp_116_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_116_in1 = valid ? eq_115_out : eq_115_out;
	end
	// controller for andOp_118.andOp_118_in0
	// controller for andOp_118.andOp_118_in1
	// Insensitive connections
	always @(*) begin
		andOp_118_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_118_in1 = valid ? eq_117_out : eq_117_out;
	end
	// controller for andOp_120.andOp_120_in0
	// controller for andOp_120.andOp_120_in1
	// Insensitive connections
	always @(*) begin
		andOp_120_in0 = valid ? bb_6_active_out_data : bb_6_active_out_data;
		andOp_120_in1 = valid ? eq_119_out : eq_119_out;
	end
	// controller for andOp_122.andOp_122_in0
	// controller for andOp_122.andOp_122_in1
	// Insensitive connections
	always @(*) begin
		andOp_122_in0 = valid ? bb_7_active_out_data : bb_7_active_out_data;
		andOp_122_in1 = valid ? eq_121_out : eq_121_out;
	end
	// controller for andOp_124.andOp_124_in0
	// controller for andOp_124.andOp_124_in1
	// Insensitive connections
	always @(*) begin
		andOp_124_in0 = valid ? bb_7_active_out_data : bb_7_active_out_data;
		andOp_124_in1 = valid ? eq_123_out : eq_123_out;
	end
	// controller for andOp_126.andOp_126_in0
	// controller for andOp_126.andOp_126_in1
	// Insensitive connections
	always @(*) begin
		andOp_126_in0 = valid ? bb_2_active_out_data : bb_2_active_out_data;
		andOp_126_in1 = valid ? eq_125_out : eq_125_out;
	end
	// controller for andOp_128.andOp_128_in0
	// controller for andOp_128.andOp_128_in1
	// Insensitive connections
	always @(*) begin
		andOp_128_in0 = valid ? bb_2_active_out_data : bb_2_active_out_data;
		andOp_128_in1 = valid ? eq_127_out : eq_127_out;
	end
	// controller for andOp_13.andOp_13_in0
	// controller for andOp_13.andOp_13_in1
	// Insensitive connections
	always @(*) begin
		andOp_13_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_13_in1 = valid ? eq_12_out : eq_12_out;
	end
	// controller for andOp_130.andOp_130_in0
	// controller for andOp_130.andOp_130_in1
	// Insensitive connections
	always @(*) begin
		andOp_130_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_130_in1 = valid ? eq_129_out : eq_129_out;
	end
	// controller for andOp_132.andOp_132_in0
	// controller for andOp_132.andOp_132_in1
	// Insensitive connections
	always @(*) begin
		andOp_132_in0 = valid ? bb_3_active_out_data : bb_3_active_out_data;
		andOp_132_in1 = valid ? eq_131_out : eq_131_out;
	end
	// controller for andOp_134.andOp_134_in0
	// controller for andOp_134.andOp_134_in1
	// Insensitive connections
	always @(*) begin
		andOp_134_in0 = valid ? notOp_133_out : notOp_133_out;
		andOp_134_in1 = valid ? andOp_130_out : andOp_130_out;
	end
	// controller for andOp_136.andOp_136_in0
	// controller for andOp_136.andOp_136_in1
	// Insensitive connections
	always @(*) begin
		andOp_136_in0 = valid ? bb_3_active_out_data : bb_3_active_out_data;
		andOp_136_in1 = valid ? eq_135_out : eq_135_out;
	end
	// controller for andOp_138.andOp_138_in0
	// controller for andOp_138.andOp_138_in1
	// Insensitive connections
	always @(*) begin
		andOp_138_in0 = valid ? bb_8_active_out_data : bb_8_active_out_data;
		andOp_138_in1 = valid ? eq_137_out : eq_137_out;
	end
	// controller for andOp_14.andOp_14_in0
	// controller for andOp_14.andOp_14_in1
	// Insensitive connections
	always @(*) begin
		andOp_14_in0 = valid ? andOp_13_out : andOp_13_out;
		andOp_14_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_140.andOp_140_in0
	// controller for andOp_140.andOp_140_in1
	// Insensitive connections
	always @(*) begin
		andOp_140_in0 = valid ? notOp_139_out : notOp_139_out;
		andOp_140_in1 = valid ? andOp_136_out : andOp_136_out;
	end
	// controller for andOp_142.andOp_142_in0
	// controller for andOp_142.andOp_142_in1
	// Insensitive connections
	always @(*) begin
		andOp_142_in0 = valid ? bb_8_active_out_data : bb_8_active_out_data;
		andOp_142_in1 = valid ? eq_141_out : eq_141_out;
	end
	// controller for andOp_144.andOp_144_in0
	// controller for andOp_144.andOp_144_in1
	// Insensitive connections
	always @(*) begin
		andOp_144_in0 = valid ? bb_9_active_out_data : bb_9_active_out_data;
		andOp_144_in1 = valid ? eq_143_out : eq_143_out;
	end
	// controller for andOp_146.andOp_146_in0
	// controller for andOp_146.andOp_146_in1
	// Insensitive connections
	always @(*) begin
		andOp_146_in0 = valid ? notOp_145_out : notOp_145_out;
		andOp_146_in1 = valid ? andOp_142_out : andOp_142_out;
	end
	// controller for andOp_148.andOp_148_in0
	// controller for andOp_148.andOp_148_in1
	// Insensitive connections
	always @(*) begin
		andOp_148_in0 = valid ? bb_9_active_out_data : bb_9_active_out_data;
		andOp_148_in1 = valid ? eq_147_out : eq_147_out;
	end
	// controller for andOp_150.andOp_150_in0
	// controller for andOp_150.andOp_150_in1
	// Insensitive connections
	always @(*) begin
		andOp_150_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_150_in1 = valid ? eq_149_out : eq_149_out;
	end
	// controller for andOp_152.andOp_152_in0
	// controller for andOp_152.andOp_152_in1
	// Insensitive connections
	always @(*) begin
		andOp_152_in0 = valid ? notOp_151_out : notOp_151_out;
		andOp_152_in1 = valid ? andOp_148_out : andOp_148_out;
	end
	// controller for andOp_154.andOp_154_in0
	// controller for andOp_154.andOp_154_in1
	// Insensitive connections
	always @(*) begin
		andOp_154_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_154_in1 = valid ? eq_153_out : eq_153_out;
	end
	// controller for andOp_156.andOp_156_in0
	// controller for andOp_156.andOp_156_in1
	// Insensitive connections
	always @(*) begin
		andOp_156_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_156_in1 = valid ? eq_155_out : eq_155_out;
	end
	// controller for andOp_158.andOp_158_in0
	// controller for andOp_158.andOp_158_in1
	// Insensitive connections
	always @(*) begin
		andOp_158_in0 = valid ? notOp_157_out : notOp_157_out;
		andOp_158_in1 = valid ? andOp_154_out : andOp_154_out;
	end
	// controller for andOp_16.andOp_16_in0
	// controller for andOp_16.andOp_16_in1
	// Insensitive connections
	always @(*) begin
		andOp_16_in0 = valid ? andOp_14_out : andOp_14_out;
		andOp_16_in1 = valid ? icmp_tmp_6 : icmp_tmp_6;
	end
	// controller for andOp_160.andOp_160_in0
	// controller for andOp_160.andOp_160_in1
	// Insensitive connections
	always @(*) begin
		andOp_160_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_160_in1 = valid ? eq_159_out : eq_159_out;
	end
	// controller for andOp_162.andOp_162_in0
	// controller for andOp_162.andOp_162_in1
	// Insensitive connections
	always @(*) begin
		andOp_162_in0 = valid ? bb_1_active_out_data : bb_1_active_out_data;
		andOp_162_in1 = valid ? eq_161_out : eq_161_out;
	end
	// controller for andOp_164.andOp_164_in0
	// controller for andOp_164.andOp_164_in1
	// Insensitive connections
	always @(*) begin
		andOp_164_in0 = valid ? notOp_163_out : notOp_163_out;
		andOp_164_in1 = valid ? andOp_160_out : andOp_160_out;
	end
	// controller for andOp_166.andOp_166_in0
	// controller for andOp_166.andOp_166_in1
	// Insensitive connections
	always @(*) begin
		andOp_166_in0 = valid ? bb_3_active_out_data : bb_3_active_out_data;
		andOp_166_in1 = valid ? eq_165_out : eq_165_out;
	end
	// controller for andOp_168.andOp_168_in0
	// controller for andOp_168.andOp_168_in1
	// Insensitive connections
	always @(*) begin
		andOp_168_in0 = valid ? notOp_167_out : notOp_167_out;
		andOp_168_in1 = valid ? andOp_164_out : andOp_164_out;
	end
	// controller for andOp_170.andOp_170_in0
	// controller for andOp_170.andOp_170_in1
	// Insensitive connections
	always @(*) begin
		andOp_170_in0 = valid ? bb_1_active_out_data : bb_1_active_out_data;
		andOp_170_in1 = valid ? eq_169_out : eq_169_out;
	end
	// controller for andOp_172.andOp_172_in0
	// controller for andOp_172.andOp_172_in1
	// Insensitive connections
	always @(*) begin
		andOp_172_in0 = valid ? bb_5_active_out_data : bb_5_active_out_data;
		andOp_172_in1 = valid ? eq_171_out : eq_171_out;
	end
	// controller for andOp_174.andOp_174_in0
	// controller for andOp_174.andOp_174_in1
	// Insensitive connections
	always @(*) begin
		andOp_174_in0 = valid ? notOp_173_out : notOp_173_out;
		andOp_174_in1 = valid ? andOp_170_out : andOp_170_out;
	end
	// controller for andOp_176.andOp_176_in0
	// controller for andOp_176.andOp_176_in1
	// Insensitive connections
	always @(*) begin
		andOp_176_in0 = valid ? bb_5_active_out_data : bb_5_active_out_data;
		andOp_176_in1 = valid ? eq_175_out : eq_175_out;
	end
	// controller for andOp_178.andOp_178_in0
	// controller for andOp_178.andOp_178_in1
	// Insensitive connections
	always @(*) begin
		andOp_178_in0 = valid ? bb_6_active_out_data : bb_6_active_out_data;
		andOp_178_in1 = valid ? eq_177_out : eq_177_out;
	end
	// controller for andOp_18.andOp_18_in0
	// controller for andOp_18.andOp_18_in1
	// Insensitive connections
	always @(*) begin
		andOp_18_in0 = valid ? andOp_14_out : andOp_14_out;
		andOp_18_in1 = valid ? notOp_17_out : notOp_17_out;
	end
	// controller for andOp_180.andOp_180_in0
	// controller for andOp_180.andOp_180_in1
	// Insensitive connections
	always @(*) begin
		andOp_180_in0 = valid ? notOp_179_out : notOp_179_out;
		andOp_180_in1 = valid ? andOp_176_out : andOp_176_out;
	end
	// controller for andOp_182.andOp_182_in0
	// controller for andOp_182.andOp_182_in1
	// Insensitive connections
	always @(*) begin
		andOp_182_in0 = valid ? bb_6_active_out_data : bb_6_active_out_data;
		andOp_182_in1 = valid ? eq_181_out : eq_181_out;
	end
	// controller for andOp_184.andOp_184_in0
	// controller for andOp_184.andOp_184_in1
	// Insensitive connections
	always @(*) begin
		andOp_184_in0 = valid ? bb_7_active_out_data : bb_7_active_out_data;
		andOp_184_in1 = valid ? eq_183_out : eq_183_out;
	end
	// controller for andOp_186.andOp_186_in0
	// controller for andOp_186.andOp_186_in1
	// Insensitive connections
	always @(*) begin
		andOp_186_in0 = valid ? notOp_185_out : notOp_185_out;
		andOp_186_in1 = valid ? andOp_182_out : andOp_182_out;
	end
	// controller for andOp_188.andOp_188_in0
	// controller for andOp_188.andOp_188_in1
	// Insensitive connections
	always @(*) begin
		andOp_188_in0 = valid ? bb_7_active_out_data : bb_7_active_out_data;
		andOp_188_in1 = valid ? eq_187_out : eq_187_out;
	end
	// controller for andOp_190.andOp_190_in0
	// controller for andOp_190.andOp_190_in1
	// Insensitive connections
	always @(*) begin
		andOp_190_in0 = valid ? bb_2_active_out_data : bb_2_active_out_data;
		andOp_190_in1 = valid ? eq_189_out : eq_189_out;
	end
	// controller for andOp_192.andOp_192_in0
	// controller for andOp_192.andOp_192_in1
	// Insensitive connections
	always @(*) begin
		andOp_192_in0 = valid ? notOp_191_out : notOp_191_out;
		andOp_192_in1 = valid ? andOp_188_out : andOp_188_out;
	end
	// controller for andOp_194.andOp_194_in0
	// controller for andOp_194.andOp_194_in1
	// Insensitive connections
	always @(*) begin
		andOp_194_in0 = valid ? bb_2_active_out_data : bb_2_active_out_data;
		andOp_194_in1 = valid ? eq_193_out : eq_193_out;
	end
	// controller for andOp_196.andOp_196_in0
	// controller for andOp_196.andOp_196_in1
	// Insensitive connections
	always @(*) begin
		andOp_196_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_196_in1 = valid ? eq_195_out : eq_195_out;
	end
	// controller for andOp_197.andOp_197_in0
	// controller for andOp_197.andOp_197_in1
	// Insensitive connections
	always @(*) begin
		andOp_197_in0 = valid ? andOp_196_out : andOp_196_out;
		andOp_197_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_199.andOp_199_in0
	// controller for andOp_199.andOp_199_in1
	// Insensitive connections
	always @(*) begin
		andOp_199_in0 = valid ? eq_198_out : eq_198_out;
		andOp_199_in1 = valid ? andOp_197_out : andOp_197_out;
	end
	// controller for andOp_2.andOp_2_in0
	// controller for andOp_2.andOp_2_in1
	// Insensitive connections
	always @(*) begin
		andOp_2_in0 = valid ? andOp_1_out : andOp_1_out;
		andOp_2_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_20.andOp_20_in0
	// controller for andOp_20.andOp_20_in1
	// Insensitive connections
	always @(*) begin
		andOp_20_in0 = valid ? bb_5_active_out_data : bb_5_active_out_data;
		andOp_20_in1 = valid ? eq_19_out : eq_19_out;
	end
	// controller for andOp_201.andOp_201_in0
	// controller for andOp_201.andOp_201_in1
	// Insensitive connections
	always @(*) begin
		andOp_201_in0 = valid ? bb_8_active_out_data : bb_8_active_out_data;
		andOp_201_in1 = valid ? eq_200_out : eq_200_out;
	end
	// controller for andOp_202.andOp_202_in0
	// controller for andOp_202.andOp_202_in1
	// Insensitive connections
	always @(*) begin
		andOp_202_in0 = valid ? andOp_201_out : andOp_201_out;
		andOp_202_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_204.andOp_204_in0
	// controller for andOp_204.andOp_204_in1
	// Insensitive connections
	always @(*) begin
		andOp_204_in0 = valid ? eq_203_out : eq_203_out;
		andOp_204_in1 = valid ? andOp_202_out : andOp_202_out;
	end
	// controller for andOp_206.andOp_206_in0
	// controller for andOp_206.andOp_206_in1
	// Insensitive connections
	always @(*) begin
		andOp_206_in0 = valid ? bb_9_active_out_data : bb_9_active_out_data;
		andOp_206_in1 = valid ? eq_205_out : eq_205_out;
	end
	// controller for andOp_207.andOp_207_in0
	// controller for andOp_207.andOp_207_in1
	// Insensitive connections
	always @(*) begin
		andOp_207_in0 = valid ? andOp_206_out : andOp_206_out;
		andOp_207_in1 = valid ? in_read_ready : in_read_ready;
	end
	// controller for andOp_209.andOp_209_in0
	// controller for andOp_209.andOp_209_in1
	// Insensitive connections
	always @(*) begin
		andOp_209_in0 = valid ? eq_208_out : eq_208_out;
		andOp_209_in1 = valid ? andOp_207_out : andOp_207_out;
	end
	// controller for andOp_21.andOp_21_in0
	// controller for andOp_21.andOp_21_in1
	// Insensitive connections
	always @(*) begin
		andOp_21_in0 = valid ? andOp_20_out : andOp_20_out;
		andOp_21_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_212.andOp_212_in0
	// controller for andOp_212.andOp_212_in1
	// Insensitive connections
	always @(*) begin
		andOp_212_in0 = valid ? bb_9_active_out_data : bb_9_active_out_data;
		andOp_212_in1 = valid ? eq_211_out : eq_211_out;
	end
	// controller for andOp_213.andOp_213_in0
	// controller for andOp_213.andOp_213_in1
	// Insensitive connections
	always @(*) begin
		andOp_213_in0 = valid ? andOp_212_out : andOp_212_out;
		andOp_213_in1 = valid ? notOp_210_out : notOp_210_out;
	end
	// controller for andOp_215.andOp_215_in0
	// controller for andOp_215.andOp_215_in1
	// Insensitive connections
	always @(*) begin
		andOp_215_in0 = valid ? eq_214_out : eq_214_out;
		andOp_215_in1 = valid ? andOp_213_out : andOp_213_out;
	end
	// controller for andOp_217.andOp_217_in0
	// controller for andOp_217.andOp_217_in1
	// Insensitive connections
	always @(*) begin
		andOp_217_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_217_in1 = valid ? eq_216_out : eq_216_out;
	end
	// controller for andOp_218.andOp_218_in0
	// controller for andOp_218.andOp_218_in1
	// Insensitive connections
	always @(*) begin
		andOp_218_in0 = valid ? andOp_217_out : andOp_217_out;
		andOp_218_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_220.andOp_220_in0
	// controller for andOp_220.andOp_220_in1
	// Insensitive connections
	always @(*) begin
		andOp_220_in0 = valid ? eq_219_out : eq_219_out;
		andOp_220_in1 = valid ? andOp_218_out : andOp_218_out;
	end
	// controller for andOp_222.andOp_222_in0
	// controller for andOp_222.andOp_222_in1
	// Insensitive connections
	always @(*) begin
		andOp_222_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_222_in1 = valid ? eq_221_out : eq_221_out;
	end
	// controller for andOp_223.andOp_223_in0
	// controller for andOp_223.andOp_223_in1
	// Insensitive connections
	always @(*) begin
		andOp_223_in0 = valid ? andOp_222_out : andOp_222_out;
		andOp_223_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_225.andOp_225_in0
	// controller for andOp_225.andOp_225_in1
	// Insensitive connections
	always @(*) begin
		andOp_225_in0 = valid ? eq_224_out : eq_224_out;
		andOp_225_in1 = valid ? andOp_223_out : andOp_223_out;
	end
	// controller for andOp_227.andOp_227_in0
	// controller for andOp_227.andOp_227_in1
	// Insensitive connections
	always @(*) begin
		andOp_227_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_227_in1 = valid ? eq_226_out : eq_226_out;
	end
	// controller for andOp_228.andOp_228_in0
	// controller for andOp_228.andOp_228_in1
	// Insensitive connections
	always @(*) begin
		andOp_228_in0 = valid ? andOp_227_out : andOp_227_out;
		andOp_228_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_230.andOp_230_in0
	// controller for andOp_230.andOp_230_in1
	// Insensitive connections
	always @(*) begin
		andOp_230_in0 = valid ? eq_229_out : eq_229_out;
		andOp_230_in1 = valid ? andOp_228_out : andOp_228_out;
	end
	// controller for andOp_233.andOp_233_in0
	// controller for andOp_233.andOp_233_in1
	// Insensitive connections
	always @(*) begin
		andOp_233_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_233_in1 = valid ? eq_232_out : eq_232_out;
	end
	// controller for andOp_234.andOp_234_in0
	// controller for andOp_234.andOp_234_in1
	// Insensitive connections
	always @(*) begin
		andOp_234_in0 = valid ? andOp_233_out : andOp_233_out;
		andOp_234_in1 = valid ? notOp_231_out : notOp_231_out;
	end
	// controller for andOp_236.andOp_236_in0
	// controller for andOp_236.andOp_236_in1
	// Insensitive connections
	always @(*) begin
		andOp_236_in0 = valid ? eq_235_out : eq_235_out;
		andOp_236_in1 = valid ? andOp_234_out : andOp_234_out;
	end
	// controller for andOp_238.andOp_238_in0
	// controller for andOp_238.andOp_238_in1
	// Insensitive connections
	always @(*) begin
		andOp_238_in0 = valid ? bb_5_active_out_data : bb_5_active_out_data;
		andOp_238_in1 = valid ? eq_237_out : eq_237_out;
	end
	// controller for andOp_239.andOp_239_in0
	// controller for andOp_239.andOp_239_in1
	// Insensitive connections
	always @(*) begin
		andOp_239_in0 = valid ? andOp_238_out : andOp_238_out;
		andOp_239_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_24.andOp_24_in0
	// controller for andOp_24.andOp_24_in1
	// Insensitive connections
	always @(*) begin
		andOp_24_in0 = valid ? bb_6_active_out_data : bb_6_active_out_data;
		andOp_24_in1 = valid ? eq_23_out : eq_23_out;
	end
	// controller for andOp_241.andOp_241_in0
	// controller for andOp_241.andOp_241_in1
	// Insensitive connections
	always @(*) begin
		andOp_241_in0 = valid ? eq_240_out : eq_240_out;
		andOp_241_in1 = valid ? andOp_239_out : andOp_239_out;
	end
	// controller for andOp_243.andOp_243_in0
	// controller for andOp_243.andOp_243_in1
	// Insensitive connections
	always @(*) begin
		andOp_243_in0 = valid ? bb_6_active_out_data : bb_6_active_out_data;
		andOp_243_in1 = valid ? eq_242_out : eq_242_out;
	end
	// controller for andOp_244.andOp_244_in0
	// controller for andOp_244.andOp_244_in1
	// Insensitive connections
	always @(*) begin
		andOp_244_in0 = valid ? andOp_243_out : andOp_243_out;
		andOp_244_in1 = valid ? out_write_ready : out_write_ready;
	end
	// controller for andOp_246.andOp_246_in0
	// controller for andOp_246.andOp_246_in1
	// Insensitive connections
	always @(*) begin
		andOp_246_in0 = valid ? eq_245_out : eq_245_out;
		andOp_246_in1 = valid ? andOp_244_out : andOp_244_out;
	end
	// controller for andOp_249.andOp_249_in0
	// controller for andOp_249.andOp_249_in1
	// Insensitive connections
	always @(*) begin
		andOp_249_in0 = valid ? bb_6_active_out_data : bb_6_active_out_data;
		andOp_249_in1 = valid ? eq_248_out : eq_248_out;
	end
	// controller for andOp_25.andOp_25_in0
	// controller for andOp_25.andOp_25_in1
	// Insensitive connections
	always @(*) begin
		andOp_25_in0 = valid ? andOp_24_out : andOp_24_out;
		andOp_25_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_250.andOp_250_in0
	// controller for andOp_250.andOp_250_in1
	// Insensitive connections
	always @(*) begin
		andOp_250_in0 = valid ? andOp_249_out : andOp_249_out;
		andOp_250_in1 = valid ? notOp_247_out : notOp_247_out;
	end
	// controller for andOp_252.andOp_252_in0
	// controller for andOp_252.andOp_252_in1
	// Insensitive connections
	always @(*) begin
		andOp_252_in0 = valid ? eq_251_out : eq_251_out;
		andOp_252_in1 = valid ? andOp_250_out : andOp_250_out;
	end
	// controller for andOp_254.andOp_254_in0
	// controller for andOp_254.andOp_254_in1
	// Insensitive connections
	always @(*) begin
		andOp_254_in0 = valid ? bb_7_active_out_data : bb_7_active_out_data;
		andOp_254_in1 = valid ? eq_253_out : eq_253_out;
	end
	// controller for andOp_255.andOp_255_in0
	// controller for andOp_255.andOp_255_in1
	// Insensitive connections
	always @(*) begin
		andOp_255_in0 = valid ? andOp_254_out : andOp_254_out;
		andOp_255_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_257.andOp_257_in0
	// controller for andOp_257.andOp_257_in1
	// Insensitive connections
	always @(*) begin
		andOp_257_in0 = valid ? eq_256_out : eq_256_out;
		andOp_257_in1 = valid ? andOp_255_out : andOp_255_out;
	end
	// controller for andOp_259.andOp_259_in0
	// controller for andOp_259.andOp_259_in1
	// Insensitive connections
	always @(*) begin
		andOp_259_in0 = valid ? bb_2_active_out_data : bb_2_active_out_data;
		andOp_259_in1 = valid ? eq_258_out : eq_258_out;
	end
	// controller for andOp_260.andOp_260_in0
	// controller for andOp_260.andOp_260_in1
	// Insensitive connections
	always @(*) begin
		andOp_260_in0 = valid ? andOp_259_out : andOp_259_out;
		andOp_260_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_262.andOp_262_in0
	// controller for andOp_262.andOp_262_in1
	// Insensitive connections
	always @(*) begin
		andOp_262_in0 = valid ? eq_261_out : eq_261_out;
		andOp_262_in1 = valid ? andOp_260_out : andOp_260_out;
	end
	// controller for andOp_264.andOp_264_in0
	// controller for andOp_264.andOp_264_in1
	// Insensitive connections
	always @(*) begin
		andOp_264_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_264_in1 = valid ? eq_263_out : eq_263_out;
	end
	// controller for andOp_266.andOp_266_in0
	// controller for andOp_266.andOp_266_in1
	// Insensitive connections
	always @(*) begin
		andOp_266_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_266_in1 = valid ? eq_265_out : eq_265_out;
	end
	// controller for andOp_268.andOp_268_in0
	// controller for andOp_268.andOp_268_in1
	// Insensitive connections
	always @(*) begin
		andOp_268_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_268_in1 = valid ? eq_267_out : eq_267_out;
	end
	// controller for andOp_27.andOp_27_in0
	// controller for andOp_27.andOp_27_in1
	// Insensitive connections
	always @(*) begin
		andOp_27_in0 = valid ? andOp_25_out : andOp_25_out;
		andOp_27_in1 = valid ? out_write_ready : out_write_ready;
	end
	// controller for andOp_270.andOp_270_in0
	// controller for andOp_270.andOp_270_in1
	// Insensitive connections
	always @(*) begin
		andOp_270_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_270_in1 = valid ? eq_269_out : eq_269_out;
	end
	// controller for andOp_272.andOp_272_in0
	// controller for andOp_272.andOp_272_in1
	// Insensitive connections
	always @(*) begin
		andOp_272_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_272_in1 = valid ? eq_271_out : eq_271_out;
	end
	// controller for andOp_274.andOp_274_in0
	// controller for andOp_274.andOp_274_in1
	// Insensitive connections
	always @(*) begin
		andOp_274_in0 = valid ? bb_3_active_out_data : bb_3_active_out_data;
		andOp_274_in1 = valid ? eq_273_out : eq_273_out;
	end
	// controller for andOp_276.andOp_276_in0
	// controller for andOp_276.andOp_276_in1
	// Insensitive connections
	always @(*) begin
		andOp_276_in0 = valid ? bb_3_active_out_data : bb_3_active_out_data;
		andOp_276_in1 = valid ? eq_275_out : eq_275_out;
	end
	// controller for andOp_277.andOp_277_in0
	// controller for andOp_277.andOp_277_in1
	// Insensitive connections
	always @(*) begin
		andOp_277_in0 = valid ? andOp_274_out : andOp_274_out;
		andOp_277_in1 = valid ? andOp_276_out : andOp_276_out;
	end
	// controller for andOp_279.andOp_279_in0
	// controller for andOp_279.andOp_279_in1
	// Insensitive connections
	always @(*) begin
		andOp_279_in0 = valid ? bb_3_active_out_data : bb_3_active_out_data;
		andOp_279_in1 = valid ? eq_278_out : eq_278_out;
	end
	// controller for andOp_281.andOp_281_in0
	// controller for andOp_281.andOp_281_in1
	// Insensitive connections
	always @(*) begin
		andOp_281_in0 = valid ? bb_8_active_out_data : bb_8_active_out_data;
		andOp_281_in1 = valid ? eq_280_out : eq_280_out;
	end
	// controller for andOp_283.andOp_283_in0
	// controller for andOp_283.andOp_283_in1
	// Insensitive connections
	always @(*) begin
		andOp_283_in0 = valid ? bb_9_active_out_data : bb_9_active_out_data;
		andOp_283_in1 = valid ? eq_282_out : eq_282_out;
	end
	// controller for andOp_285.andOp_285_in0
	// controller for andOp_285.andOp_285_in1
	// Insensitive connections
	always @(*) begin
		andOp_285_in0 = valid ? bb_9_active_out_data : bb_9_active_out_data;
		andOp_285_in1 = valid ? eq_284_out : eq_284_out;
	end
	// controller for andOp_287.andOp_287_in0
	// controller for andOp_287.andOp_287_in1
	// Insensitive connections
	always @(*) begin
		andOp_287_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_287_in1 = valid ? eq_286_out : eq_286_out;
	end
	// controller for andOp_289.andOp_289_in0
	// controller for andOp_289.andOp_289_in1
	// Insensitive connections
	always @(*) begin
		andOp_289_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_289_in1 = valid ? eq_288_out : eq_288_out;
	end
	// controller for andOp_29.andOp_29_in0
	// controller for andOp_29.andOp_29_in1
	// Insensitive connections
	always @(*) begin
		andOp_29_in0 = valid ? andOp_25_out : andOp_25_out;
		andOp_29_in1 = valid ? notOp_28_out : notOp_28_out;
	end
	// controller for andOp_291.andOp_291_in0
	// controller for andOp_291.andOp_291_in1
	// Insensitive connections
	always @(*) begin
		andOp_291_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_291_in1 = valid ? eq_290_out : eq_290_out;
	end
	// controller for andOp_293.andOp_293_in0
	// controller for andOp_293.andOp_293_in1
	// Insensitive connections
	always @(*) begin
		andOp_293_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_293_in1 = valid ? eq_292_out : eq_292_out;
	end
	// controller for andOp_294.andOp_294_in0
	// controller for andOp_294.andOp_294_in1
	// Insensitive connections
	always @(*) begin
		andOp_294_in0 = valid ? andOp_291_out : andOp_291_out;
		andOp_294_in1 = valid ? andOp_293_out : andOp_293_out;
	end
	// controller for andOp_296.andOp_296_in0
	// controller for andOp_296.andOp_296_in1
	// Insensitive connections
	always @(*) begin
		andOp_296_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_296_in1 = valid ? eq_295_out : eq_295_out;
	end
	// controller for andOp_298.andOp_298_in0
	// controller for andOp_298.andOp_298_in1
	// Insensitive connections
	always @(*) begin
		andOp_298_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_298_in1 = valid ? eq_297_out : eq_297_out;
	end
	// controller for andOp_300.andOp_300_in0
	// controller for andOp_300.andOp_300_in1
	// Insensitive connections
	always @(*) begin
		andOp_300_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_300_in1 = valid ? eq_299_out : eq_299_out;
	end
	// controller for andOp_302.andOp_302_in0
	// controller for andOp_302.andOp_302_in1
	// Insensitive connections
	always @(*) begin
		andOp_302_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_302_in1 = valid ? eq_301_out : eq_301_out;
	end
	// controller for andOp_303.andOp_303_in0
	// controller for andOp_303.andOp_303_in1
	// Insensitive connections
	always @(*) begin
		andOp_303_in0 = valid ? andOp_300_out : andOp_300_out;
		andOp_303_in1 = valid ? andOp_302_out : andOp_302_out;
	end
	// controller for andOp_305.andOp_305_in0
	// controller for andOp_305.andOp_305_in1
	// Insensitive connections
	always @(*) begin
		andOp_305_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_305_in1 = valid ? eq_304_out : eq_304_out;
	end
	// controller for andOp_307.andOp_307_in0
	// controller for andOp_307.andOp_307_in1
	// Insensitive connections
	always @(*) begin
		andOp_307_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_307_in1 = valid ? eq_306_out : eq_306_out;
	end
	// controller for andOp_308.andOp_308_in0
	// controller for andOp_308.andOp_308_in1
	// Insensitive connections
	always @(*) begin
		andOp_308_in0 = valid ? andOp_305_out : andOp_305_out;
		andOp_308_in1 = valid ? andOp_307_out : andOp_307_out;
	end
	// controller for andOp_31.andOp_31_in0
	// controller for andOp_31.andOp_31_in1
	// Insensitive connections
	always @(*) begin
		andOp_31_in0 = valid ? bb_7_active_out_data : bb_7_active_out_data;
		andOp_31_in1 = valid ? eq_30_out : eq_30_out;
	end
	// controller for andOp_310.andOp_310_in0
	// controller for andOp_310.andOp_310_in1
	// Insensitive connections
	always @(*) begin
		andOp_310_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_310_in1 = valid ? eq_309_out : eq_309_out;
	end
	// controller for andOp_312.andOp_312_in0
	// controller for andOp_312.andOp_312_in1
	// Insensitive connections
	always @(*) begin
		andOp_312_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_312_in1 = valid ? eq_311_out : eq_311_out;
	end
	// controller for andOp_314.andOp_314_in0
	// controller for andOp_314.andOp_314_in1
	// Insensitive connections
	always @(*) begin
		andOp_314_in0 = valid ? bb_1_active_out_data : bb_1_active_out_data;
		andOp_314_in1 = valid ? eq_313_out : eq_313_out;
	end
	// controller for andOp_316.andOp_316_in0
	// controller for andOp_316.andOp_316_in1
	// Insensitive connections
	always @(*) begin
		andOp_316_in0 = valid ? bb_5_active_out_data : bb_5_active_out_data;
		andOp_316_in1 = valid ? eq_315_out : eq_315_out;
	end
	// controller for andOp_318.andOp_318_in0
	// controller for andOp_318.andOp_318_in1
	// Insensitive connections
	always @(*) begin
		andOp_318_in0 = valid ? bb_6_active_out_data : bb_6_active_out_data;
		andOp_318_in1 = valid ? eq_317_out : eq_317_out;
	end
	// controller for andOp_32.andOp_32_in0
	// controller for andOp_32.andOp_32_in1
	// Insensitive connections
	always @(*) begin
		andOp_32_in0 = valid ? andOp_31_out : andOp_31_out;
		andOp_32_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_320.andOp_320_in0
	// controller for andOp_320.andOp_320_in1
	// Insensitive connections
	always @(*) begin
		andOp_320_in0 = valid ? bb_6_active_out_data : bb_6_active_out_data;
		andOp_320_in1 = valid ? eq_319_out : eq_319_out;
	end
	// controller for andOp_322.andOp_322_in0
	// controller for andOp_322.andOp_322_in1
	// Insensitive connections
	always @(*) begin
		andOp_322_in0 = valid ? bb_7_active_out_data : bb_7_active_out_data;
		andOp_322_in1 = valid ? eq_321_out : eq_321_out;
	end
	// controller for andOp_324.andOp_324_in0
	// controller for andOp_324.andOp_324_in1
	// Insensitive connections
	always @(*) begin
		andOp_324_in0 = valid ? bb_7_active_out_data : bb_7_active_out_data;
		andOp_324_in1 = valid ? eq_323_out : eq_323_out;
	end
	// controller for andOp_326.andOp_326_in0
	// controller for andOp_326.andOp_326_in1
	// Insensitive connections
	always @(*) begin
		andOp_326_in0 = valid ? bb_7_active_out_data : bb_7_active_out_data;
		andOp_326_in1 = valid ? eq_325_out : eq_325_out;
	end
	// controller for andOp_328.andOp_328_in0
	// controller for andOp_328.andOp_328_in1
	// Insensitive connections
	always @(*) begin
		andOp_328_in0 = valid ? bb_7_active_out_data : bb_7_active_out_data;
		andOp_328_in1 = valid ? eq_327_out : eq_327_out;
	end
	// controller for andOp_330.andOp_330_in0
	// controller for andOp_330.andOp_330_in1
	// Insensitive connections
	always @(*) begin
		andOp_330_in0 = valid ? bb_2_active_out_data : bb_2_active_out_data;
		andOp_330_in1 = valid ? eq_329_out : eq_329_out;
	end
	// controller for andOp_332.andOp_332_in0
	// controller for andOp_332.andOp_332_in1
	// Insensitive connections
	always @(*) begin
		andOp_332_in0 = valid ? bb_2_active_out_data : bb_2_active_out_data;
		andOp_332_in1 = valid ? eq_331_out : eq_331_out;
	end
	// controller for andOp_35.andOp_35_in0
	// controller for andOp_35.andOp_35_in1
	// Insensitive connections
	always @(*) begin
		andOp_35_in0 = valid ? bb_8_active_out_data : bb_8_active_out_data;
		andOp_35_in1 = valid ? eq_34_out : eq_34_out;
	end
	// controller for andOp_36.andOp_36_in0
	// controller for andOp_36.andOp_36_in1
	// Insensitive connections
	always @(*) begin
		andOp_36_in0 = valid ? andOp_35_out : andOp_35_out;
		andOp_36_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_39.andOp_39_in0
	// controller for andOp_39.andOp_39_in1
	// Insensitive connections
	always @(*) begin
		andOp_39_in0 = valid ? bb_9_active_out_data : bb_9_active_out_data;
		andOp_39_in1 = valid ? eq_38_out : eq_38_out;
	end
	// controller for andOp_40.andOp_40_in0
	// controller for andOp_40.andOp_40_in1
	// Insensitive connections
	always @(*) begin
		andOp_40_in0 = valid ? andOp_39_out : andOp_39_out;
		andOp_40_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_42.andOp_42_in0
	// controller for andOp_42.andOp_42_in1
	// Insensitive connections
	always @(*) begin
		andOp_42_in0 = valid ? andOp_40_out : andOp_40_out;
		andOp_42_in1 = valid ? in_read_ready : in_read_ready;
	end
	// controller for andOp_44.andOp_44_in0
	// controller for andOp_44.andOp_44_in1
	// Insensitive connections
	always @(*) begin
		andOp_44_in0 = valid ? andOp_40_out : andOp_40_out;
		andOp_44_in1 = valid ? notOp_43_out : notOp_43_out;
	end
	// controller for andOp_46.andOp_46_in0
	// controller for andOp_46.andOp_46_in1
	// Insensitive connections
	always @(*) begin
		andOp_46_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_46_in1 = valid ? eq_45_out : eq_45_out;
	end
	// controller for andOp_47.andOp_47_in0
	// controller for andOp_47.andOp_47_in1
	// Insensitive connections
	always @(*) begin
		andOp_47_in0 = valid ? andOp_46_out : andOp_46_out;
		andOp_47_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_5.andOp_5_in0
	// controller for andOp_5.andOp_5_in1
	// Insensitive connections
	always @(*) begin
		andOp_5_in0 = valid ? bb_1_active_out_data : bb_1_active_out_data;
		andOp_5_in1 = valid ? eq_4_out : eq_4_out;
	end
	// controller for andOp_6.andOp_6_in0
	// controller for andOp_6.andOp_6_in1
	// Insensitive connections
	always @(*) begin
		andOp_6_in0 = valid ? andOp_5_out : andOp_5_out;
		andOp_6_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_65.andOp_65_in0
	// controller for andOp_65.andOp_65_in1
	// Insensitive connections
	always @(*) begin
		andOp_65_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_65_in1 = valid ? eq_64_out : eq_64_out;
	end
	// controller for andOp_67.andOp_67_in0
	// controller for andOp_67.andOp_67_in1
	// Insensitive connections
	always @(*) begin
		andOp_67_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_67_in1 = valid ? eq_66_out : eq_66_out;
	end
	// controller for andOp_69.andOp_69_in0
	// controller for andOp_69.andOp_69_in1
	// Insensitive connections
	always @(*) begin
		andOp_69_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_69_in1 = valid ? eq_68_out : eq_68_out;
	end
	// controller for andOp_71.andOp_71_in0
	// controller for andOp_71.andOp_71_in1
	// Insensitive connections
	always @(*) begin
		andOp_71_in0 = valid ? bb_2_active_out_data : bb_2_active_out_data;
		andOp_71_in1 = valid ? eq_70_out : eq_70_out;
	end
	// controller for andOp_75.andOp_75_in0
	// controller for andOp_75.andOp_75_in1
	// Insensitive connections
	always @(*) begin
		andOp_75_in0 = valid ? notOp_74_out : notOp_74_out;
		andOp_75_in1 = valid ? andOp_16_out : andOp_16_out;
	end
	// controller for andOp_79.andOp_79_in0
	// controller for andOp_79.andOp_79_in1
	// Insensitive connections
	always @(*) begin
		andOp_79_in0 = valid ? notOp_78_out : notOp_78_out;
		andOp_79_in1 = valid ? andOp_2_out : andOp_2_out;
	end
	// controller for andOp_83.andOp_83_in0
	// controller for andOp_83.andOp_83_in1
	// Insensitive connections
	always @(*) begin
		andOp_83_in0 = valid ? notOp_82_out : notOp_82_out;
		andOp_83_in1 = valid ? andOp_6_out : andOp_6_out;
	end
	// controller for andOp_88.andOp_88_in0
	// controller for andOp_88.andOp_88_in1
	// Insensitive connections
	always @(*) begin
		andOp_88_in0 = valid ? notOp_87_out : notOp_87_out;
		andOp_88_in1 = valid ? andOp_10_out : andOp_10_out;
	end
	// controller for andOp_9.andOp_9_in0
	// controller for andOp_9.andOp_9_in1
	// Insensitive connections
	always @(*) begin
		andOp_9_in0 = valid ? bb_3_active_out_data : bb_3_active_out_data;
		andOp_9_in1 = valid ? eq_8_out : eq_8_out;
	end
	// controller for andOp_92.andOp_92_in0
	// controller for andOp_92.andOp_92_in1
	// Insensitive connections
	always @(*) begin
		andOp_92_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_92_in1 = valid ? eq_91_out : eq_91_out;
	end
	// controller for andOp_94.andOp_94_in0
	// controller for andOp_94.andOp_94_in1
	// Insensitive connections
	always @(*) begin
		andOp_94_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_94_in1 = valid ? eq_93_out : eq_93_out;
	end
	// controller for andOp_96.andOp_96_in0
	// controller for andOp_96.andOp_96_in1
	// Insensitive connections
	always @(*) begin
		andOp_96_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_96_in1 = valid ? eq_95_out : eq_95_out;
	end
	// controller for andOp_98.andOp_98_in0
	// controller for andOp_98.andOp_98_in1
	// Insensitive connections
	always @(*) begin
		andOp_98_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_98_in1 = valid ? eq_97_out : eq_97_out;
	end
	// controller for bb_0_active.bb_0_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_data = eq_49_out;
		end else begin
			bb_0_active_in_data = 0;
		end
	end
	// controller for bb_0_predecessor.bb_0_predecessor_in_data
	always @(*) begin
		if (eq_72_out) begin 
			bb_0_predecessor_in_data = last_BB_reg;
		end else begin
			bb_0_predecessor_in_data = 0;
		end
	end
	// controller for bb_10_active.bb_10_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_data = eq_63_out;
		end else begin
			bb_10_active_in_data = 0;
		end
	end
	// controller for bb_10_predecessor.bb_10_predecessor_in_data
	always @(*) begin
		if (eq_90_out) begin 
			bb_10_predecessor_in_data = last_BB_reg;
		end else begin
			bb_10_predecessor_in_data = 0;
		end
	end
	// controller for bb_1_active.bb_1_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_data = orOp_51_out;
		end else begin
			bb_1_active_in_data = 0;
		end
	end
	// controller for bb_1_predecessor.bb_1_predecessor_in_data
	always @(*) begin
		if (andOp_75_out) begin 
			bb_1_predecessor_in_data = 32'd4;
		end else if (eq_73_out) begin 
			bb_1_predecessor_in_data = last_BB_reg;
		end else begin
			bb_1_predecessor_in_data = 0;
		end
	end
	// controller for bb_2_active.bb_2_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_data = eq_52_out;
		end else begin
			bb_2_active_in_data = 0;
		end
	end
	// controller for bb_2_predecessor.bb_2_predecessor_in_data
	always @(*) begin
		if (eq_76_out) begin 
			bb_2_predecessor_in_data = last_BB_reg;
		end else begin
			bb_2_predecessor_in_data = 0;
		end
	end
	// controller for bb_3_active.bb_3_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_data = orOp_54_out;
		end else begin
			bb_3_active_in_data = 0;
		end
	end
	// controller for bb_3_predecessor.bb_3_predecessor_in_data
	always @(*) begin
		if (andOp_79_out) begin 
			bb_3_predecessor_in_data = 32'd0;
		end else if (eq_77_out) begin 
			bb_3_predecessor_in_data = last_BB_reg;
		end else begin
			bb_3_predecessor_in_data = 0;
		end
	end
	// controller for bb_4_active.bb_4_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_data = eq_55_out;
		end else begin
			bb_4_active_in_data = 0;
		end
	end
	// controller for bb_4_predecessor.bb_4_predecessor_in_data
	always @(*) begin
		if (eq_80_out) begin 
			bb_4_predecessor_in_data = last_BB_reg;
		end else begin
			bb_4_predecessor_in_data = 0;
		end
	end
	// controller for bb_5_active.bb_5_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_5_active_in_data = orOp_57_out;
		end else begin
			bb_5_active_in_data = 0;
		end
	end
	// controller for bb_5_predecessor.bb_5_predecessor_in_data
	always @(*) begin
		if (andOp_83_out) begin 
			bb_5_predecessor_in_data = 32'd1;
		end else if (eq_81_out) begin 
			bb_5_predecessor_in_data = last_BB_reg;
		end else begin
			bb_5_predecessor_in_data = 0;
		end
	end
	// controller for bb_6_active.bb_6_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_6_active_in_data = eq_58_out;
		end else begin
			bb_6_active_in_data = 0;
		end
	end
	// controller for bb_6_predecessor.bb_6_predecessor_in_data
	always @(*) begin
		if (eq_84_out) begin 
			bb_6_predecessor_in_data = last_BB_reg;
		end else begin
			bb_6_predecessor_in_data = 0;
		end
	end
	// controller for bb_7_active.bb_7_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_7_active_in_data = eq_59_out;
		end else begin
			bb_7_active_in_data = 0;
		end
	end
	// controller for bb_7_predecessor.bb_7_predecessor_in_data
	always @(*) begin
		if (eq_85_out) begin 
			bb_7_predecessor_in_data = last_BB_reg;
		end else begin
			bb_7_predecessor_in_data = 0;
		end
	end
	// controller for bb_8_active.bb_8_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_data = orOp_61_out;
		end else begin
			bb_8_active_in_data = 0;
		end
	end
	// controller for bb_8_predecessor.bb_8_predecessor_in_data
	always @(*) begin
		if (andOp_88_out) begin 
			bb_8_predecessor_in_data = 32'd3;
		end else if (eq_86_out) begin 
			bb_8_predecessor_in_data = last_BB_reg;
		end else begin
			bb_8_predecessor_in_data = 0;
		end
	end
	// controller for bb_9_active.bb_9_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_9_active_in_data = eq_62_out;
		end else begin
			bb_9_active_in_data = 0;
		end
	end
	// controller for bb_9_predecessor.bb_9_predecessor_in_data
	always @(*) begin
		if (eq_89_out) begin 
			bb_9_predecessor_in_data = last_BB_reg;
		end else begin
			bb_9_predecessor_in_data = 0;
		end
	end
	// controller for br_0_happened.br_0_happened_in_data
	always @(*) begin
		if (andOp_2_out) begin 
			br_0_happened_in_data = 1'd1;
		end else if (notOp_3_out) begin 
			br_0_happened_in_data = 1'd0;
		end else begin
			br_0_happened_in_data = 0;
		end
	end
	// controller for br_10_happened.br_10_happened_in_data
	always @(*) begin
		if (andOp_47_out) begin 
			br_10_happened_in_data = 1'd1;
		end else if (notOp_48_out) begin 
			br_10_happened_in_data = 1'd0;
		end else begin
			br_10_happened_in_data = 0;
		end
	end
	// controller for br_1_happened.br_1_happened_in_data
	always @(*) begin
		if (andOp_6_out) begin 
			br_1_happened_in_data = 1'd1;
		end else if (notOp_7_out) begin 
			br_1_happened_in_data = 1'd0;
		end else begin
			br_1_happened_in_data = 0;
		end
	end
	// controller for br_3_happened.br_3_happened_in_data
	always @(*) begin
		if (andOp_10_out) begin 
			br_3_happened_in_data = 1'd1;
		end else if (notOp_11_out) begin 
			br_3_happened_in_data = 1'd0;
		end else begin
			br_3_happened_in_data = 0;
		end
	end
	// controller for br_4_happened.br_4_happened_in_data
	always @(*) begin
		if (andOp_14_out) begin 
			br_4_happened_in_data = 1'd1;
		end else if (notOp_15_out) begin 
			br_4_happened_in_data = 1'd0;
		end else begin
			br_4_happened_in_data = 0;
		end
	end
	// controller for br_5_happened.br_5_happened_in_data
	always @(*) begin
		if (andOp_21_out) begin 
			br_5_happened_in_data = 1'd1;
		end else if (notOp_22_out) begin 
			br_5_happened_in_data = 1'd0;
		end else begin
			br_5_happened_in_data = 0;
		end
	end
	// controller for br_6_happened.br_6_happened_in_data
	always @(*) begin
		if (andOp_25_out) begin 
			br_6_happened_in_data = 1'd1;
		end else if (notOp_26_out) begin 
			br_6_happened_in_data = 1'd0;
		end else begin
			br_6_happened_in_data = 0;
		end
	end
	// controller for br_7_happened.br_7_happened_in_data
	always @(*) begin
		if (andOp_32_out) begin 
			br_7_happened_in_data = 1'd1;
		end else if (notOp_33_out) begin 
			br_7_happened_in_data = 1'd0;
		end else begin
			br_7_happened_in_data = 0;
		end
	end
	// controller for br_8_happened.br_8_happened_in_data
	always @(*) begin
		if (andOp_36_out) begin 
			br_8_happened_in_data = 1'd1;
		end else if (notOp_37_out) begin 
			br_8_happened_in_data = 1'd0;
		end else begin
			br_8_happened_in_data = 0;
		end
	end
	// controller for br_9_happened.br_9_happened_in_data
	always @(*) begin
		if (andOp_40_out) begin 
			br_9_happened_in_data = 1'd1;
		end else if (notOp_41_out) begin 
			br_9_happened_in_data = 1'd0;
		end else begin
			br_9_happened_in_data = 0;
		end
	end
	// controller for eq_0.eq_0_in0
	// controller for eq_0.eq_0_in1
	// Insensitive connections
	always @(*) begin
		eq_0_in0 = valid ? 32'd1 : 32'd1;
		eq_0_in1 = valid ? global_state : global_state;
	end
	// controller for eq_101.eq_101_in0
	// controller for eq_101.eq_101_in1
	// Insensitive connections
	always @(*) begin
		eq_101_in0 = valid ? 32'd5 : 32'd5;
		eq_101_in1 = valid ? global_state : global_state;
	end
	// controller for eq_103.eq_103_in0
	// controller for eq_103.eq_103_in1
	// Insensitive connections
	always @(*) begin
		eq_103_in0 = valid ? 32'd8 : 32'd8;
		eq_103_in1 = valid ? global_state : global_state;
	end
	// controller for eq_105.eq_105_in0
	// controller for eq_105.eq_105_in1
	// Insensitive connections
	always @(*) begin
		eq_105_in0 = valid ? 32'd1 : 32'd1;
		eq_105_in1 = valid ? global_state : global_state;
	end
	// controller for eq_107.eq_107_in0
	// controller for eq_107.eq_107_in1
	// Insensitive connections
	always @(*) begin
		eq_107_in0 = valid ? 32'd2 : 32'd2;
		eq_107_in1 = valid ? global_state : global_state;
	end
	// controller for eq_109.eq_109_in0
	// controller for eq_109.eq_109_in1
	// Insensitive connections
	always @(*) begin
		eq_109_in0 = valid ? 32'd3 : 32'd3;
		eq_109_in1 = valid ? global_state : global_state;
	end
	// controller for eq_111.eq_111_in0
	// controller for eq_111.eq_111_in1
	// Insensitive connections
	always @(*) begin
		eq_111_in0 = valid ? 32'd4 : 32'd4;
		eq_111_in1 = valid ? global_state : global_state;
	end
	// controller for eq_113.eq_113_in0
	// controller for eq_113.eq_113_in1
	// Insensitive connections
	always @(*) begin
		eq_113_in0 = valid ? 32'd5 : 32'd5;
		eq_113_in1 = valid ? global_state : global_state;
	end
	// controller for eq_115.eq_115_in0
	// controller for eq_115.eq_115_in1
	// Insensitive connections
	always @(*) begin
		eq_115_in0 = valid ? 32'd5 : 32'd5;
		eq_115_in1 = valid ? global_state : global_state;
	end
	// controller for eq_117.eq_117_in0
	// controller for eq_117.eq_117_in1
	// Insensitive connections
	always @(*) begin
		eq_117_in0 = valid ? 32'd5 : 32'd5;
		eq_117_in1 = valid ? global_state : global_state;
	end
	// controller for eq_119.eq_119_in0
	// controller for eq_119.eq_119_in1
	// Insensitive connections
	always @(*) begin
		eq_119_in0 = valid ? 32'd7 : 32'd7;
		eq_119_in1 = valid ? global_state : global_state;
	end
	// controller for eq_12.eq_12_in0
	// controller for eq_12.eq_12_in1
	// Insensitive connections
	always @(*) begin
		eq_12_in0 = valid ? 32'd6 : 32'd6;
		eq_12_in1 = valid ? global_state : global_state;
	end
	// controller for eq_121.eq_121_in0
	// controller for eq_121.eq_121_in1
	// Insensitive connections
	always @(*) begin
		eq_121_in0 = valid ? 32'd8 : 32'd8;
		eq_121_in1 = valid ? global_state : global_state;
	end
	// controller for eq_123.eq_123_in0
	// controller for eq_123.eq_123_in1
	// Insensitive connections
	always @(*) begin
		eq_123_in0 = valid ? 32'd8 : 32'd8;
		eq_123_in1 = valid ? global_state : global_state;
	end
	// controller for eq_125.eq_125_in0
	// controller for eq_125.eq_125_in1
	// Insensitive connections
	always @(*) begin
		eq_125_in0 = valid ? 32'd9 : 32'd9;
		eq_125_in1 = valid ? global_state : global_state;
	end
	// controller for eq_127.eq_127_in0
	// controller for eq_127.eq_127_in1
	// Insensitive connections
	always @(*) begin
		eq_127_in0 = valid ? 32'd9 : 32'd9;
		eq_127_in1 = valid ? global_state : global_state;
	end
	// controller for eq_129.eq_129_in0
	// controller for eq_129.eq_129_in1
	// Insensitive connections
	always @(*) begin
		eq_129_in0 = valid ? 32'd1 : 32'd1;
		eq_129_in1 = valid ? global_state : global_state;
	end
	// controller for eq_131.eq_131_in0
	// controller for eq_131.eq_131_in1
	// Insensitive connections
	always @(*) begin
		eq_131_in0 = valid ? 32'd1 : 32'd1;
		eq_131_in1 = valid ? global_state : global_state;
	end
	// controller for eq_135.eq_135_in0
	// controller for eq_135.eq_135_in1
	// Insensitive connections
	always @(*) begin
		eq_135_in0 = valid ? 32'd1 : 32'd1;
		eq_135_in1 = valid ? global_state : global_state;
	end
	// controller for eq_137.eq_137_in0
	// controller for eq_137.eq_137_in1
	// Insensitive connections
	always @(*) begin
		eq_137_in0 = valid ? 32'd1 : 32'd1;
		eq_137_in1 = valid ? global_state : global_state;
	end
	// controller for eq_141.eq_141_in0
	// controller for eq_141.eq_141_in1
	// Insensitive connections
	always @(*) begin
		eq_141_in0 = valid ? 32'd1 : 32'd1;
		eq_141_in1 = valid ? global_state : global_state;
	end
	// controller for eq_143.eq_143_in0
	// controller for eq_143.eq_143_in1
	// Insensitive connections
	always @(*) begin
		eq_143_in0 = valid ? 32'd1 : 32'd1;
		eq_143_in1 = valid ? global_state : global_state;
	end
	// controller for eq_147.eq_147_in0
	// controller for eq_147.eq_147_in1
	// Insensitive connections
	always @(*) begin
		eq_147_in0 = valid ? 32'd2 : 32'd2;
		eq_147_in1 = valid ? global_state : global_state;
	end
	// controller for eq_149.eq_149_in0
	// controller for eq_149.eq_149_in1
	// Insensitive connections
	always @(*) begin
		eq_149_in0 = valid ? 32'd2 : 32'd2;
		eq_149_in1 = valid ? global_state : global_state;
	end
	// controller for eq_153.eq_153_in0
	// controller for eq_153.eq_153_in1
	// Insensitive connections
	always @(*) begin
		eq_153_in0 = valid ? 32'd4 : 32'd4;
		eq_153_in1 = valid ? global_state : global_state;
	end
	// controller for eq_155.eq_155_in0
	// controller for eq_155.eq_155_in1
	// Insensitive connections
	always @(*) begin
		eq_155_in0 = valid ? 32'd4 : 32'd4;
		eq_155_in1 = valid ? global_state : global_state;
	end
	// controller for eq_159.eq_159_in0
	// controller for eq_159.eq_159_in1
	// Insensitive connections
	always @(*) begin
		eq_159_in0 = valid ? 32'd6 : 32'd6;
		eq_159_in1 = valid ? global_state : global_state;
	end
	// controller for eq_161.eq_161_in0
	// controller for eq_161.eq_161_in1
	// Insensitive connections
	always @(*) begin
		eq_161_in0 = valid ? 32'd6 : 32'd6;
		eq_161_in1 = valid ? global_state : global_state;
	end
	// controller for eq_165.eq_165_in0
	// controller for eq_165.eq_165_in1
	// Insensitive connections
	always @(*) begin
		eq_165_in0 = valid ? 32'd6 : 32'd6;
		eq_165_in1 = valid ? global_state : global_state;
	end
	// controller for eq_169.eq_169_in0
	// controller for eq_169.eq_169_in1
	// Insensitive connections
	always @(*) begin
		eq_169_in0 = valid ? 32'd6 : 32'd6;
		eq_169_in1 = valid ? global_state : global_state;
	end
	// controller for eq_171.eq_171_in0
	// controller for eq_171.eq_171_in1
	// Insensitive connections
	always @(*) begin
		eq_171_in0 = valid ? 32'd6 : 32'd6;
		eq_171_in1 = valid ? global_state : global_state;
	end
	// controller for eq_175.eq_175_in0
	// controller for eq_175.eq_175_in1
	// Insensitive connections
	always @(*) begin
		eq_175_in0 = valid ? 32'd6 : 32'd6;
		eq_175_in1 = valid ? global_state : global_state;
	end
	// controller for eq_177.eq_177_in0
	// controller for eq_177.eq_177_in1
	// Insensitive connections
	always @(*) begin
		eq_177_in0 = valid ? 32'd6 : 32'd6;
		eq_177_in1 = valid ? global_state : global_state;
	end
	// controller for eq_181.eq_181_in0
	// controller for eq_181.eq_181_in1
	// Insensitive connections
	always @(*) begin
		eq_181_in0 = valid ? 32'd7 : 32'd7;
		eq_181_in1 = valid ? global_state : global_state;
	end
	// controller for eq_183.eq_183_in0
	// controller for eq_183.eq_183_in1
	// Insensitive connections
	always @(*) begin
		eq_183_in0 = valid ? 32'd7 : 32'd7;
		eq_183_in1 = valid ? global_state : global_state;
	end
	// controller for eq_187.eq_187_in0
	// controller for eq_187.eq_187_in1
	// Insensitive connections
	always @(*) begin
		eq_187_in0 = valid ? 32'd8 : 32'd8;
		eq_187_in1 = valid ? global_state : global_state;
	end
	// controller for eq_189.eq_189_in0
	// controller for eq_189.eq_189_in1
	// Insensitive connections
	always @(*) begin
		eq_189_in0 = valid ? 32'd8 : 32'd8;
		eq_189_in1 = valid ? global_state : global_state;
	end
	// controller for eq_19.eq_19_in0
	// controller for eq_19.eq_19_in1
	// Insensitive connections
	always @(*) begin
		eq_19_in0 = valid ? 32'd6 : 32'd6;
		eq_19_in1 = valid ? global_state : global_state;
	end
	// controller for eq_193.eq_193_in0
	// controller for eq_193.eq_193_in1
	// Insensitive connections
	always @(*) begin
		eq_193_in0 = valid ? 32'd9 : 32'd9;
		eq_193_in1 = valid ? global_state : global_state;
	end
	// controller for eq_195.eq_195_in0
	// controller for eq_195.eq_195_in1
	// Insensitive connections
	always @(*) begin
		eq_195_in0 = valid ? 32'd0 : 32'd0;
		eq_195_in1 = valid ? global_state : global_state;
	end
	// controller for eq_198.eq_198_in0
	// controller for eq_198.eq_198_in1
	// Insensitive connections
	always @(*) begin
		eq_198_in0 = valid ? 32'd0 : 32'd0;
		eq_198_in1 = valid ? global_state : global_state;
	end
	// controller for eq_200.eq_200_in0
	// controller for eq_200.eq_200_in1
	// Insensitive connections
	always @(*) begin
		eq_200_in0 = valid ? 32'd1 : 32'd1;
		eq_200_in1 = valid ? global_state : global_state;
	end
	// controller for eq_203.eq_203_in0
	// controller for eq_203.eq_203_in1
	// Insensitive connections
	always @(*) begin
		eq_203_in0 = valid ? 32'd1 : 32'd1;
		eq_203_in1 = valid ? global_state : global_state;
	end
	// controller for eq_205.eq_205_in0
	// controller for eq_205.eq_205_in1
	// Insensitive connections
	always @(*) begin
		eq_205_in0 = valid ? 32'd2 : 32'd2;
		eq_205_in1 = valid ? global_state : global_state;
	end
	// controller for eq_208.eq_208_in0
	// controller for eq_208.eq_208_in1
	// Insensitive connections
	always @(*) begin
		eq_208_in0 = valid ? 32'd2 : 32'd2;
		eq_208_in1 = valid ? global_state : global_state;
	end
	// controller for eq_211.eq_211_in0
	// controller for eq_211.eq_211_in1
	// Insensitive connections
	always @(*) begin
		eq_211_in0 = valid ? 32'd2 : 32'd2;
		eq_211_in1 = valid ? global_state : global_state;
	end
	// controller for eq_214.eq_214_in0
	// controller for eq_214.eq_214_in1
	// Insensitive connections
	always @(*) begin
		eq_214_in0 = valid ? 32'd2 : 32'd2;
		eq_214_in1 = valid ? global_state : global_state;
	end
	// controller for eq_216.eq_216_in0
	// controller for eq_216.eq_216_in1
	// Insensitive connections
	always @(*) begin
		eq_216_in0 = valid ? 32'd3 : 32'd3;
		eq_216_in1 = valid ? global_state : global_state;
	end
	// controller for eq_219.eq_219_in0
	// controller for eq_219.eq_219_in1
	// Insensitive connections
	always @(*) begin
		eq_219_in0 = valid ? 32'd3 : 32'd3;
		eq_219_in1 = valid ? global_state : global_state;
	end
	// controller for eq_221.eq_221_in0
	// controller for eq_221.eq_221_in1
	// Insensitive connections
	always @(*) begin
		eq_221_in0 = valid ? 32'd4 : 32'd4;
		eq_221_in1 = valid ? global_state : global_state;
	end
	// controller for eq_224.eq_224_in0
	// controller for eq_224.eq_224_in1
	// Insensitive connections
	always @(*) begin
		eq_224_in0 = valid ? 32'd4 : 32'd4;
		eq_224_in1 = valid ? global_state : global_state;
	end
	// controller for eq_226.eq_226_in0
	// controller for eq_226.eq_226_in1
	// Insensitive connections
	always @(*) begin
		eq_226_in0 = valid ? 32'd5 : 32'd5;
		eq_226_in1 = valid ? global_state : global_state;
	end
	// controller for eq_229.eq_229_in0
	// controller for eq_229.eq_229_in1
	// Insensitive connections
	always @(*) begin
		eq_229_in0 = valid ? 32'd5 : 32'd5;
		eq_229_in1 = valid ? global_state : global_state;
	end
	// controller for eq_23.eq_23_in0
	// controller for eq_23.eq_23_in1
	// Insensitive connections
	always @(*) begin
		eq_23_in0 = valid ? 32'd7 : 32'd7;
		eq_23_in1 = valid ? global_state : global_state;
	end
	// controller for eq_232.eq_232_in0
	// controller for eq_232.eq_232_in1
	// Insensitive connections
	always @(*) begin
		eq_232_in0 = valid ? 32'd6 : 32'd6;
		eq_232_in1 = valid ? global_state : global_state;
	end
	// controller for eq_235.eq_235_in0
	// controller for eq_235.eq_235_in1
	// Insensitive connections
	always @(*) begin
		eq_235_in0 = valid ? 32'd6 : 32'd6;
		eq_235_in1 = valid ? global_state : global_state;
	end
	// controller for eq_237.eq_237_in0
	// controller for eq_237.eq_237_in1
	// Insensitive connections
	always @(*) begin
		eq_237_in0 = valid ? 32'd6 : 32'd6;
		eq_237_in1 = valid ? global_state : global_state;
	end
	// controller for eq_240.eq_240_in0
	// controller for eq_240.eq_240_in1
	// Insensitive connections
	always @(*) begin
		eq_240_in0 = valid ? 32'd6 : 32'd6;
		eq_240_in1 = valid ? global_state : global_state;
	end
	// controller for eq_242.eq_242_in0
	// controller for eq_242.eq_242_in1
	// Insensitive connections
	always @(*) begin
		eq_242_in0 = valid ? 32'd7 : 32'd7;
		eq_242_in1 = valid ? global_state : global_state;
	end
	// controller for eq_245.eq_245_in0
	// controller for eq_245.eq_245_in1
	// Insensitive connections
	always @(*) begin
		eq_245_in0 = valid ? 32'd7 : 32'd7;
		eq_245_in1 = valid ? global_state : global_state;
	end
	// controller for eq_248.eq_248_in0
	// controller for eq_248.eq_248_in1
	// Insensitive connections
	always @(*) begin
		eq_248_in0 = valid ? 32'd7 : 32'd7;
		eq_248_in1 = valid ? global_state : global_state;
	end
	// controller for eq_251.eq_251_in0
	// controller for eq_251.eq_251_in1
	// Insensitive connections
	always @(*) begin
		eq_251_in0 = valid ? 32'd7 : 32'd7;
		eq_251_in1 = valid ? global_state : global_state;
	end
	// controller for eq_253.eq_253_in0
	// controller for eq_253.eq_253_in1
	// Insensitive connections
	always @(*) begin
		eq_253_in0 = valid ? 32'd8 : 32'd8;
		eq_253_in1 = valid ? global_state : global_state;
	end
	// controller for eq_256.eq_256_in0
	// controller for eq_256.eq_256_in1
	// Insensitive connections
	always @(*) begin
		eq_256_in0 = valid ? 32'd8 : 32'd8;
		eq_256_in1 = valid ? global_state : global_state;
	end
	// controller for eq_258.eq_258_in0
	// controller for eq_258.eq_258_in1
	// Insensitive connections
	always @(*) begin
		eq_258_in0 = valid ? 32'd9 : 32'd9;
		eq_258_in1 = valid ? global_state : global_state;
	end
	// controller for eq_261.eq_261_in0
	// controller for eq_261.eq_261_in1
	// Insensitive connections
	always @(*) begin
		eq_261_in0 = valid ? 32'd9 : 32'd9;
		eq_261_in1 = valid ? global_state : global_state;
	end
	// controller for eq_263.eq_263_in0
	// controller for eq_263.eq_263_in1
	// Insensitive connections
	always @(*) begin
		eq_263_in0 = valid ? 32'd0 : 32'd0;
		eq_263_in1 = valid ? global_state : global_state;
	end
	// controller for eq_265.eq_265_in0
	// controller for eq_265.eq_265_in1
	// Insensitive connections
	always @(*) begin
		eq_265_in0 = valid ? 32'd0 : 32'd0;
		eq_265_in1 = valid ? global_state : global_state;
	end
	// controller for eq_267.eq_267_in0
	// controller for eq_267.eq_267_in1
	// Insensitive connections
	always @(*) begin
		eq_267_in0 = valid ? 32'd0 : 32'd0;
		eq_267_in1 = valid ? global_state : global_state;
	end
	// controller for eq_269.eq_269_in0
	// controller for eq_269.eq_269_in1
	// Insensitive connections
	always @(*) begin
		eq_269_in0 = valid ? 32'd1 : 32'd1;
		eq_269_in1 = valid ? global_state : global_state;
	end
	// controller for eq_271.eq_271_in0
	// controller for eq_271.eq_271_in1
	// Insensitive connections
	always @(*) begin
		eq_271_in0 = valid ? 32'd1 : 32'd1;
		eq_271_in1 = valid ? global_state : global_state;
	end
	// controller for eq_273.eq_273_in0
	// controller for eq_273.eq_273_in1
	// Insensitive connections
	always @(*) begin
		eq_273_in0 = valid ? 32'd1 : 32'd1;
		eq_273_in1 = valid ? global_state : global_state;
	end
	// controller for eq_275.eq_275_in0
	// controller for eq_275.eq_275_in1
	// Insensitive connections
	always @(*) begin
		eq_275_in0 = valid ? 32'd1 : 32'd1;
		eq_275_in1 = valid ? global_state : global_state;
	end
	// controller for eq_278.eq_278_in0
	// controller for eq_278.eq_278_in1
	// Insensitive connections
	always @(*) begin
		eq_278_in0 = valid ? 32'd1 : 32'd1;
		eq_278_in1 = valid ? global_state : global_state;
	end
	// controller for eq_280.eq_280_in0
	// controller for eq_280.eq_280_in1
	// Insensitive connections
	always @(*) begin
		eq_280_in0 = valid ? 32'd1 : 32'd1;
		eq_280_in1 = valid ? global_state : global_state;
	end
	// controller for eq_282.eq_282_in0
	// controller for eq_282.eq_282_in1
	// Insensitive connections
	always @(*) begin
		eq_282_in0 = valid ? 32'd2 : 32'd2;
		eq_282_in1 = valid ? global_state : global_state;
	end
	// controller for eq_284.eq_284_in0
	// controller for eq_284.eq_284_in1
	// Insensitive connections
	always @(*) begin
		eq_284_in0 = valid ? 32'd2 : 32'd2;
		eq_284_in1 = valid ? global_state : global_state;
	end
	// controller for eq_286.eq_286_in0
	// controller for eq_286.eq_286_in1
	// Insensitive connections
	always @(*) begin
		eq_286_in0 = valid ? 32'd3 : 32'd3;
		eq_286_in1 = valid ? global_state : global_state;
	end
	// controller for eq_288.eq_288_in0
	// controller for eq_288.eq_288_in1
	// Insensitive connections
	always @(*) begin
		eq_288_in0 = valid ? 32'd4 : 32'd4;
		eq_288_in1 = valid ? global_state : global_state;
	end
	// controller for eq_290.eq_290_in0
	// controller for eq_290.eq_290_in1
	// Insensitive connections
	always @(*) begin
		eq_290_in0 = valid ? 32'd4 : 32'd4;
		eq_290_in1 = valid ? global_state : global_state;
	end
	// controller for eq_292.eq_292_in0
	// controller for eq_292.eq_292_in1
	// Insensitive connections
	always @(*) begin
		eq_292_in0 = valid ? 32'd4 : 32'd4;
		eq_292_in1 = valid ? global_state : global_state;
	end
	// controller for eq_295.eq_295_in0
	// controller for eq_295.eq_295_in1
	// Insensitive connections
	always @(*) begin
		eq_295_in0 = valid ? 32'd5 : 32'd5;
		eq_295_in1 = valid ? global_state : global_state;
	end
	// controller for eq_297.eq_297_in0
	// controller for eq_297.eq_297_in1
	// Insensitive connections
	always @(*) begin
		eq_297_in0 = valid ? 32'd5 : 32'd5;
		eq_297_in1 = valid ? global_state : global_state;
	end
	// controller for eq_299.eq_299_in0
	// controller for eq_299.eq_299_in1
	// Insensitive connections
	always @(*) begin
		eq_299_in0 = valid ? 32'd5 : 32'd5;
		eq_299_in1 = valid ? global_state : global_state;
	end
	// controller for eq_30.eq_30_in0
	// controller for eq_30.eq_30_in1
	// Insensitive connections
	always @(*) begin
		eq_30_in0 = valid ? 32'd8 : 32'd8;
		eq_30_in1 = valid ? global_state : global_state;
	end
	// controller for eq_301.eq_301_in0
	// controller for eq_301.eq_301_in1
	// Insensitive connections
	always @(*) begin
		eq_301_in0 = valid ? 32'd5 : 32'd5;
		eq_301_in1 = valid ? global_state : global_state;
	end
	// controller for eq_304.eq_304_in0
	// controller for eq_304.eq_304_in1
	// Insensitive connections
	always @(*) begin
		eq_304_in0 = valid ? 32'd5 : 32'd5;
		eq_304_in1 = valid ? global_state : global_state;
	end
	// controller for eq_306.eq_306_in0
	// controller for eq_306.eq_306_in1
	// Insensitive connections
	always @(*) begin
		eq_306_in0 = valid ? 32'd5 : 32'd5;
		eq_306_in1 = valid ? global_state : global_state;
	end
	// controller for eq_309.eq_309_in0
	// controller for eq_309.eq_309_in1
	// Insensitive connections
	always @(*) begin
		eq_309_in0 = valid ? 32'd6 : 32'd6;
		eq_309_in1 = valid ? global_state : global_state;
	end
	// controller for eq_311.eq_311_in0
	// controller for eq_311.eq_311_in1
	// Insensitive connections
	always @(*) begin
		eq_311_in0 = valid ? 32'd6 : 32'd6;
		eq_311_in1 = valid ? global_state : global_state;
	end
	// controller for eq_313.eq_313_in0
	// controller for eq_313.eq_313_in1
	// Insensitive connections
	always @(*) begin
		eq_313_in0 = valid ? 32'd6 : 32'd6;
		eq_313_in1 = valid ? global_state : global_state;
	end
	// controller for eq_315.eq_315_in0
	// controller for eq_315.eq_315_in1
	// Insensitive connections
	always @(*) begin
		eq_315_in0 = valid ? 32'd6 : 32'd6;
		eq_315_in1 = valid ? global_state : global_state;
	end
	// controller for eq_317.eq_317_in0
	// controller for eq_317.eq_317_in1
	// Insensitive connections
	always @(*) begin
		eq_317_in0 = valid ? 32'd7 : 32'd7;
		eq_317_in1 = valid ? global_state : global_state;
	end
	// controller for eq_319.eq_319_in0
	// controller for eq_319.eq_319_in1
	// Insensitive connections
	always @(*) begin
		eq_319_in0 = valid ? 32'd7 : 32'd7;
		eq_319_in1 = valid ? global_state : global_state;
	end
	// controller for eq_321.eq_321_in0
	// controller for eq_321.eq_321_in1
	// Insensitive connections
	always @(*) begin
		eq_321_in0 = valid ? 32'd8 : 32'd8;
		eq_321_in1 = valid ? global_state : global_state;
	end
	// controller for eq_323.eq_323_in0
	// controller for eq_323.eq_323_in1
	// Insensitive connections
	always @(*) begin
		eq_323_in0 = valid ? 32'd8 : 32'd8;
		eq_323_in1 = valid ? global_state : global_state;
	end
	// controller for eq_325.eq_325_in0
	// controller for eq_325.eq_325_in1
	// Insensitive connections
	always @(*) begin
		eq_325_in0 = valid ? 32'd8 : 32'd8;
		eq_325_in1 = valid ? global_state : global_state;
	end
	// controller for eq_327.eq_327_in0
	// controller for eq_327.eq_327_in1
	// Insensitive connections
	always @(*) begin
		eq_327_in0 = valid ? 32'd8 : 32'd8;
		eq_327_in1 = valid ? global_state : global_state;
	end
	// controller for eq_329.eq_329_in0
	// controller for eq_329.eq_329_in1
	// Insensitive connections
	always @(*) begin
		eq_329_in0 = valid ? 32'd9 : 32'd9;
		eq_329_in1 = valid ? global_state : global_state;
	end
	// controller for eq_331.eq_331_in0
	// controller for eq_331.eq_331_in1
	// Insensitive connections
	always @(*) begin
		eq_331_in0 = valid ? 32'd9 : 32'd9;
		eq_331_in1 = valid ? global_state : global_state;
	end
	// controller for eq_34.eq_34_in0
	// controller for eq_34.eq_34_in1
	// Insensitive connections
	always @(*) begin
		eq_34_in0 = valid ? 32'd1 : 32'd1;
		eq_34_in1 = valid ? global_state : global_state;
	end
	// controller for eq_38.eq_38_in0
	// controller for eq_38.eq_38_in1
	// Insensitive connections
	always @(*) begin
		eq_38_in0 = valid ? 32'd2 : 32'd2;
		eq_38_in1 = valid ? global_state : global_state;
	end
	// controller for eq_4.eq_4_in0
	// controller for eq_4.eq_4_in1
	// Insensitive connections
	always @(*) begin
		eq_4_in0 = valid ? 32'd6 : 32'd6;
		eq_4_in1 = valid ? global_state : global_state;
	end
	// controller for eq_45.eq_45_in0
	// controller for eq_45.eq_45_in1
	// Insensitive connections
	always @(*) begin
		eq_45_in0 = valid ? 32'd4 : 32'd4;
		eq_45_in1 = valid ? global_state : global_state;
	end
	// controller for eq_49.eq_49_in0
	// controller for eq_49.eq_49_in1
	// Insensitive connections
	always @(*) begin
		eq_49_in0 = valid ? 32'd0 : 32'd0;
		eq_49_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_50.eq_50_in0
	// controller for eq_50.eq_50_in1
	// Insensitive connections
	always @(*) begin
		eq_50_in0 = valid ? 32'd1 : 32'd1;
		eq_50_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_52.eq_52_in0
	// controller for eq_52.eq_52_in1
	// Insensitive connections
	always @(*) begin
		eq_52_in0 = valid ? 32'd2 : 32'd2;
		eq_52_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_53.eq_53_in0
	// controller for eq_53.eq_53_in1
	// Insensitive connections
	always @(*) begin
		eq_53_in0 = valid ? 32'd3 : 32'd3;
		eq_53_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_55.eq_55_in0
	// controller for eq_55.eq_55_in1
	// Insensitive connections
	always @(*) begin
		eq_55_in0 = valid ? 32'd4 : 32'd4;
		eq_55_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_56.eq_56_in0
	// controller for eq_56.eq_56_in1
	// Insensitive connections
	always @(*) begin
		eq_56_in0 = valid ? 32'd5 : 32'd5;
		eq_56_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_58.eq_58_in0
	// controller for eq_58.eq_58_in1
	// Insensitive connections
	always @(*) begin
		eq_58_in0 = valid ? 32'd6 : 32'd6;
		eq_58_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_59.eq_59_in0
	// controller for eq_59.eq_59_in1
	// Insensitive connections
	always @(*) begin
		eq_59_in0 = valid ? 32'd7 : 32'd7;
		eq_59_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_60.eq_60_in0
	// controller for eq_60.eq_60_in1
	// Insensitive connections
	always @(*) begin
		eq_60_in0 = valid ? 32'd8 : 32'd8;
		eq_60_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_62.eq_62_in0
	// controller for eq_62.eq_62_in1
	// Insensitive connections
	always @(*) begin
		eq_62_in0 = valid ? 32'd9 : 32'd9;
		eq_62_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_63.eq_63_in0
	// controller for eq_63.eq_63_in1
	// Insensitive connections
	always @(*) begin
		eq_63_in0 = valid ? 32'd10 : 32'd10;
		eq_63_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_64.eq_64_in0
	// controller for eq_64.eq_64_in1
	// Insensitive connections
	always @(*) begin
		eq_64_in0 = valid ? 32'd0 : 32'd0;
		eq_64_in1 = valid ? global_state : global_state;
	end
	// controller for eq_66.eq_66_in0
	// controller for eq_66.eq_66_in1
	// Insensitive connections
	always @(*) begin
		eq_66_in0 = valid ? 32'd3 : 32'd3;
		eq_66_in1 = valid ? global_state : global_state;
	end
	// controller for eq_68.eq_68_in0
	// controller for eq_68.eq_68_in1
	// Insensitive connections
	always @(*) begin
		eq_68_in0 = valid ? 32'd5 : 32'd5;
		eq_68_in1 = valid ? global_state : global_state;
	end
	// controller for eq_70.eq_70_in0
	// controller for eq_70.eq_70_in1
	// Insensitive connections
	always @(*) begin
		eq_70_in0 = valid ? 32'd9 : 32'd9;
		eq_70_in1 = valid ? global_state : global_state;
	end
	// controller for eq_72.eq_72_in0
	// controller for eq_72.eq_72_in1
	// Insensitive connections
	always @(*) begin
		eq_72_in0 = valid ? 32'd0 : 32'd0;
		eq_72_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_73.eq_73_in0
	// controller for eq_73.eq_73_in1
	// Insensitive connections
	always @(*) begin
		eq_73_in0 = valid ? 32'd1 : 32'd1;
		eq_73_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_76.eq_76_in0
	// controller for eq_76.eq_76_in1
	// Insensitive connections
	always @(*) begin
		eq_76_in0 = valid ? 32'd2 : 32'd2;
		eq_76_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_77.eq_77_in0
	// controller for eq_77.eq_77_in1
	// Insensitive connections
	always @(*) begin
		eq_77_in0 = valid ? 32'd3 : 32'd3;
		eq_77_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_8.eq_8_in0
	// controller for eq_8.eq_8_in1
	// Insensitive connections
	always @(*) begin
		eq_8_in0 = valid ? 32'd1 : 32'd1;
		eq_8_in1 = valid ? global_state : global_state;
	end
	// controller for eq_80.eq_80_in0
	// controller for eq_80.eq_80_in1
	// Insensitive connections
	always @(*) begin
		eq_80_in0 = valid ? 32'd4 : 32'd4;
		eq_80_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_81.eq_81_in0
	// controller for eq_81.eq_81_in1
	// Insensitive connections
	always @(*) begin
		eq_81_in0 = valid ? 32'd5 : 32'd5;
		eq_81_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_84.eq_84_in0
	// controller for eq_84.eq_84_in1
	// Insensitive connections
	always @(*) begin
		eq_84_in0 = valid ? 32'd6 : 32'd6;
		eq_84_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_85.eq_85_in0
	// controller for eq_85.eq_85_in1
	// Insensitive connections
	always @(*) begin
		eq_85_in0 = valid ? 32'd7 : 32'd7;
		eq_85_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_86.eq_86_in0
	// controller for eq_86.eq_86_in1
	// Insensitive connections
	always @(*) begin
		eq_86_in0 = valid ? 32'd8 : 32'd8;
		eq_86_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_89.eq_89_in0
	// controller for eq_89.eq_89_in1
	// Insensitive connections
	always @(*) begin
		eq_89_in0 = valid ? 32'd9 : 32'd9;
		eq_89_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_90.eq_90_in0
	// controller for eq_90.eq_90_in1
	// Insensitive connections
	always @(*) begin
		eq_90_in0 = valid ? 32'd10 : 32'd10;
		eq_90_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_91.eq_91_in0
	// controller for eq_91.eq_91_in1
	// Insensitive connections
	always @(*) begin
		eq_91_in0 = valid ? 32'd0 : 32'd0;
		eq_91_in1 = valid ? global_state : global_state;
	end
	// controller for eq_93.eq_93_in0
	// controller for eq_93.eq_93_in1
	// Insensitive connections
	always @(*) begin
		eq_93_in0 = valid ? 32'd0 : 32'd0;
		eq_93_in1 = valid ? global_state : global_state;
	end
	// controller for eq_95.eq_95_in0
	// controller for eq_95.eq_95_in1
	// Insensitive connections
	always @(*) begin
		eq_95_in0 = valid ? 32'd0 : 32'd0;
		eq_95_in1 = valid ? global_state : global_state;
	end
	// controller for eq_97.eq_97_in0
	// controller for eq_97.eq_97_in1
	// Insensitive connections
	always @(*) begin
		eq_97_in0 = valid ? 32'd0 : 32'd0;
		eq_97_in1 = valid ? global_state : global_state;
	end
	// controller for eq_99.eq_99_in0
	// controller for eq_99.eq_99_in1
	// Insensitive connections
	always @(*) begin
		eq_99_in0 = valid ? 32'd5 : 32'd5;
		eq_99_in1 = valid ? global_state : global_state;
	end
	// controller for icmp_17.cmp_in0_icmp_17
	// controller for icmp_17.cmp_in1_icmp_17
	// Insensitive connections
	always @(*) begin
		cmp_in0_icmp_17 = valid ? add_out_add_16 : add_out_add_16;
		cmp_in1_icmp_17 = valid ? (32'd4) : (32'd4);
	end
	// controller for in.in_read_valid_reg
	always @(*) begin
		if (andOp_110_out) begin 
			in_read_valid_reg = -(1'd1);
		end else begin
			in_read_valid_reg = 0;
		end
	end
	// controller for notOp_11.notOp_11_in0
	// Insensitive connections
	always @(*) begin
		notOp_11_in0 = valid ? andOp_10_out : andOp_10_out;
	end
	// controller for notOp_133.notOp_133_in0
	// Insensitive connections
	always @(*) begin
		notOp_133_in0 = valid ? andOp_132_out : andOp_132_out;
	end
	// controller for notOp_139.notOp_139_in0
	// Insensitive connections
	always @(*) begin
		notOp_139_in0 = valid ? andOp_138_out : andOp_138_out;
	end
	// controller for notOp_145.notOp_145_in0
	// Insensitive connections
	always @(*) begin
		notOp_145_in0 = valid ? andOp_144_out : andOp_144_out;
	end
	// controller for notOp_15.notOp_15_in0
	// Insensitive connections
	always @(*) begin
		notOp_15_in0 = valid ? andOp_14_out : andOp_14_out;
	end
	// controller for notOp_151.notOp_151_in0
	// Insensitive connections
	always @(*) begin
		notOp_151_in0 = valid ? andOp_150_out : andOp_150_out;
	end
	// controller for notOp_157.notOp_157_in0
	// Insensitive connections
	always @(*) begin
		notOp_157_in0 = valid ? andOp_156_out : andOp_156_out;
	end
	// controller for notOp_163.notOp_163_in0
	// Insensitive connections
	always @(*) begin
		notOp_163_in0 = valid ? andOp_162_out : andOp_162_out;
	end
	// controller for notOp_167.notOp_167_in0
	// Insensitive connections
	always @(*) begin
		notOp_167_in0 = valid ? andOp_166_out : andOp_166_out;
	end
	// controller for notOp_17.notOp_17_in0
	// Insensitive connections
	always @(*) begin
		notOp_17_in0 = valid ? icmp_tmp_6 : icmp_tmp_6;
	end
	// controller for notOp_173.notOp_173_in0
	// Insensitive connections
	always @(*) begin
		notOp_173_in0 = valid ? andOp_172_out : andOp_172_out;
	end
	// controller for notOp_179.notOp_179_in0
	// Insensitive connections
	always @(*) begin
		notOp_179_in0 = valid ? andOp_178_out : andOp_178_out;
	end
	// controller for notOp_185.notOp_185_in0
	// Insensitive connections
	always @(*) begin
		notOp_185_in0 = valid ? andOp_184_out : andOp_184_out;
	end
	// controller for notOp_191.notOp_191_in0
	// Insensitive connections
	always @(*) begin
		notOp_191_in0 = valid ? andOp_190_out : andOp_190_out;
	end
	// controller for notOp_210.notOp_210_in0
	// Insensitive connections
	always @(*) begin
		notOp_210_in0 = valid ? in_read_ready : in_read_ready;
	end
	// controller for notOp_22.notOp_22_in0
	// Insensitive connections
	always @(*) begin
		notOp_22_in0 = valid ? andOp_21_out : andOp_21_out;
	end
	// controller for notOp_231.notOp_231_in0
	// Insensitive connections
	always @(*) begin
		notOp_231_in0 = valid ? icmp_tmp_6 : icmp_tmp_6;
	end
	// controller for notOp_247.notOp_247_in0
	// Insensitive connections
	always @(*) begin
		notOp_247_in0 = valid ? out_write_ready : out_write_ready;
	end
	// controller for notOp_26.notOp_26_in0
	// Insensitive connections
	always @(*) begin
		notOp_26_in0 = valid ? andOp_25_out : andOp_25_out;
	end
	// controller for notOp_28.notOp_28_in0
	// Insensitive connections
	always @(*) begin
		notOp_28_in0 = valid ? out_write_ready : out_write_ready;
	end
	// controller for notOp_3.notOp_3_in0
	// Insensitive connections
	always @(*) begin
		notOp_3_in0 = valid ? andOp_2_out : andOp_2_out;
	end
	// controller for notOp_33.notOp_33_in0
	// Insensitive connections
	always @(*) begin
		notOp_33_in0 = valid ? andOp_32_out : andOp_32_out;
	end
	// controller for notOp_37.notOp_37_in0
	// Insensitive connections
	always @(*) begin
		notOp_37_in0 = valid ? andOp_36_out : andOp_36_out;
	end
	// controller for notOp_41.notOp_41_in0
	// Insensitive connections
	always @(*) begin
		notOp_41_in0 = valid ? andOp_40_out : andOp_40_out;
	end
	// controller for notOp_43.notOp_43_in0
	// Insensitive connections
	always @(*) begin
		notOp_43_in0 = valid ? in_read_ready : in_read_ready;
	end
	// controller for notOp_48.notOp_48_in0
	// Insensitive connections
	always @(*) begin
		notOp_48_in0 = valid ? andOp_47_out : andOp_47_out;
	end
	// controller for notOp_7.notOp_7_in0
	// Insensitive connections
	always @(*) begin
		notOp_7_in0 = valid ? andOp_6_out : andOp_6_out;
	end
	// controller for notOp_74.notOp_74_in0
	// Insensitive connections
	always @(*) begin
		notOp_74_in0 = valid ? eq_73_out : eq_73_out;
	end
	// controller for notOp_78.notOp_78_in0
	// Insensitive connections
	always @(*) begin
		notOp_78_in0 = valid ? eq_77_out : eq_77_out;
	end
	// controller for notOp_82.notOp_82_in0
	// Insensitive connections
	always @(*) begin
		notOp_82_in0 = valid ? eq_81_out : eq_81_out;
	end
	// controller for notOp_87.notOp_87_in0
	// Insensitive connections
	always @(*) begin
		notOp_87_in0 = valid ? eq_86_out : eq_86_out;
	end
	// controller for orOp_51.orOp_51_in0
	// controller for orOp_51.orOp_51_in1
	// Insensitive connections
	always @(*) begin
		orOp_51_in0 = valid ? eq_50_out : eq_50_out;
		orOp_51_in1 = valid ? andOp_16_out : andOp_16_out;
	end
	// controller for orOp_54.orOp_54_in0
	// controller for orOp_54.orOp_54_in1
	// Insensitive connections
	always @(*) begin
		orOp_54_in0 = valid ? eq_53_out : eq_53_out;
		orOp_54_in1 = valid ? andOp_2_out : andOp_2_out;
	end
	// controller for orOp_57.orOp_57_in0
	// controller for orOp_57.orOp_57_in1
	// Insensitive connections
	always @(*) begin
		orOp_57_in0 = valid ? eq_56_out : eq_56_out;
		orOp_57_in1 = valid ? andOp_6_out : andOp_6_out;
	end
	// controller for orOp_61.orOp_61_in0
	// controller for orOp_61.orOp_61_in1
	// Insensitive connections
	always @(*) begin
		orOp_61_in0 = valid ? eq_60_out : eq_60_out;
		orOp_61_in1 = valid ? andOp_10_out : andOp_10_out;
	end
	// controller for out.out_in_data_reg
	always @(*) begin
		if (andOp_124_out) begin 
			out_in_data_reg = rdata_ram_0;
		end else begin
			out_in_data_reg = 0;
		end
	end
	// controller for out.out_write_valid_reg
	always @(*) begin
		if (andOp_122_out) begin 
			out_write_valid_reg = -(1'd1);
		end else begin
			out_write_valid_reg = 0;
		end
	end
	// controller for phi_5.phi_in_phi_5
	// controller for phi_5.phi_last_block_phi_5
	// controller for phi_5.phi_s_phi_5
	// Insensitive connections
	always @(*) begin
		phi_in_phi_5 = valid ? {(32'd0), add_tmp_5} : {(32'd0), add_tmp_5};
		phi_last_block_phi_5 = valid ? bb_3_predecessor_out_data : bb_3_predecessor_out_data;
		phi_s_phi_5 = valid ? {32'd0, 32'd4} : {32'd0, 32'd4};
	end
	// controller for ram_0.raddr_ram_0_reg
	always @(*) begin
		if (andOp_100_out) begin 
			raddr_ram_0_reg = 0;
		end else if (andOp_104_out) begin 
			raddr_ram_0_reg = 0;
		end else begin
			raddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.waddr_ram_0_reg
	always @(*) begin
		if (andOp_102_out) begin 
			waddr_ram_0_reg = 0;
		end else if (andOp_98_out) begin 
			waddr_ram_0_reg = 0;
		end else begin
			waddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wdata_ram_0_reg
	always @(*) begin
		if (andOp_102_out) begin 
			wdata_ram_0_reg = add_out_add_14;
		end else if (andOp_98_out) begin 
			wdata_ram_0_reg = (32'd0);
		end else begin
			wdata_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wen_ram_0_reg
	always @(*) begin
		if (andOp_102_out) begin 
			wen_ram_0_reg = 1;
		end else if (andOp_98_out) begin 
			wen_ram_0_reg = 1;
		end else begin
			wen_ram_0_reg = 0;
		end
	end
	// controller for ret_28.valid_reg
	always @(*) begin
		if (andOp_128_out) begin 
			valid_reg = 1;
		end else begin
			valid_reg = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			add_tmp_5 <= 0;
		end else begin
			if (andOp_303_out) begin
				add_tmp_5 <= add_out_add_16;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			call_tmp_2 <= 0;
		end else begin
			if (andOp_294_out) begin
				call_tmp_2 <= in_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_next_block <= 0;
		end else begin
			if (andOp_18_out) begin
				global_next_block <= 3;
			end
			if (andOp_27_out) begin
				global_next_block <= 7;
			end
			if (andOp_29_out) begin
				global_next_block <= 6;
			end
			if (andOp_42_out) begin
				global_next_block <= 10;
			end
			if (andOp_44_out) begin
				global_next_block <= 9;
			end
			if (andOp_65_out) begin
				global_next_block <= 0;
			end
			if (andOp_67_out) begin
				global_next_block <= 10;
			end
			if (andOp_69_out) begin
				global_next_block <= 4;
			end
			if (andOp_71_out) begin
				global_next_block <= 2;
			end
			if (br_10_happened_out_data) begin
				global_next_block <= 4;
			end
			if (br_5_happened_out_data) begin
				global_next_block <= 6;
			end
			if (br_7_happened_out_data) begin
				global_next_block <= 2;
			end
			if (br_8_happened_out_data) begin
				global_next_block <= 9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_199_out) begin
				global_state <= 1;
			end
			if (andOp_204_out) begin
				global_state <= 2;
			end
			if (andOp_209_out) begin
				global_state <= 3;
			end
			if (andOp_215_out) begin
				global_state <= 2;
			end
			if (andOp_220_out) begin
				global_state <= 4;
			end
			if (andOp_225_out) begin
				global_state <= 5;
			end
			if (andOp_230_out) begin
				global_state <= 6;
			end
			if (andOp_236_out) begin
				global_state <= 1;
			end
			if (andOp_241_out) begin
				global_state <= 7;
			end
			if (andOp_246_out) begin
				global_state <= 8;
			end
			if (andOp_252_out) begin
				global_state <= 7;
			end
			if (andOp_257_out) begin
				global_state <= 9;
			end
			if (andOp_262_out) begin
				global_state <= 9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			icmp_tmp_6 <= 0;
		end else begin
			if (andOp_308_out) begin
				icmp_tmp_6 <= cmp_out_icmp_17;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			last_BB_reg <= 0;
		end else begin
			if (andOp_134_out) begin
				last_BB_reg <= 0;
			end
			if (andOp_140_out) begin
				last_BB_reg <= 3;
			end
			if (andOp_146_out) begin
				last_BB_reg <= 8;
			end
			if (andOp_152_out) begin
				last_BB_reg <= 9;
			end
			if (andOp_158_out) begin
				last_BB_reg <= 10;
			end
			if (andOp_168_out) begin
				last_BB_reg <= 4;
			end
			if (andOp_174_out) begin
				last_BB_reg <= 1;
			end
			if (andOp_180_out) begin
				last_BB_reg <= 5;
			end
			if (andOp_186_out) begin
				last_BB_reg <= 6;
			end
			if (andOp_192_out) begin
				last_BB_reg <= 7;
			end
			if (andOp_194_out) begin
				last_BB_reg <= 2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			phi_tmp_0 <= 0;
		end else begin
			if (andOp_277_out) begin
				phi_tmp_0 <= phi_out_phi_5;
			end
		end
	end

endmodule

