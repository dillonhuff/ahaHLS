module vadd_smul_fifo(input [0:0] clk, input [0:0] rst, output [0:0] valid, output [31:0] arg_0_in_data, input [31:0] arg_0_out_data, input [0:0] arg_0_read_ready, output [0:0] arg_0_read_valid, input [0:0] arg_0_write_ready, output [0:0] arg_0_write_valid, output [31:0] arg_1_in_data, input [31:0] arg_1_out_data, input [0:0] arg_1_read_ready, output [0:0] arg_1_read_valid, input [0:0] arg_1_write_ready, output [0:0] arg_1_write_valid, output [31:0] arg_2_in_data, input [31:0] arg_2_out_data, input [0:0] arg_2_read_ready, output [0:0] arg_2_read_valid, input [0:0] arg_2_write_ready, output [0:0] arg_2_write_valid);

	reg [0:0] valid_reg;
	reg [31:0] arg_0_in_data_reg;
	reg [0:0] arg_0_read_valid_reg;
	reg [0:0] arg_0_write_valid_reg;
	reg [31:0] arg_1_in_data_reg;
	reg [0:0] arg_1_read_valid_reg;
	reg [0:0] arg_1_write_valid_reg;
	reg [31:0] arg_2_in_data_reg;
	reg [0:0] arg_2_read_valid_reg;
	reg [0:0] arg_2_write_valid_reg;

	assign valid = valid_reg;
	assign arg_0_in_data = arg_0_in_data_reg;
	assign arg_0_read_valid = arg_0_read_valid_reg;
	assign arg_0_write_valid = arg_0_write_valid_reg;
	assign arg_1_in_data = arg_1_in_data_reg;
	assign arg_1_read_valid = arg_1_read_valid_reg;
	assign arg_1_write_valid = arg_1_write_valid_reg;
	assign arg_2_in_data = arg_2_in_data_reg;
	assign arg_2_read_valid = arg_2_read_valid_reg;
	assign arg_2_write_valid = arg_2_write_valid_reg;

	// Start debug wires and ports

	initial begin
	end






	// End debug wires and ports

	// Start Functional Units
	reg [31:0] _____dlr_0___eq___alloca___dlr_builtin_fifo_32_in_data;
	reg [0:0] _____dlr_0___eq___alloca___dlr_builtin_fifo_32_read_valid;
	reg [0:0] _____dlr_0___eq___alloca___dlr_builtin_fifo_32_write_valid;
	wire [31:0] _____dlr_0___eq___alloca___dlr_builtin_fifo_32_out_data;
	wire [0:0] _____dlr_0___eq___alloca___dlr_builtin_fifo_32_read_ready;
	wire [0:0] _____dlr_0___eq___alloca___dlr_builtin_fifo_32_write_ready;
	fifo #(.DEPTH(16), .WIDTH(32)) _____dlr_0___eq___alloca___dlr_builtin_fifo_32(.clk(clk), .in_data(_____dlr_0___eq___alloca___dlr_builtin_fifo_32_in_data), .out_data(_____dlr_0___eq___alloca___dlr_builtin_fifo_32_out_data), .read_ready(_____dlr_0___eq___alloca___dlr_builtin_fifo_32_read_ready), .read_valid(_____dlr_0___eq___alloca___dlr_builtin_fifo_32_read_valid), .rst(rst), .write_ready(_____dlr_0___eq___alloca___dlr_builtin_fifo_32_write_ready), .write_valid(_____dlr_0___eq___alloca___dlr_builtin_fifo_32_write_valid));

	br_dummy br_unit();

	wire [31:0] add_add22_in0;
	wire [31:0] add_add22_in1;
	wire [31:0] add_add22_out;
	add #(.WIDTH(32)) add_add22(.in0(add_add22_in0), .in1(add_add22_in1), .out(add_add22_out));

	wire [31:0] icmp_icmp26_in0;
	wire [31:0] icmp_icmp26_in1;
	wire [0:0] icmp_icmp26_out;
	ne #(.WIDTH(32)) icmp_icmp26(.in0(icmp_icmp26_in0), .in1(icmp_icmp26_in1), .out(icmp_icmp26_out));

	wire [63:0] phi_phi31_in;
	wire [31:0] phi_phi31_last_block;
	wire [63:0] phi_phi31_s;
	wire [31:0] phi_phi31_out;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_phi31(.in(phi_phi31_in), .last_block(phi_phi31_last_block), .out(phi_phi31_out), .s(phi_phi31_s));

	wire [31:0] add_add32_in0;
	wire [31:0] add_add32_in1;
	wire [31:0] add_add32_out;
	add #(.WIDTH(32)) add_add32(.in0(add_add32_in0), .in1(add_add32_in1), .out(add_add32_out));

	wire [31:0] mul_mul41_in0;
	wire [31:0] mul_mul41_in1;
	wire [31:0] mul_mul41_out;
	mul #(.WIDTH(32)) mul_mul41(.in0(mul_mul41_in0), .in1(mul_mul41_in1), .out(mul_mul41_out));

	wire [31:0] icmp_icmp45_in0;
	wire [31:0] icmp_icmp45_in1;
	wire [0:0] icmp_icmp45_out;
	ne #(.WIDTH(32)) icmp_icmp45(.in0(icmp_icmp45_in0), .in1(icmp_icmp45_in1), .out(icmp_icmp45_out));

	wire [63:0] phi_phi6_in;
	wire [31:0] phi_phi6_last_block;
	wire [63:0] phi_phi6_s;
	wire [31:0] phi_phi6_out;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_phi6(.in(phi_phi6_in), .last_block(phi_phi6_last_block), .out(phi_phi6_out), .s(phi_phi6_s));

	wire [31:0] add_add7_in0;
	wire [31:0] add_add7_in1;
	wire [31:0] add_add7_out;
	add #(.WIDTH(32)) add_add7(.in0(add_add7_in0), .in1(add_add7_in1), .out(add_add7_out));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] bb_16_active_in_state_1_in_data;
	wire [0:0] bb_16_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_16_active_in_state_1(.in_data(bb_16_active_in_state_1_in_data), .out_data(bb_16_active_in_state_1_out_data));

	reg [31:0] bb_16_predecessor_in_state_1_in_data;
	wire [31:0] bb_16_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_16_predecessor_in_state_1(.in_data(bb_16_predecessor_in_state_1_in_data), .out_data(bb_16_predecessor_in_state_1_out_data));

	reg [0:0] br_16_happened_in_state_1_in_data;
	wire [0:0] br_16_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_16_happened_in_state_1(.in_data(br_16_happened_in_state_1_in_data), .out_data(br_16_happened_in_state_1_out_data));

	reg [0:0] bb_15_active_in_state_1_in_data;
	wire [0:0] bb_15_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_15_active_in_state_1(.in_data(bb_15_active_in_state_1_in_data), .out_data(bb_15_active_in_state_1_out_data));

	reg [31:0] bb_15_predecessor_in_state_1_in_data;
	wire [31:0] bb_15_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_15_predecessor_in_state_1(.in_data(bb_15_predecessor_in_state_1_in_data), .out_data(bb_15_predecessor_in_state_1_out_data));

	reg [0:0] br_15_happened_in_state_1_in_data;
	wire [0:0] br_15_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_15_happened_in_state_1(.in_data(br_15_happened_in_state_1_in_data), .out_data(br_15_happened_in_state_1_out_data));

	reg [0:0] bb_4_active_in_state_1_in_data;
	wire [0:0] bb_4_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_1(.in_data(bb_4_active_in_state_1_in_data), .out_data(bb_4_active_in_state_1_out_data));

	reg [31:0] bb_4_predecessor_in_state_1_in_data;
	wire [31:0] bb_4_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_1(.in_data(bb_4_predecessor_in_state_1_in_data), .out_data(bb_4_predecessor_in_state_1_out_data));

	reg [0:0] br_4_happened_in_state_1_in_data;
	wire [0:0] br_4_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_1(.in_data(br_4_happened_in_state_1_in_data), .out_data(br_4_happened_in_state_1_out_data));

	reg [0:0] bb_17_active_in_state_2_in_data;
	wire [0:0] bb_17_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_17_active_in_state_2(.in_data(bb_17_active_in_state_2_in_data), .out_data(bb_17_active_in_state_2_out_data));

	reg [31:0] bb_17_predecessor_in_state_2_in_data;
	wire [31:0] bb_17_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_17_predecessor_in_state_2(.in_data(bb_17_predecessor_in_state_2_in_data), .out_data(bb_17_predecessor_in_state_2_out_data));

	reg [0:0] br_17_happened_in_state_2_in_data;
	wire [0:0] br_17_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_17_happened_in_state_2(.in_data(br_17_happened_in_state_2_in_data), .out_data(br_17_happened_in_state_2_out_data));

	reg [0:0] bb_18_active_in_state_3_in_data;
	wire [0:0] bb_18_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_18_active_in_state_3(.in_data(bb_18_active_in_state_3_in_data), .out_data(bb_18_active_in_state_3_out_data));

	reg [31:0] bb_18_predecessor_in_state_3_in_data;
	wire [31:0] bb_18_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_18_predecessor_in_state_3(.in_data(bb_18_predecessor_in_state_3_in_data), .out_data(bb_18_predecessor_in_state_3_out_data));

	reg [0:0] br_18_happened_in_state_3_in_data;
	wire [0:0] br_18_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_18_happened_in_state_3(.in_data(br_18_happened_in_state_3_in_data), .out_data(br_18_happened_in_state_3_out_data));

	reg [0:0] bb_17_active_in_state_3_in_data;
	wire [0:0] bb_17_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_17_active_in_state_3(.in_data(bb_17_active_in_state_3_in_data), .out_data(bb_17_active_in_state_3_out_data));

	reg [31:0] bb_17_predecessor_in_state_3_in_data;
	wire [31:0] bb_17_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_17_predecessor_in_state_3(.in_data(bb_17_predecessor_in_state_3_in_data), .out_data(bb_17_predecessor_in_state_3_out_data));

	reg [0:0] br_17_happened_in_state_3_in_data;
	wire [0:0] br_17_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_17_happened_in_state_3(.in_data(br_17_happened_in_state_3_in_data), .out_data(br_17_happened_in_state_3_out_data));

	reg [0:0] bb_5_active_in_state_3_in_data;
	wire [0:0] bb_5_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_5_active_in_state_3(.in_data(bb_5_active_in_state_3_in_data), .out_data(bb_5_active_in_state_3_out_data));

	reg [31:0] bb_5_predecessor_in_state_3_in_data;
	wire [31:0] bb_5_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_5_predecessor_in_state_3(.in_data(bb_5_predecessor_in_state_3_in_data), .out_data(bb_5_predecessor_in_state_3_out_data));

	reg [0:0] br_5_happened_in_state_3_in_data;
	wire [0:0] br_5_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_5_happened_in_state_3(.in_data(br_5_happened_in_state_3_in_data), .out_data(br_5_happened_in_state_3_out_data));

	reg [0:0] bb_19_active_in_state_3_in_data;
	wire [0:0] bb_19_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_19_active_in_state_3(.in_data(bb_19_active_in_state_3_in_data), .out_data(bb_19_active_in_state_3_out_data));

	reg [31:0] bb_19_predecessor_in_state_3_in_data;
	wire [31:0] bb_19_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_19_predecessor_in_state_3(.in_data(bb_19_predecessor_in_state_3_in_data), .out_data(bb_19_predecessor_in_state_3_out_data));

	reg [0:0] br_19_happened_in_state_3_in_data;
	wire [0:0] br_19_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_19_happened_in_state_3(.in_data(br_19_happened_in_state_3_in_data), .out_data(br_19_happened_in_state_3_out_data));

	reg [0:0] bb_20_active_in_state_4_in_data;
	wire [0:0] bb_20_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_20_active_in_state_4(.in_data(bb_20_active_in_state_4_in_data), .out_data(bb_20_active_in_state_4_out_data));

	reg [31:0] bb_20_predecessor_in_state_4_in_data;
	wire [31:0] bb_20_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_20_predecessor_in_state_4(.in_data(bb_20_predecessor_in_state_4_in_data), .out_data(bb_20_predecessor_in_state_4_out_data));

	reg [0:0] br_20_happened_in_state_4_in_data;
	wire [0:0] br_20_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_20_happened_in_state_4(.in_data(br_20_happened_in_state_4_in_data), .out_data(br_20_happened_in_state_4_out_data));

	reg [0:0] bb_20_active_in_state_5_in_data;
	wire [0:0] bb_20_active_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) bb_20_active_in_state_5(.in_data(bb_20_active_in_state_5_in_data), .out_data(bb_20_active_in_state_5_out_data));

	reg [31:0] bb_20_predecessor_in_state_5_in_data;
	wire [31:0] bb_20_predecessor_in_state_5_out_data;
	hls_wire #(.WIDTH(32)) bb_20_predecessor_in_state_5(.in_data(bb_20_predecessor_in_state_5_in_data), .out_data(bb_20_predecessor_in_state_5_out_data));

	reg [0:0] br_20_happened_in_state_5_in_data;
	wire [0:0] br_20_happened_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) br_20_happened_in_state_5(.in_data(br_20_happened_in_state_5_in_data), .out_data(br_20_happened_in_state_5_out_data));

	reg [0:0] bb_21_active_in_state_6_in_data;
	wire [0:0] bb_21_active_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) bb_21_active_in_state_6(.in_data(bb_21_active_in_state_6_in_data), .out_data(bb_21_active_in_state_6_out_data));

	reg [31:0] bb_21_predecessor_in_state_6_in_data;
	wire [31:0] bb_21_predecessor_in_state_6_out_data;
	hls_wire #(.WIDTH(32)) bb_21_predecessor_in_state_6(.in_data(bb_21_predecessor_in_state_6_in_data), .out_data(bb_21_predecessor_in_state_6_out_data));

	reg [0:0] br_21_happened_in_state_6_in_data;
	wire [0:0] br_21_happened_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) br_21_happened_in_state_6(.in_data(br_21_happened_in_state_6_in_data), .out_data(br_21_happened_in_state_6_out_data));

	reg [0:0] bb_6_active_in_state_6_in_data;
	wire [0:0] bb_6_active_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) bb_6_active_in_state_6(.in_data(bb_6_active_in_state_6_in_data), .out_data(bb_6_active_in_state_6_out_data));

	reg [31:0] bb_6_predecessor_in_state_6_in_data;
	wire [31:0] bb_6_predecessor_in_state_6_out_data;
	hls_wire #(.WIDTH(32)) bb_6_predecessor_in_state_6(.in_data(bb_6_predecessor_in_state_6_in_data), .out_data(bb_6_predecessor_in_state_6_out_data));

	reg [0:0] br_6_happened_in_state_6_in_data;
	wire [0:0] br_6_happened_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) br_6_happened_in_state_6(.in_data(br_6_happened_in_state_6_in_data), .out_data(br_6_happened_in_state_6_out_data));

	reg [0:0] bb_20_active_in_state_6_in_data;
	wire [0:0] bb_20_active_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) bb_20_active_in_state_6(.in_data(bb_20_active_in_state_6_in_data), .out_data(bb_20_active_in_state_6_out_data));

	reg [31:0] bb_20_predecessor_in_state_6_in_data;
	wire [31:0] bb_20_predecessor_in_state_6_out_data;
	hls_wire #(.WIDTH(32)) bb_20_predecessor_in_state_6(.in_data(bb_20_predecessor_in_state_6_in_data), .out_data(bb_20_predecessor_in_state_6_out_data));

	reg [0:0] br_20_happened_in_state_6_in_data;
	wire [0:0] br_20_happened_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) br_20_happened_in_state_6(.in_data(br_20_happened_in_state_6_in_data), .out_data(br_20_happened_in_state_6_out_data));

	reg [0:0] bb_22_active_in_state_6_in_data;
	wire [0:0] bb_22_active_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) bb_22_active_in_state_6(.in_data(bb_22_active_in_state_6_in_data), .out_data(bb_22_active_in_state_6_out_data));

	reg [31:0] bb_22_predecessor_in_state_6_in_data;
	wire [31:0] bb_22_predecessor_in_state_6_out_data;
	hls_wire #(.WIDTH(32)) bb_22_predecessor_in_state_6(.in_data(bb_22_predecessor_in_state_6_in_data), .out_data(bb_22_predecessor_in_state_6_out_data));

	reg [0:0] br_22_happened_in_state_6_in_data;
	wire [0:0] br_22_happened_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) br_22_happened_in_state_6(.in_data(br_22_happened_in_state_6_in_data), .out_data(br_22_happened_in_state_6_out_data));

	reg [0:0] bb_7_active_in_state_7_in_data;
	wire [0:0] bb_7_active_in_state_7_out_data;
	hls_wire #(.WIDTH(1)) bb_7_active_in_state_7(.in_data(bb_7_active_in_state_7_in_data), .out_data(bb_7_active_in_state_7_out_data));

	reg [31:0] bb_7_predecessor_in_state_7_in_data;
	wire [31:0] bb_7_predecessor_in_state_7_out_data;
	hls_wire #(.WIDTH(32)) bb_7_predecessor_in_state_7(.in_data(bb_7_predecessor_in_state_7_in_data), .out_data(bb_7_predecessor_in_state_7_out_data));

	reg [0:0] br_7_happened_in_state_7_in_data;
	wire [0:0] br_7_happened_in_state_7_out_data;
	hls_wire #(.WIDTH(1)) br_7_happened_in_state_7(.in_data(br_7_happened_in_state_7_in_data), .out_data(br_7_happened_in_state_7_out_data));

	reg [0:0] bb_23_active_in_state_7_in_data;
	wire [0:0] bb_23_active_in_state_7_out_data;
	hls_wire #(.WIDTH(1)) bb_23_active_in_state_7(.in_data(bb_23_active_in_state_7_in_data), .out_data(bb_23_active_in_state_7_out_data));

	reg [31:0] bb_23_predecessor_in_state_7_in_data;
	wire [31:0] bb_23_predecessor_in_state_7_out_data;
	hls_wire #(.WIDTH(32)) bb_23_predecessor_in_state_7(.in_data(bb_23_predecessor_in_state_7_in_data), .out_data(bb_23_predecessor_in_state_7_out_data));

	reg [0:0] br_23_happened_in_state_7_in_data;
	wire [0:0] br_23_happened_in_state_7_out_data;
	hls_wire #(.WIDTH(1)) br_23_happened_in_state_7(.in_data(br_23_happened_in_state_7_in_data), .out_data(br_23_happened_in_state_7_out_data));

	reg [0:0] bb_1_active_in_state_8_in_data;
	wire [0:0] bb_1_active_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_8(.in_data(bb_1_active_in_state_8_in_data), .out_data(bb_1_active_in_state_8_out_data));

	reg [31:0] bb_1_predecessor_in_state_8_in_data;
	wire [31:0] bb_1_predecessor_in_state_8_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_8(.in_data(bb_1_predecessor_in_state_8_in_data), .out_data(bb_1_predecessor_in_state_8_out_data));

	reg [0:0] br_1_happened_in_state_8_in_data;
	wire [0:0] br_1_happened_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened_in_state_8(.in_data(br_1_happened_in_state_8_in_data), .out_data(br_1_happened_in_state_8_out_data));

	reg [0:0] bb_9_active_in_state_8_in_data;
	wire [0:0] bb_9_active_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) bb_9_active_in_state_8(.in_data(bb_9_active_in_state_8_in_data), .out_data(bb_9_active_in_state_8_out_data));

	reg [31:0] bb_9_predecessor_in_state_8_in_data;
	wire [31:0] bb_9_predecessor_in_state_8_out_data;
	hls_wire #(.WIDTH(32)) bb_9_predecessor_in_state_8(.in_data(bb_9_predecessor_in_state_8_in_data), .out_data(bb_9_predecessor_in_state_8_out_data));

	reg [0:0] br_9_happened_in_state_8_in_data;
	wire [0:0] br_9_happened_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) br_9_happened_in_state_8(.in_data(br_9_happened_in_state_8_in_data), .out_data(br_9_happened_in_state_8_out_data));

	reg [0:0] bb_10_active_in_state_8_in_data;
	wire [0:0] bb_10_active_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_8(.in_data(bb_10_active_in_state_8_in_data), .out_data(bb_10_active_in_state_8_out_data));

	reg [31:0] bb_10_predecessor_in_state_8_in_data;
	wire [31:0] bb_10_predecessor_in_state_8_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_8(.in_data(bb_10_predecessor_in_state_8_in_data), .out_data(bb_10_predecessor_in_state_8_out_data));

	reg [0:0] br_10_happened_in_state_8_in_data;
	wire [0:0] br_10_happened_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_8(.in_data(br_10_happened_in_state_8_in_data), .out_data(br_10_happened_in_state_8_out_data));

	reg [0:0] bb_11_active_in_state_9_in_data;
	wire [0:0] bb_11_active_in_state_9_out_data;
	hls_wire #(.WIDTH(1)) bb_11_active_in_state_9(.in_data(bb_11_active_in_state_9_in_data), .out_data(bb_11_active_in_state_9_out_data));

	reg [31:0] bb_11_predecessor_in_state_9_in_data;
	wire [31:0] bb_11_predecessor_in_state_9_out_data;
	hls_wire #(.WIDTH(32)) bb_11_predecessor_in_state_9(.in_data(bb_11_predecessor_in_state_9_in_data), .out_data(bb_11_predecessor_in_state_9_out_data));

	reg [0:0] br_11_happened_in_state_9_in_data;
	wire [0:0] br_11_happened_in_state_9_out_data;
	hls_wire #(.WIDTH(1)) br_11_happened_in_state_9(.in_data(br_11_happened_in_state_9_in_data), .out_data(br_11_happened_in_state_9_out_data));

	reg [0:0] bb_11_active_in_state_10_in_data;
	wire [0:0] bb_11_active_in_state_10_out_data;
	hls_wire #(.WIDTH(1)) bb_11_active_in_state_10(.in_data(bb_11_active_in_state_10_in_data), .out_data(bb_11_active_in_state_10_out_data));

	reg [31:0] bb_11_predecessor_in_state_10_in_data;
	wire [31:0] bb_11_predecessor_in_state_10_out_data;
	hls_wire #(.WIDTH(32)) bb_11_predecessor_in_state_10(.in_data(bb_11_predecessor_in_state_10_in_data), .out_data(bb_11_predecessor_in_state_10_out_data));

	reg [0:0] br_11_happened_in_state_10_in_data;
	wire [0:0] br_11_happened_in_state_10_out_data;
	hls_wire #(.WIDTH(1)) br_11_happened_in_state_10(.in_data(br_11_happened_in_state_10_in_data), .out_data(br_11_happened_in_state_10_out_data));

	reg [0:0] bb_12_active_in_state_11_in_data;
	wire [0:0] bb_12_active_in_state_11_out_data;
	hls_wire #(.WIDTH(1)) bb_12_active_in_state_11(.in_data(bb_12_active_in_state_11_in_data), .out_data(bb_12_active_in_state_11_out_data));

	reg [31:0] bb_12_predecessor_in_state_11_in_data;
	wire [31:0] bb_12_predecessor_in_state_11_out_data;
	hls_wire #(.WIDTH(32)) bb_12_predecessor_in_state_11(.in_data(bb_12_predecessor_in_state_11_in_data), .out_data(bb_12_predecessor_in_state_11_out_data));

	reg [0:0] br_12_happened_in_state_11_in_data;
	wire [0:0] br_12_happened_in_state_11_out_data;
	hls_wire #(.WIDTH(1)) br_12_happened_in_state_11(.in_data(br_12_happened_in_state_11_in_data), .out_data(br_12_happened_in_state_11_out_data));

	reg [0:0] bb_13_active_in_state_11_in_data;
	wire [0:0] bb_13_active_in_state_11_out_data;
	hls_wire #(.WIDTH(1)) bb_13_active_in_state_11(.in_data(bb_13_active_in_state_11_in_data), .out_data(bb_13_active_in_state_11_out_data));

	reg [31:0] bb_13_predecessor_in_state_11_in_data;
	wire [31:0] bb_13_predecessor_in_state_11_out_data;
	hls_wire #(.WIDTH(32)) bb_13_predecessor_in_state_11(.in_data(bb_13_predecessor_in_state_11_in_data), .out_data(bb_13_predecessor_in_state_11_out_data));

	reg [0:0] br_13_happened_in_state_11_in_data;
	wire [0:0] br_13_happened_in_state_11_out_data;
	hls_wire #(.WIDTH(1)) br_13_happened_in_state_11(.in_data(br_13_happened_in_state_11_in_data), .out_data(br_13_happened_in_state_11_out_data));

	reg [0:0] bb_2_active_in_state_11_in_data;
	wire [0:0] bb_2_active_in_state_11_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_11(.in_data(bb_2_active_in_state_11_in_data), .out_data(bb_2_active_in_state_11_out_data));

	reg [31:0] bb_2_predecessor_in_state_11_in_data;
	wire [31:0] bb_2_predecessor_in_state_11_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_11(.in_data(bb_2_predecessor_in_state_11_in_data), .out_data(bb_2_predecessor_in_state_11_out_data));

	reg [0:0] br_2_happened_in_state_11_in_data;
	wire [0:0] br_2_happened_in_state_11_out_data;
	hls_wire #(.WIDTH(1)) br_2_happened_in_state_11(.in_data(br_2_happened_in_state_11_in_data), .out_data(br_2_happened_in_state_11_out_data));

	reg [0:0] bb_3_active_in_state_12_in_data;
	wire [0:0] bb_3_active_in_state_12_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_12(.in_data(bb_3_active_in_state_12_in_data), .out_data(bb_3_active_in_state_12_out_data));

	reg [31:0] bb_3_predecessor_in_state_12_in_data;
	wire [31:0] bb_3_predecessor_in_state_12_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_12(.in_data(bb_3_predecessor_in_state_12_in_data), .out_data(bb_3_predecessor_in_state_12_out_data));

	reg [0:0] br_3_happened_in_state_12_in_data;
	wire [0:0] br_3_happened_in_state_12_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_12(.in_data(br_3_happened_in_state_12_in_data), .out_data(br_3_happened_in_state_12_out_data));

	reg [0:0] bb_14_active_in_state_12_in_data;
	wire [0:0] bb_14_active_in_state_12_out_data;
	hls_wire #(.WIDTH(1)) bb_14_active_in_state_12(.in_data(bb_14_active_in_state_12_in_data), .out_data(bb_14_active_in_state_12_out_data));

	reg [31:0] bb_14_predecessor_in_state_12_in_data;
	wire [31:0] bb_14_predecessor_in_state_12_out_data;
	hls_wire #(.WIDTH(32)) bb_14_predecessor_in_state_12(.in_data(bb_14_predecessor_in_state_12_in_data), .out_data(bb_14_predecessor_in_state_12_out_data));

	reg [0:0] br_14_happened_in_state_12_in_data;
	wire [0:0] br_14_happened_in_state_12_out_data;
	hls_wire #(.WIDTH(1)) br_14_happened_in_state_12(.in_data(br_14_happened_in_state_12_in_data), .out_data(br_14_happened_in_state_12_out_data));

	reg [0:0] bb_8_active_in_state_13_in_data;
	wire [0:0] bb_8_active_in_state_13_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active_in_state_13(.in_data(bb_8_active_in_state_13_in_data), .out_data(bb_8_active_in_state_13_out_data));

	reg [31:0] bb_8_predecessor_in_state_13_in_data;
	wire [31:0] bb_8_predecessor_in_state_13_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor_in_state_13(.in_data(bb_8_predecessor_in_state_13_in_data), .out_data(bb_8_predecessor_in_state_13_out_data));

	reg [31:0] data_in_1_1_in_data;
	wire [31:0] data_in_1_1_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_1(.in_data(data_in_1_1_in_data), .out_data(data_in_1_1_out_data));

	reg [31:0] data_in_1_3_in_data;
	wire [31:0] data_in_1_3_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_3(.in_data(data_in_1_3_in_data), .out_data(data_in_1_3_out_data));

	reg [31:0] data_in_1_5_in_data;
	wire [31:0] data_in_1_5_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_5(.in_data(data_in_1_5_in_data), .out_data(data_in_1_5_out_data));

	reg [31:0] data_in_2_7_in_data;
	wire [31:0] data_in_2_7_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_7(.in_data(data_in_2_7_in_data), .out_data(data_in_2_7_out_data));

	reg [31:0] data_in_2_9_in_data;
	wire [31:0] data_in_2_9_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_9(.in_data(data_in_2_9_in_data), .out_data(data_in_2_9_out_data));

	reg [31:0] data_in_2_11_in_data;
	wire [31:0] data_in_2_11_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_11(.in_data(data_in_2_11_in_data), .out_data(data_in_2_11_out_data));

	reg [31:0] data_in_3_13_in_data;
	wire [31:0] data_in_3_13_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_13(.in_data(data_in_3_13_in_data), .out_data(data_in_3_13_out_data));

	reg [31:0] data_in_3_15_in_data;
	wire [31:0] data_in_3_15_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_15(.in_data(data_in_3_15_in_data), .out_data(data_in_3_15_out_data));

	reg [31:0] data_in_3_17_in_data;
	wire [31:0] data_in_3_17_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_17(.in_data(data_in_3_17_in_data), .out_data(data_in_3_17_out_data));

	reg [31:0] data_in_4_19_in_data;
	wire [31:0] data_in_4_19_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_19(.in_data(data_in_4_19_in_data), .out_data(data_in_4_19_out_data));

	reg [31:0] data_in_4_21_in_data;
	wire [31:0] data_in_4_21_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_21(.in_data(data_in_4_21_in_data), .out_data(data_in_4_21_out_data));

	reg [31:0] data_in_4_23_in_data;
	wire [31:0] data_in_4_23_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_23(.in_data(data_in_4_23_in_data), .out_data(data_in_4_23_out_data));

	reg [31:0] data_in_5_26_in_data;
	wire [31:0] data_in_5_26_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_26(.in_data(data_in_5_26_in_data), .out_data(data_in_5_26_out_data));

	reg [31:0] data_in_5_28_in_data;
	wire [31:0] data_in_5_28_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_28(.in_data(data_in_5_28_in_data), .out_data(data_in_5_28_out_data));

	reg [31:0] data_in_5_30_in_data;
	wire [31:0] data_in_5_30_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_30(.in_data(data_in_5_30_in_data), .out_data(data_in_5_30_out_data));

	reg [31:0] data_in_6_32_in_data;
	wire [31:0] data_in_6_32_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_32(.in_data(data_in_6_32_in_data), .out_data(data_in_6_32_out_data));

	reg [31:0] data_in_6_34_in_data;
	wire [31:0] data_in_6_34_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_34(.in_data(data_in_6_34_in_data), .out_data(data_in_6_34_out_data));

	reg [31:0] data_in_6_36_in_data;
	wire [31:0] data_in_6_36_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_36(.in_data(data_in_6_36_in_data), .out_data(data_in_6_36_out_data));

	reg [31:0] data_in_6_38_in_data;
	wire [31:0] data_in_6_38_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_38(.in_data(data_in_6_38_in_data), .out_data(data_in_6_38_out_data));

	reg [31:0] data_in_7_40_in_data;
	wire [31:0] data_in_7_40_out_data;
	hls_wire #(.WIDTH(32)) data_in_7_40(.in_data(data_in_7_40_in_data), .out_data(data_in_7_40_out_data));

	reg [31:0] data_in_7_42_in_data;
	wire [31:0] data_in_7_42_out_data;
	hls_wire #(.WIDTH(32)) data_in_7_42(.in_data(data_in_7_42_in_data), .out_data(data_in_7_42_out_data));

	reg [31:0] data_in_7_44_in_data;
	wire [31:0] data_in_7_44_out_data;
	hls_wire #(.WIDTH(32)) data_in_7_44(.in_data(data_in_7_44_in_data), .out_data(data_in_7_44_out_data));

	reg [31:0] data_in_8_46_in_data;
	wire [31:0] data_in_8_46_out_data;
	hls_wire #(.WIDTH(32)) data_in_8_46(.in_data(data_in_8_46_in_data), .out_data(data_in_8_46_out_data));

	reg [31:0] data_in_8_48_in_data;
	wire [31:0] data_in_8_48_out_data;
	hls_wire #(.WIDTH(32)) data_in_8_48(.in_data(data_in_8_48_in_data), .out_data(data_in_8_48_out_data));

	reg [31:0] data_in_9_50_in_data;
	wire [31:0] data_in_9_50_out_data;
	hls_wire #(.WIDTH(32)) data_in_9_50(.in_data(data_in_9_50_in_data), .out_data(data_in_9_50_out_data));

	reg [31:0] data_in_9_52_in_data;
	wire [31:0] data_in_9_52_out_data;
	hls_wire #(.WIDTH(32)) data_in_9_52(.in_data(data_in_9_52_in_data), .out_data(data_in_9_52_out_data));

	reg [31:0] data_in_10_55_in_data;
	wire [31:0] data_in_10_55_out_data;
	hls_wire #(.WIDTH(32)) data_in_10_55(.in_data(data_in_10_55_in_data), .out_data(data_in_10_55_out_data));

	reg [31:0] data_in_10_57_in_data;
	wire [31:0] data_in_10_57_out_data;
	hls_wire #(.WIDTH(32)) data_in_10_57(.in_data(data_in_10_57_in_data), .out_data(data_in_10_57_out_data));

	reg [31:0] data_in_11_59_in_data;
	wire [31:0] data_in_11_59_out_data;
	hls_wire #(.WIDTH(32)) data_in_11_59(.in_data(data_in_11_59_in_data), .out_data(data_in_11_59_out_data));

	reg [31:0] data_in_11_61_in_data;
	wire [31:0] data_in_11_61_out_data;
	hls_wire #(.WIDTH(32)) data_in_11_61(.in_data(data_in_11_61_in_data), .out_data(data_in_11_61_out_data));

	reg [31:0] data_in_11_63_in_data;
	wire [31:0] data_in_11_63_out_data;
	hls_wire #(.WIDTH(32)) data_in_11_63(.in_data(data_in_11_63_in_data), .out_data(data_in_11_63_out_data));

	reg [31:0] data_in_12_65_in_data;
	wire [31:0] data_in_12_65_out_data;
	hls_wire #(.WIDTH(32)) data_in_12_65(.in_data(data_in_12_65_in_data), .out_data(data_in_12_65_out_data));

	reg [31:0] data_in_12_67_in_data;
	wire [31:0] data_in_12_67_out_data;
	hls_wire #(.WIDTH(32)) data_in_12_67(.in_data(data_in_12_67_in_data), .out_data(data_in_12_67_out_data));

	wire [0:0] andOp_68_in0;
	wire [0:0] andOp_68_in1;
	wire [0:0] andOp_68_out;
	andOp #(.WIDTH(1)) andOp_68(.in0(andOp_68_in0), .in1(andOp_68_in1), .out(andOp_68_out));

	wire [0:0] notOp_69_in0;
	wire [0:0] notOp_69_out;
	notOp #(.WIDTH(1)) notOp_69(.in(notOp_69_in0), .out(notOp_69_out));

	wire [0:0] andOp_70_in0;
	wire [0:0] andOp_70_in1;
	wire [0:0] andOp_70_out;
	andOp #(.WIDTH(1)) andOp_70(.in0(andOp_70_in0), .in1(andOp_70_in1), .out(andOp_70_out));

	wire [0:0] notOp_71_in0;
	wire [0:0] notOp_71_out;
	notOp #(.WIDTH(1)) notOp_71(.in(notOp_71_in0), .out(notOp_71_out));

	wire [0:0] andOp_72_in0;
	wire [0:0] andOp_72_in1;
	wire [0:0] andOp_72_out;
	andOp #(.WIDTH(1)) andOp_72(.in0(andOp_72_in0), .in1(andOp_72_in1), .out(andOp_72_out));

	wire [0:0] notOp_73_in0;
	wire [0:0] notOp_73_out;
	notOp #(.WIDTH(1)) notOp_73(.in(notOp_73_in0), .out(notOp_73_out));

	wire [0:0] andOp_74_in0;
	wire [0:0] andOp_74_in1;
	wire [0:0] andOp_74_out;
	andOp #(.WIDTH(1)) andOp_74(.in0(andOp_74_in0), .in1(andOp_74_in1), .out(andOp_74_out));

	wire [0:0] andOp_75_in0;
	wire [0:0] andOp_75_in1;
	wire [0:0] andOp_75_out;
	andOp #(.WIDTH(1)) andOp_75(.in0(andOp_75_in0), .in1(andOp_75_in1), .out(andOp_75_out));

	wire [0:0] notOp_76_in0;
	wire [0:0] notOp_76_out;
	notOp #(.WIDTH(1)) notOp_76(.in(notOp_76_in0), .out(notOp_76_out));

	wire [0:0] andOp_77_in0;
	wire [0:0] andOp_77_in1;
	wire [0:0] andOp_77_out;
	andOp #(.WIDTH(1)) andOp_77(.in0(andOp_77_in0), .in1(andOp_77_in1), .out(andOp_77_out));

	wire [0:0] notOp_78_in0;
	wire [0:0] notOp_78_out;
	notOp #(.WIDTH(1)) notOp_78(.in(notOp_78_in0), .out(notOp_78_out));

	wire [0:0] andOp_79_in0;
	wire [0:0] andOp_79_in1;
	wire [0:0] andOp_79_out;
	andOp #(.WIDTH(1)) andOp_79(.in0(andOp_79_in0), .in1(andOp_79_in1), .out(andOp_79_out));

	wire [0:0] notOp_80_in0;
	wire [0:0] notOp_80_out;
	notOp #(.WIDTH(1)) notOp_80(.in(notOp_80_in0), .out(notOp_80_out));

	wire [0:0] andOp_81_in0;
	wire [0:0] andOp_81_in1;
	wire [0:0] andOp_81_out;
	andOp #(.WIDTH(1)) andOp_81(.in0(andOp_81_in0), .in1(andOp_81_in1), .out(andOp_81_out));

	wire [0:0] notOp_82_in0;
	wire [0:0] notOp_82_out;
	notOp #(.WIDTH(1)) notOp_82(.in(notOp_82_in0), .out(notOp_82_out));

	wire [0:0] andOp_83_in0;
	wire [0:0] andOp_83_in1;
	wire [0:0] andOp_83_out;
	andOp #(.WIDTH(1)) andOp_83(.in0(andOp_83_in0), .in1(andOp_83_in1), .out(andOp_83_out));

	wire [0:0] notOp_84_in0;
	wire [0:0] notOp_84_out;
	notOp #(.WIDTH(1)) notOp_84(.in(notOp_84_in0), .out(notOp_84_out));

	wire [0:0] andOp_85_in0;
	wire [0:0] andOp_85_in1;
	wire [0:0] andOp_85_out;
	andOp #(.WIDTH(1)) andOp_85(.in0(andOp_85_in0), .in1(andOp_85_in1), .out(andOp_85_out));

	wire [0:0] notOp_86_in0;
	wire [0:0] notOp_86_out;
	notOp #(.WIDTH(1)) notOp_86(.in(notOp_86_in0), .out(notOp_86_out));

	wire [0:0] andOp_87_in0;
	wire [0:0] andOp_87_in1;
	wire [0:0] andOp_87_out;
	andOp #(.WIDTH(1)) andOp_87(.in0(andOp_87_in0), .in1(andOp_87_in1), .out(andOp_87_out));

	wire [0:0] notOp_88_in0;
	wire [0:0] notOp_88_out;
	notOp #(.WIDTH(1)) notOp_88(.in(notOp_88_in0), .out(notOp_88_out));

	wire [0:0] andOp_89_in0;
	wire [0:0] andOp_89_in1;
	wire [0:0] andOp_89_out;
	andOp #(.WIDTH(1)) andOp_89(.in0(andOp_89_in0), .in1(andOp_89_in1), .out(andOp_89_out));

	wire [0:0] notOp_90_in0;
	wire [0:0] notOp_90_out;
	notOp #(.WIDTH(1)) notOp_90(.in(notOp_90_in0), .out(notOp_90_out));

	wire [0:0] andOp_91_in0;
	wire [0:0] andOp_91_in1;
	wire [0:0] andOp_91_out;
	andOp #(.WIDTH(1)) andOp_91(.in0(andOp_91_in0), .in1(andOp_91_in1), .out(andOp_91_out));

	wire [0:0] andOp_92_in0;
	wire [0:0] andOp_92_in1;
	wire [0:0] andOp_92_out;
	andOp #(.WIDTH(1)) andOp_92(.in0(andOp_92_in0), .in1(andOp_92_in1), .out(andOp_92_out));

	wire [0:0] notOp_93_in0;
	wire [0:0] notOp_93_out;
	notOp #(.WIDTH(1)) notOp_93(.in(notOp_93_in0), .out(notOp_93_out));

	wire [0:0] andOp_94_in0;
	wire [0:0] andOp_94_in1;
	wire [0:0] andOp_94_out;
	andOp #(.WIDTH(1)) andOp_94(.in0(andOp_94_in0), .in1(andOp_94_in1), .out(andOp_94_out));

	wire [0:0] notOp_95_in0;
	wire [0:0] notOp_95_out;
	notOp #(.WIDTH(1)) notOp_95(.in(notOp_95_in0), .out(notOp_95_out));

	wire [0:0] andOp_96_in0;
	wire [0:0] andOp_96_in1;
	wire [0:0] andOp_96_out;
	andOp #(.WIDTH(1)) andOp_96(.in0(andOp_96_in0), .in1(andOp_96_in1), .out(andOp_96_out));

	wire [0:0] notOp_97_in0;
	wire [0:0] notOp_97_out;
	notOp #(.WIDTH(1)) notOp_97(.in(notOp_97_in0), .out(notOp_97_out));

	wire [0:0] andOp_98_in0;
	wire [0:0] andOp_98_in1;
	wire [0:0] andOp_98_out;
	andOp #(.WIDTH(1)) andOp_98(.in0(andOp_98_in0), .in1(andOp_98_in1), .out(andOp_98_out));

	wire [0:0] notOp_99_in0;
	wire [0:0] notOp_99_out;
	notOp #(.WIDTH(1)) notOp_99(.in(notOp_99_in0), .out(notOp_99_out));

	wire [0:0] andOp_100_in0;
	wire [0:0] andOp_100_in1;
	wire [0:0] andOp_100_out;
	andOp #(.WIDTH(1)) andOp_100(.in0(andOp_100_in0), .in1(andOp_100_in1), .out(andOp_100_out));

	wire [0:0] notOp_101_in0;
	wire [0:0] notOp_101_out;
	notOp #(.WIDTH(1)) notOp_101(.in(notOp_101_in0), .out(notOp_101_out));

	wire [0:0] andOp_102_in0;
	wire [0:0] andOp_102_in1;
	wire [0:0] andOp_102_out;
	andOp #(.WIDTH(1)) andOp_102(.in0(andOp_102_in0), .in1(andOp_102_in1), .out(andOp_102_out));

	wire [0:0] notOp_103_in0;
	wire [0:0] notOp_103_out;
	notOp #(.WIDTH(1)) notOp_103(.in(notOp_103_in0), .out(notOp_103_out));

	wire [0:0] andOp_104_in0;
	wire [0:0] andOp_104_in1;
	wire [0:0] andOp_104_out;
	andOp #(.WIDTH(1)) andOp_104(.in0(andOp_104_in0), .in1(andOp_104_in1), .out(andOp_104_out));

	wire [0:0] notOp_105_in0;
	wire [0:0] notOp_105_out;
	notOp #(.WIDTH(1)) notOp_105(.in(notOp_105_in0), .out(notOp_105_out));

	wire [0:0] andOp_106_in0;
	wire [0:0] andOp_106_in1;
	wire [0:0] andOp_106_out;
	andOp #(.WIDTH(1)) andOp_106(.in0(andOp_106_in0), .in1(andOp_106_in1), .out(andOp_106_out));

	wire [0:0] andOp_107_in0;
	wire [0:0] andOp_107_in1;
	wire [0:0] andOp_107_out;
	andOp #(.WIDTH(1)) andOp_107(.in0(andOp_107_in0), .in1(andOp_107_in1), .out(andOp_107_out));

	wire [0:0] notOp_108_in0;
	wire [0:0] notOp_108_out;
	notOp #(.WIDTH(1)) notOp_108(.in(notOp_108_in0), .out(notOp_108_out));

	wire [0:0] andOp_109_in0;
	wire [0:0] andOp_109_in1;
	wire [0:0] andOp_109_out;
	andOp #(.WIDTH(1)) andOp_109(.in0(andOp_109_in0), .in1(andOp_109_in1), .out(andOp_109_out));

	wire [0:0] notOp_110_in0;
	wire [0:0] notOp_110_out;
	notOp #(.WIDTH(1)) notOp_110(.in(notOp_110_in0), .out(notOp_110_out));

	wire [0:0] andOp_111_in0;
	wire [0:0] andOp_111_in1;
	wire [0:0] andOp_111_out;
	andOp #(.WIDTH(1)) andOp_111(.in0(andOp_111_in0), .in1(andOp_111_in1), .out(andOp_111_out));

	wire [0:0] andOp_112_in0;
	wire [0:0] andOp_112_in1;
	wire [0:0] andOp_112_out;
	andOp #(.WIDTH(1)) andOp_112(.in0(andOp_112_in0), .in1(andOp_112_in1), .out(andOp_112_out));

	wire [0:0] notOp_113_in0;
	wire [0:0] notOp_113_out;
	notOp #(.WIDTH(1)) notOp_113(.in(notOp_113_in0), .out(notOp_113_out));

	wire [0:0] andOp_114_in0;
	wire [0:0] andOp_114_in1;
	wire [0:0] andOp_114_out;
	andOp #(.WIDTH(1)) andOp_114(.in0(andOp_114_in0), .in1(andOp_114_in1), .out(andOp_114_out));

	wire [0:0] notOp_115_in0;
	wire [0:0] notOp_115_out;
	notOp #(.WIDTH(1)) notOp_115(.in(notOp_115_in0), .out(notOp_115_out));

	wire [0:0] andOp_116_in0;
	wire [0:0] andOp_116_in1;
	wire [0:0] andOp_116_out;
	andOp #(.WIDTH(1)) andOp_116(.in0(andOp_116_in0), .in1(andOp_116_in1), .out(andOp_116_out));

	wire [0:0] notOp_117_in0;
	wire [0:0] notOp_117_out;
	notOp #(.WIDTH(1)) notOp_117(.in(notOp_117_in0), .out(notOp_117_out));

	wire [0:0] andOp_118_in0;
	wire [0:0] andOp_118_in1;
	wire [0:0] andOp_118_out;
	andOp #(.WIDTH(1)) andOp_118(.in0(andOp_118_in0), .in1(andOp_118_in1), .out(andOp_118_out));

	wire [0:0] notOp_119_in0;
	wire [0:0] notOp_119_out;
	notOp #(.WIDTH(1)) notOp_119(.in(notOp_119_in0), .out(notOp_119_out));

	wire [0:0] andOp_120_in0;
	wire [0:0] andOp_120_in1;
	wire [0:0] andOp_120_out;
	andOp #(.WIDTH(1)) andOp_120(.in0(andOp_120_in0), .in1(andOp_120_in1), .out(andOp_120_out));

	wire [0:0] notOp_121_in0;
	wire [0:0] notOp_121_out;
	notOp #(.WIDTH(1)) notOp_121(.in(notOp_121_in0), .out(notOp_121_out));

	wire [0:0] andOp_122_in0;
	wire [0:0] andOp_122_in1;
	wire [0:0] andOp_122_out;
	andOp #(.WIDTH(1)) andOp_122(.in0(andOp_122_in0), .in1(andOp_122_in1), .out(andOp_122_out));

	wire [0:0] andOp_123_in0;
	wire [0:0] andOp_123_in1;
	wire [0:0] andOp_123_out;
	andOp #(.WIDTH(1)) andOp_123(.in0(andOp_123_in0), .in1(andOp_123_in1), .out(andOp_123_out));

	wire [0:0] notOp_124_in0;
	wire [0:0] notOp_124_out;
	notOp #(.WIDTH(1)) notOp_124(.in(notOp_124_in0), .out(notOp_124_out));

	wire [0:0] andOp_125_in0;
	wire [0:0] andOp_125_in1;
	wire [0:0] andOp_125_out;
	andOp #(.WIDTH(1)) andOp_125(.in0(andOp_125_in0), .in1(andOp_125_in1), .out(andOp_125_out));

	wire [0:0] notOp_126_in0;
	wire [0:0] notOp_126_out;
	notOp #(.WIDTH(1)) notOp_126(.in(notOp_126_in0), .out(notOp_126_out));

	wire [0:0] andOp_127_in0;
	wire [0:0] andOp_127_in1;
	wire [0:0] andOp_127_out;
	andOp #(.WIDTH(1)) andOp_127(.in0(andOp_127_in0), .in1(andOp_127_in1), .out(andOp_127_out));

	wire [0:0] notOp_128_in0;
	wire [0:0] notOp_128_out;
	notOp #(.WIDTH(1)) notOp_128(.in(notOp_128_in0), .out(notOp_128_out));

	wire [0:0] andOp_129_in0;
	wire [0:0] andOp_129_in1;
	wire [0:0] andOp_129_out;
	andOp #(.WIDTH(1)) andOp_129(.in0(andOp_129_in0), .in1(andOp_129_in1), .out(andOp_129_out));

	wire [0:0] notOp_130_in0;
	wire [0:0] notOp_130_out;
	notOp #(.WIDTH(1)) notOp_130(.in(notOp_130_in0), .out(notOp_130_out));

	wire [0:0] andOp_131_in0;
	wire [0:0] andOp_131_in1;
	wire [0:0] andOp_131_out;
	andOp #(.WIDTH(1)) andOp_131(.in0(andOp_131_in0), .in1(andOp_131_in1), .out(andOp_131_out));

	wire [0:0] notOp_132_in0;
	wire [0:0] notOp_132_out;
	notOp #(.WIDTH(1)) notOp_132(.in(notOp_132_in0), .out(notOp_132_out));

	wire [0:0] andOp_133_in0;
	wire [0:0] andOp_133_in1;
	wire [0:0] andOp_133_out;
	andOp #(.WIDTH(1)) andOp_133(.in0(andOp_133_in0), .in1(andOp_133_in1), .out(andOp_133_out));

	wire [0:0] andOp_134_in0;
	wire [0:0] andOp_134_in1;
	wire [0:0] andOp_134_out;
	andOp #(.WIDTH(1)) andOp_134(.in0(andOp_134_in0), .in1(andOp_134_in1), .out(andOp_134_out));

	wire [0:0] notOp_135_in0;
	wire [0:0] notOp_135_out;
	notOp #(.WIDTH(1)) notOp_135(.in(notOp_135_in0), .out(notOp_135_out));

	wire [0:0] andOp_136_in0;
	wire [0:0] andOp_136_in1;
	wire [0:0] andOp_136_out;
	andOp #(.WIDTH(1)) andOp_136(.in0(andOp_136_in0), .in1(andOp_136_in1), .out(andOp_136_out));

	wire [0:0] notOp_137_in0;
	wire [0:0] notOp_137_out;
	notOp #(.WIDTH(1)) notOp_137(.in(notOp_137_in0), .out(notOp_137_out));

	wire [0:0] andOp_138_in0;
	wire [0:0] andOp_138_in1;
	wire [0:0] andOp_138_out;
	andOp #(.WIDTH(1)) andOp_138(.in0(andOp_138_in0), .in1(andOp_138_in1), .out(andOp_138_out));

	wire [0:0] notOp_139_in0;
	wire [0:0] notOp_139_out;
	notOp #(.WIDTH(1)) notOp_139(.in(notOp_139_in0), .out(notOp_139_out));

	wire [0:0] andOp_140_in0;
	wire [0:0] andOp_140_in1;
	wire [0:0] andOp_140_out;
	andOp #(.WIDTH(1)) andOp_140(.in0(andOp_140_in0), .in1(andOp_140_in1), .out(andOp_140_out));

	wire [0:0] andOp_141_in0;
	wire [0:0] andOp_141_in1;
	wire [0:0] andOp_141_out;
	andOp #(.WIDTH(1)) andOp_141(.in0(andOp_141_in0), .in1(andOp_141_in1), .out(andOp_141_out));

	wire [0:0] notOp_142_in0;
	wire [0:0] notOp_142_out;
	notOp #(.WIDTH(1)) notOp_142(.in(notOp_142_in0), .out(notOp_142_out));

	wire [31:0] eq_143_in0;
	wire [31:0] eq_143_in1;
	wire [0:0] eq_143_out;
	eq #(.WIDTH(32)) eq_143(.in0(eq_143_in0), .in1(eq_143_in1), .out(eq_143_out));

	wire [31:0] eq_144_in0;
	wire [31:0] eq_144_in1;
	wire [0:0] eq_144_out;
	eq #(.WIDTH(32)) eq_144(.in0(eq_144_in0), .in1(eq_144_in1), .out(eq_144_out));

	wire [0:0] orOp_145_in0;
	wire [0:0] orOp_145_in1;
	wire [0:0] orOp_145_out;
	orOp #(.WIDTH(1)) orOp_145(.in0(orOp_145_in0), .in1(orOp_145_in1), .out(orOp_145_out));

	wire [31:0] eq_146_in0;
	wire [31:0] eq_146_in1;
	wire [0:0] eq_146_out;
	eq #(.WIDTH(32)) eq_146(.in0(eq_146_in0), .in1(eq_146_in1), .out(eq_146_out));

	wire [0:0] orOp_147_in0;
	wire [0:0] orOp_147_in1;
	wire [0:0] orOp_147_out;
	orOp #(.WIDTH(1)) orOp_147(.in0(orOp_147_in0), .in1(orOp_147_in1), .out(orOp_147_out));

	wire [31:0] eq_148_in0;
	wire [31:0] eq_148_in1;
	wire [0:0] eq_148_out;
	eq #(.WIDTH(32)) eq_148(.in0(eq_148_in0), .in1(eq_148_in1), .out(eq_148_out));

	wire [31:0] eq_149_in0;
	wire [31:0] eq_149_in1;
	wire [0:0] eq_149_out;
	eq #(.WIDTH(32)) eq_149(.in0(eq_149_in0), .in1(eq_149_in1), .out(eq_149_out));

	wire [31:0] eq_150_in0;
	wire [31:0] eq_150_in1;
	wire [0:0] eq_150_out;
	eq #(.WIDTH(32)) eq_150(.in0(eq_150_in0), .in1(eq_150_in1), .out(eq_150_out));

	wire [0:0] orOp_151_in0;
	wire [0:0] orOp_151_in1;
	wire [0:0] orOp_151_out;
	orOp #(.WIDTH(1)) orOp_151(.in0(orOp_151_in0), .in1(orOp_151_in1), .out(orOp_151_out));

	wire [31:0] eq_152_in0;
	wire [31:0] eq_152_in1;
	wire [0:0] eq_152_out;
	eq #(.WIDTH(32)) eq_152(.in0(eq_152_in0), .in1(eq_152_in1), .out(eq_152_out));

	wire [31:0] eq_153_in0;
	wire [31:0] eq_153_in1;
	wire [0:0] eq_153_out;
	eq #(.WIDTH(32)) eq_153(.in0(eq_153_in0), .in1(eq_153_in1), .out(eq_153_out));

	wire [0:0] orOp_154_in0;
	wire [0:0] orOp_154_in1;
	wire [0:0] orOp_154_out;
	orOp #(.WIDTH(1)) orOp_154(.in0(orOp_154_in0), .in1(orOp_154_in1), .out(orOp_154_out));

	wire [31:0] eq_155_in0;
	wire [31:0] eq_155_in1;
	wire [0:0] eq_155_out;
	eq #(.WIDTH(32)) eq_155(.in0(eq_155_in0), .in1(eq_155_in1), .out(eq_155_out));

	wire [0:0] orOp_156_in0;
	wire [0:0] orOp_156_in1;
	wire [0:0] orOp_156_out;
	orOp #(.WIDTH(1)) orOp_156(.in0(orOp_156_in0), .in1(orOp_156_in1), .out(orOp_156_out));

	wire [31:0] eq_157_in0;
	wire [31:0] eq_157_in1;
	wire [0:0] eq_157_out;
	eq #(.WIDTH(32)) eq_157(.in0(eq_157_in0), .in1(eq_157_in1), .out(eq_157_out));

	wire [31:0] eq_158_in0;
	wire [31:0] eq_158_in1;
	wire [0:0] eq_158_out;
	eq #(.WIDTH(32)) eq_158(.in0(eq_158_in0), .in1(eq_158_in1), .out(eq_158_out));

	wire [31:0] eq_159_in0;
	wire [31:0] eq_159_in1;
	wire [0:0] eq_159_out;
	eq #(.WIDTH(32)) eq_159(.in0(eq_159_in0), .in1(eq_159_in1), .out(eq_159_out));

	wire [0:0] orOp_160_in0;
	wire [0:0] orOp_160_in1;
	wire [0:0] orOp_160_out;
	orOp #(.WIDTH(1)) orOp_160(.in0(orOp_160_in0), .in1(orOp_160_in1), .out(orOp_160_out));

	wire [31:0] eq_161_in0;
	wire [31:0] eq_161_in1;
	wire [0:0] eq_161_out;
	eq #(.WIDTH(32)) eq_161(.in0(eq_161_in0), .in1(eq_161_in1), .out(eq_161_out));

	wire [0:0] orOp_162_in0;
	wire [0:0] orOp_162_in1;
	wire [0:0] orOp_162_out;
	orOp #(.WIDTH(1)) orOp_162(.in0(orOp_162_in0), .in1(orOp_162_in1), .out(orOp_162_out));

	wire [31:0] eq_163_in0;
	wire [31:0] eq_163_in1;
	wire [0:0] eq_163_out;
	eq #(.WIDTH(32)) eq_163(.in0(eq_163_in0), .in1(eq_163_in1), .out(eq_163_out));

	wire [31:0] eq_164_in0;
	wire [31:0] eq_164_in1;
	wire [0:0] eq_164_out;
	eq #(.WIDTH(32)) eq_164(.in0(eq_164_in0), .in1(eq_164_in1), .out(eq_164_out));

	wire [0:0] orOp_165_in0;
	wire [0:0] orOp_165_in1;
	wire [0:0] orOp_165_out;
	orOp #(.WIDTH(1)) orOp_165(.in0(orOp_165_in0), .in1(orOp_165_in1), .out(orOp_165_out));

	wire [31:0] eq_166_in0;
	wire [31:0] eq_166_in1;
	wire [0:0] eq_166_out;
	eq #(.WIDTH(32)) eq_166(.in0(eq_166_in0), .in1(eq_166_in1), .out(eq_166_out));

	wire [0:0] orOp_167_in0;
	wire [0:0] orOp_167_in1;
	wire [0:0] orOp_167_out;
	orOp #(.WIDTH(1)) orOp_167(.in0(orOp_167_in0), .in1(orOp_167_in1), .out(orOp_167_out));

	wire [31:0] eq_168_in0;
	wire [31:0] eq_168_in1;
	wire [0:0] eq_168_out;
	eq #(.WIDTH(32)) eq_168(.in0(eq_168_in0), .in1(eq_168_in1), .out(eq_168_out));

	wire [31:0] eq_169_in0;
	wire [31:0] eq_169_in1;
	wire [0:0] eq_169_out;
	eq #(.WIDTH(32)) eq_169(.in0(eq_169_in0), .in1(eq_169_in1), .out(eq_169_out));

	wire [31:0] eq_170_in0;
	wire [31:0] eq_170_in1;
	wire [0:0] eq_170_out;
	eq #(.WIDTH(32)) eq_170(.in0(eq_170_in0), .in1(eq_170_in1), .out(eq_170_out));

	wire [0:0] orOp_171_in0;
	wire [0:0] orOp_171_in1;
	wire [0:0] orOp_171_out;
	orOp #(.WIDTH(1)) orOp_171(.in0(orOp_171_in0), .in1(orOp_171_in1), .out(orOp_171_out));

	wire [31:0] eq_172_in0;
	wire [31:0] eq_172_in1;
	wire [0:0] eq_172_out;
	eq #(.WIDTH(32)) eq_172(.in0(eq_172_in0), .in1(eq_172_in1), .out(eq_172_out));

	wire [0:0] orOp_173_in0;
	wire [0:0] orOp_173_in1;
	wire [0:0] orOp_173_out;
	orOp #(.WIDTH(1)) orOp_173(.in0(orOp_173_in0), .in1(orOp_173_in1), .out(orOp_173_out));

	wire [31:0] eq_174_in0;
	wire [31:0] eq_174_in1;
	wire [0:0] eq_174_out;
	eq #(.WIDTH(32)) eq_174(.in0(eq_174_in0), .in1(eq_174_in1), .out(eq_174_out));

	wire [31:0] eq_175_in0;
	wire [31:0] eq_175_in1;
	wire [0:0] eq_175_out;
	eq #(.WIDTH(32)) eq_175(.in0(eq_175_in0), .in1(eq_175_in1), .out(eq_175_out));

	wire [31:0] eq_176_in0;
	wire [31:0] eq_176_in1;
	wire [0:0] eq_176_out;
	eq #(.WIDTH(32)) eq_176(.in0(eq_176_in0), .in1(eq_176_in1), .out(eq_176_out));

	wire [0:0] orOp_177_in0;
	wire [0:0] orOp_177_in1;
	wire [0:0] orOp_177_out;
	orOp #(.WIDTH(1)) orOp_177(.in0(orOp_177_in0), .in1(orOp_177_in1), .out(orOp_177_out));

	wire [31:0] eq_178_in0;
	wire [31:0] eq_178_in1;
	wire [0:0] eq_178_out;
	eq #(.WIDTH(32)) eq_178(.in0(eq_178_in0), .in1(eq_178_in1), .out(eq_178_out));

	wire [0:0] orOp_179_in0;
	wire [0:0] orOp_179_in1;
	wire [0:0] orOp_179_out;
	orOp #(.WIDTH(1)) orOp_179(.in0(orOp_179_in0), .in1(orOp_179_in1), .out(orOp_179_out));

	wire [31:0] eq_180_in0;
	wire [31:0] eq_180_in1;
	wire [0:0] eq_180_out;
	eq #(.WIDTH(32)) eq_180(.in0(eq_180_in0), .in1(eq_180_in1), .out(eq_180_out));

	wire [31:0] eq_181_in0;
	wire [31:0] eq_181_in1;
	wire [0:0] eq_181_out;
	eq #(.WIDTH(32)) eq_181(.in0(eq_181_in0), .in1(eq_181_in1), .out(eq_181_out));

	wire [0:0] orOp_182_in0;
	wire [0:0] orOp_182_in1;
	wire [0:0] orOp_182_out;
	orOp #(.WIDTH(1)) orOp_182(.in0(orOp_182_in0), .in1(orOp_182_in1), .out(orOp_182_out));

	wire [31:0] eq_183_in0;
	wire [31:0] eq_183_in1;
	wire [0:0] eq_183_out;
	eq #(.WIDTH(32)) eq_183(.in0(eq_183_in0), .in1(eq_183_in1), .out(eq_183_out));

	wire [31:0] eq_184_in0;
	wire [31:0] eq_184_in1;
	wire [0:0] eq_184_out;
	eq #(.WIDTH(32)) eq_184(.in0(eq_184_in0), .in1(eq_184_in1), .out(eq_184_out));

	wire [31:0] eq_185_in0;
	wire [31:0] eq_185_in1;
	wire [0:0] eq_185_out;
	eq #(.WIDTH(32)) eq_185(.in0(eq_185_in0), .in1(eq_185_in1), .out(eq_185_out));

	wire [31:0] eq_186_in0;
	wire [31:0] eq_186_in1;
	wire [0:0] eq_186_out;
	eq #(.WIDTH(32)) eq_186(.in0(eq_186_in0), .in1(eq_186_in1), .out(eq_186_out));

	wire [0:0] notOp_187_in0;
	wire [0:0] notOp_187_out;
	notOp #(.WIDTH(1)) notOp_187(.in(notOp_187_in0), .out(notOp_187_out));

	wire [0:0] andOp_188_in0;
	wire [0:0] andOp_188_in1;
	wire [0:0] andOp_188_out;
	andOp #(.WIDTH(1)) andOp_188(.in0(andOp_188_in0), .in1(andOp_188_in1), .out(andOp_188_out));

	wire [31:0] eq_189_in0;
	wire [31:0] eq_189_in1;
	wire [0:0] eq_189_out;
	eq #(.WIDTH(32)) eq_189(.in0(eq_189_in0), .in1(eq_189_in1), .out(eq_189_out));

	wire [0:0] notOp_190_in0;
	wire [0:0] notOp_190_out;
	notOp #(.WIDTH(1)) notOp_190(.in(notOp_190_in0), .out(notOp_190_out));

	wire [0:0] andOp_191_in0;
	wire [0:0] andOp_191_in1;
	wire [0:0] andOp_191_out;
	andOp #(.WIDTH(1)) andOp_191(.in0(andOp_191_in0), .in1(andOp_191_in1), .out(andOp_191_out));

	wire [31:0] eq_192_in0;
	wire [31:0] eq_192_in1;
	wire [0:0] eq_192_out;
	eq #(.WIDTH(32)) eq_192(.in0(eq_192_in0), .in1(eq_192_in1), .out(eq_192_out));

	wire [31:0] eq_193_in0;
	wire [31:0] eq_193_in1;
	wire [0:0] eq_193_out;
	eq #(.WIDTH(32)) eq_193(.in0(eq_193_in0), .in1(eq_193_in1), .out(eq_193_out));

	wire [31:0] eq_194_in0;
	wire [31:0] eq_194_in1;
	wire [0:0] eq_194_out;
	eq #(.WIDTH(32)) eq_194(.in0(eq_194_in0), .in1(eq_194_in1), .out(eq_194_out));

	wire [0:0] notOp_195_in0;
	wire [0:0] notOp_195_out;
	notOp #(.WIDTH(1)) notOp_195(.in(notOp_195_in0), .out(notOp_195_out));

	wire [0:0] andOp_196_in0;
	wire [0:0] andOp_196_in1;
	wire [0:0] andOp_196_out;
	andOp #(.WIDTH(1)) andOp_196(.in0(andOp_196_in0), .in1(andOp_196_in1), .out(andOp_196_out));

	wire [31:0] eq_197_in0;
	wire [31:0] eq_197_in1;
	wire [0:0] eq_197_out;
	eq #(.WIDTH(32)) eq_197(.in0(eq_197_in0), .in1(eq_197_in1), .out(eq_197_out));

	wire [31:0] eq_198_in0;
	wire [31:0] eq_198_in1;
	wire [0:0] eq_198_out;
	eq #(.WIDTH(32)) eq_198(.in0(eq_198_in0), .in1(eq_198_in1), .out(eq_198_out));

	wire [0:0] notOp_199_in0;
	wire [0:0] notOp_199_out;
	notOp #(.WIDTH(1)) notOp_199(.in(notOp_199_in0), .out(notOp_199_out));

	wire [0:0] andOp_200_in0;
	wire [0:0] andOp_200_in1;
	wire [0:0] andOp_200_out;
	andOp #(.WIDTH(1)) andOp_200(.in0(andOp_200_in0), .in1(andOp_200_in1), .out(andOp_200_out));

	wire [31:0] eq_201_in0;
	wire [31:0] eq_201_in1;
	wire [0:0] eq_201_out;
	eq #(.WIDTH(32)) eq_201(.in0(eq_201_in0), .in1(eq_201_in1), .out(eq_201_out));

	wire [0:0] notOp_202_in0;
	wire [0:0] notOp_202_out;
	notOp #(.WIDTH(1)) notOp_202(.in(notOp_202_in0), .out(notOp_202_out));

	wire [0:0] andOp_203_in0;
	wire [0:0] andOp_203_in1;
	wire [0:0] andOp_203_out;
	andOp #(.WIDTH(1)) andOp_203(.in0(andOp_203_in0), .in1(andOp_203_in1), .out(andOp_203_out));

	wire [31:0] eq_204_in0;
	wire [31:0] eq_204_in1;
	wire [0:0] eq_204_out;
	eq #(.WIDTH(32)) eq_204(.in0(eq_204_in0), .in1(eq_204_in1), .out(eq_204_out));

	wire [31:0] eq_205_in0;
	wire [31:0] eq_205_in1;
	wire [0:0] eq_205_out;
	eq #(.WIDTH(32)) eq_205(.in0(eq_205_in0), .in1(eq_205_in1), .out(eq_205_out));

	wire [31:0] eq_206_in0;
	wire [31:0] eq_206_in1;
	wire [0:0] eq_206_out;
	eq #(.WIDTH(32)) eq_206(.in0(eq_206_in0), .in1(eq_206_in1), .out(eq_206_out));

	wire [0:0] notOp_207_in0;
	wire [0:0] notOp_207_out;
	notOp #(.WIDTH(1)) notOp_207(.in(notOp_207_in0), .out(notOp_207_out));

	wire [0:0] andOp_208_in0;
	wire [0:0] andOp_208_in1;
	wire [0:0] andOp_208_out;
	andOp #(.WIDTH(1)) andOp_208(.in0(andOp_208_in0), .in1(andOp_208_in1), .out(andOp_208_out));

	wire [31:0] eq_209_in0;
	wire [31:0] eq_209_in1;
	wire [0:0] eq_209_out;
	eq #(.WIDTH(32)) eq_209(.in0(eq_209_in0), .in1(eq_209_in1), .out(eq_209_out));

	wire [0:0] notOp_210_in0;
	wire [0:0] notOp_210_out;
	notOp #(.WIDTH(1)) notOp_210(.in(notOp_210_in0), .out(notOp_210_out));

	wire [0:0] andOp_211_in0;
	wire [0:0] andOp_211_in1;
	wire [0:0] andOp_211_out;
	andOp #(.WIDTH(1)) andOp_211(.in0(andOp_211_in0), .in1(andOp_211_in1), .out(andOp_211_out));

	wire [31:0] eq_212_in0;
	wire [31:0] eq_212_in1;
	wire [0:0] eq_212_out;
	eq #(.WIDTH(32)) eq_212(.in0(eq_212_in0), .in1(eq_212_in1), .out(eq_212_out));

	wire [31:0] eq_213_in0;
	wire [31:0] eq_213_in1;
	wire [0:0] eq_213_out;
	eq #(.WIDTH(32)) eq_213(.in0(eq_213_in0), .in1(eq_213_in1), .out(eq_213_out));

	wire [0:0] notOp_214_in0;
	wire [0:0] notOp_214_out;
	notOp #(.WIDTH(1)) notOp_214(.in(notOp_214_in0), .out(notOp_214_out));

	wire [0:0] andOp_215_in0;
	wire [0:0] andOp_215_in1;
	wire [0:0] andOp_215_out;
	andOp #(.WIDTH(1)) andOp_215(.in0(andOp_215_in0), .in1(andOp_215_in1), .out(andOp_215_out));

	wire [31:0] eq_216_in0;
	wire [31:0] eq_216_in1;
	wire [0:0] eq_216_out;
	eq #(.WIDTH(32)) eq_216(.in0(eq_216_in0), .in1(eq_216_in1), .out(eq_216_out));

	wire [0:0] notOp_217_in0;
	wire [0:0] notOp_217_out;
	notOp #(.WIDTH(1)) notOp_217(.in(notOp_217_in0), .out(notOp_217_out));

	wire [0:0] andOp_218_in0;
	wire [0:0] andOp_218_in1;
	wire [0:0] andOp_218_out;
	andOp #(.WIDTH(1)) andOp_218(.in0(andOp_218_in0), .in1(andOp_218_in1), .out(andOp_218_out));

	wire [31:0] eq_219_in0;
	wire [31:0] eq_219_in1;
	wire [0:0] eq_219_out;
	eq #(.WIDTH(32)) eq_219(.in0(eq_219_in0), .in1(eq_219_in1), .out(eq_219_out));

	wire [31:0] eq_220_in0;
	wire [31:0] eq_220_in1;
	wire [0:0] eq_220_out;
	eq #(.WIDTH(32)) eq_220(.in0(eq_220_in0), .in1(eq_220_in1), .out(eq_220_out));

	wire [31:0] eq_221_in0;
	wire [31:0] eq_221_in1;
	wire [0:0] eq_221_out;
	eq #(.WIDTH(32)) eq_221(.in0(eq_221_in0), .in1(eq_221_in1), .out(eq_221_out));

	wire [0:0] notOp_222_in0;
	wire [0:0] notOp_222_out;
	notOp #(.WIDTH(1)) notOp_222(.in(notOp_222_in0), .out(notOp_222_out));

	wire [0:0] andOp_223_in0;
	wire [0:0] andOp_223_in1;
	wire [0:0] andOp_223_out;
	andOp #(.WIDTH(1)) andOp_223(.in0(andOp_223_in0), .in1(andOp_223_in1), .out(andOp_223_out));

	wire [31:0] eq_224_in0;
	wire [31:0] eq_224_in1;
	wire [0:0] eq_224_out;
	eq #(.WIDTH(32)) eq_224(.in0(eq_224_in0), .in1(eq_224_in1), .out(eq_224_out));

	wire [0:0] notOp_225_in0;
	wire [0:0] notOp_225_out;
	notOp #(.WIDTH(1)) notOp_225(.in(notOp_225_in0), .out(notOp_225_out));

	wire [0:0] andOp_226_in0;
	wire [0:0] andOp_226_in1;
	wire [0:0] andOp_226_out;
	andOp #(.WIDTH(1)) andOp_226(.in0(andOp_226_in0), .in1(andOp_226_in1), .out(andOp_226_out));

	wire [31:0] eq_227_in0;
	wire [31:0] eq_227_in1;
	wire [0:0] eq_227_out;
	eq #(.WIDTH(32)) eq_227(.in0(eq_227_in0), .in1(eq_227_in1), .out(eq_227_out));

	wire [31:0] eq_228_in0;
	wire [31:0] eq_228_in1;
	wire [0:0] eq_228_out;
	eq #(.WIDTH(32)) eq_228(.in0(eq_228_in0), .in1(eq_228_in1), .out(eq_228_out));

	wire [31:0] eq_229_in0;
	wire [31:0] eq_229_in1;
	wire [0:0] eq_229_out;
	eq #(.WIDTH(32)) eq_229(.in0(eq_229_in0), .in1(eq_229_in1), .out(eq_229_out));

	wire [0:0] notOp_230_in0;
	wire [0:0] notOp_230_out;
	notOp #(.WIDTH(1)) notOp_230(.in(notOp_230_in0), .out(notOp_230_out));

	wire [0:0] andOp_231_in0;
	wire [0:0] andOp_231_in1;
	wire [0:0] andOp_231_out;
	andOp #(.WIDTH(1)) andOp_231(.in0(andOp_231_in0), .in1(andOp_231_in1), .out(andOp_231_out));

	wire [31:0] eq_232_in0;
	wire [31:0] eq_232_in1;
	wire [0:0] eq_232_out;
	eq #(.WIDTH(32)) eq_232(.in0(eq_232_in0), .in1(eq_232_in1), .out(eq_232_out));

	wire [0:0] notOp_233_in0;
	wire [0:0] notOp_233_out;
	notOp #(.WIDTH(1)) notOp_233(.in(notOp_233_in0), .out(notOp_233_out));

	wire [0:0] andOp_234_in0;
	wire [0:0] andOp_234_in1;
	wire [0:0] andOp_234_out;
	andOp #(.WIDTH(1)) andOp_234(.in0(andOp_234_in0), .in1(andOp_234_in1), .out(andOp_234_out));

	wire [31:0] eq_235_in0;
	wire [31:0] eq_235_in1;
	wire [0:0] eq_235_out;
	eq #(.WIDTH(32)) eq_235(.in0(eq_235_in0), .in1(eq_235_in1), .out(eq_235_out));

	wire [31:0] eq_236_in0;
	wire [31:0] eq_236_in1;
	wire [0:0] eq_236_out;
	eq #(.WIDTH(32)) eq_236(.in0(eq_236_in0), .in1(eq_236_in1), .out(eq_236_out));

	wire [0:0] notOp_237_in0;
	wire [0:0] notOp_237_out;
	notOp #(.WIDTH(1)) notOp_237(.in(notOp_237_in0), .out(notOp_237_out));

	wire [0:0] andOp_238_in0;
	wire [0:0] andOp_238_in1;
	wire [0:0] andOp_238_out;
	andOp #(.WIDTH(1)) andOp_238(.in0(andOp_238_in0), .in1(andOp_238_in1), .out(andOp_238_out));

	wire [31:0] eq_239_in0;
	wire [31:0] eq_239_in1;
	wire [0:0] eq_239_out;
	eq #(.WIDTH(32)) eq_239(.in0(eq_239_in0), .in1(eq_239_in1), .out(eq_239_out));

	wire [31:0] eq_240_in0;
	wire [31:0] eq_240_in1;
	wire [0:0] eq_240_out;
	eq #(.WIDTH(32)) eq_240(.in0(eq_240_in0), .in1(eq_240_in1), .out(eq_240_out));

	wire [0:0] andOp_241_in0;
	wire [0:0] andOp_241_in1;
	wire [0:0] andOp_241_out;
	andOp #(.WIDTH(1)) andOp_241(.in0(andOp_241_in0), .in1(andOp_241_in1), .out(andOp_241_out));

	wire [0:0] andOp_242_in0;
	wire [0:0] andOp_242_in1;
	wire [0:0] andOp_242_out;
	andOp #(.WIDTH(1)) andOp_242(.in0(andOp_242_in0), .in1(andOp_242_in1), .out(andOp_242_out));

	wire [0:0] andOp_243_in0;
	wire [0:0] andOp_243_in1;
	wire [0:0] andOp_243_out;
	andOp #(.WIDTH(1)) andOp_243(.in0(andOp_243_in0), .in1(andOp_243_in1), .out(andOp_243_out));

	wire [0:0] andOp_244_in0;
	wire [0:0] andOp_244_in1;
	wire [0:0] andOp_244_out;
	andOp #(.WIDTH(1)) andOp_244(.in0(andOp_244_in0), .in1(andOp_244_in1), .out(andOp_244_out));

	wire [0:0] andOp_245_in0;
	wire [0:0] andOp_245_in1;
	wire [0:0] andOp_245_out;
	andOp #(.WIDTH(1)) andOp_245(.in0(andOp_245_in0), .in1(andOp_245_in1), .out(andOp_245_out));

	wire [0:0] andOp_246_in0;
	wire [0:0] andOp_246_in1;
	wire [0:0] andOp_246_out;
	andOp #(.WIDTH(1)) andOp_246(.in0(andOp_246_in0), .in1(andOp_246_in1), .out(andOp_246_out));

	wire [0:0] andOp_247_in0;
	wire [0:0] andOp_247_in1;
	wire [0:0] andOp_247_out;
	andOp #(.WIDTH(1)) andOp_247(.in0(andOp_247_in0), .in1(andOp_247_in1), .out(andOp_247_out));

	wire [0:0] andOp_248_in0;
	wire [0:0] andOp_248_in1;
	wire [0:0] andOp_248_out;
	andOp #(.WIDTH(1)) andOp_248(.in0(andOp_248_in0), .in1(andOp_248_in1), .out(andOp_248_out));

	wire [0:0] andOp_249_in0;
	wire [0:0] andOp_249_in1;
	wire [0:0] andOp_249_out;
	andOp #(.WIDTH(1)) andOp_249(.in0(andOp_249_in0), .in1(andOp_249_in1), .out(andOp_249_out));

	wire [0:0] andOp_250_in0;
	wire [0:0] andOp_250_in1;
	wire [0:0] andOp_250_out;
	andOp #(.WIDTH(1)) andOp_250(.in0(andOp_250_in0), .in1(andOp_250_in1), .out(andOp_250_out));

	wire [0:0] andOp_251_in0;
	wire [0:0] andOp_251_in1;
	wire [0:0] andOp_251_out;
	andOp #(.WIDTH(1)) andOp_251(.in0(andOp_251_in0), .in1(andOp_251_in1), .out(andOp_251_out));

	wire [31:0] concat_252_in0;
	wire [31:0] concat_252_in1;
	wire [63:0] concat_252_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_252(.in0(concat_252_in0), .in1(concat_252_in1), .out(concat_252_out));

	wire [31:0] concat_253_in0;
	wire [31:0] concat_253_in1;
	wire [63:0] concat_253_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_253(.in0(concat_253_in0), .in1(concat_253_in1), .out(concat_253_out));

	wire [0:0] andOp_254_in0;
	wire [0:0] andOp_254_in1;
	wire [0:0] andOp_254_out;
	andOp #(.WIDTH(1)) andOp_254(.in0(andOp_254_in0), .in1(andOp_254_in1), .out(andOp_254_out));

	wire [0:0] andOp_255_in0;
	wire [0:0] andOp_255_in1;
	wire [0:0] andOp_255_out;
	andOp #(.WIDTH(1)) andOp_255(.in0(andOp_255_in0), .in1(andOp_255_in1), .out(andOp_255_out));

	wire [0:0] andOp_256_in0;
	wire [0:0] andOp_256_in1;
	wire [0:0] andOp_256_out;
	andOp #(.WIDTH(1)) andOp_256(.in0(andOp_256_in0), .in1(andOp_256_in1), .out(andOp_256_out));

	wire [0:0] andOp_257_in0;
	wire [0:0] andOp_257_in1;
	wire [0:0] andOp_257_out;
	andOp #(.WIDTH(1)) andOp_257(.in0(andOp_257_in0), .in1(andOp_257_in1), .out(andOp_257_out));

	wire [0:0] andOp_258_in0;
	wire [0:0] andOp_258_in1;
	wire [0:0] andOp_258_out;
	andOp #(.WIDTH(1)) andOp_258(.in0(andOp_258_in0), .in1(andOp_258_in1), .out(andOp_258_out));

	wire [0:0] andOp_259_in0;
	wire [0:0] andOp_259_in1;
	wire [0:0] andOp_259_out;
	andOp #(.WIDTH(1)) andOp_259(.in0(andOp_259_in0), .in1(andOp_259_in1), .out(andOp_259_out));

	wire [0:0] andOp_260_in0;
	wire [0:0] andOp_260_in1;
	wire [0:0] andOp_260_out;
	andOp #(.WIDTH(1)) andOp_260(.in0(andOp_260_in0), .in1(andOp_260_in1), .out(andOp_260_out));

	wire [31:0] concat_261_in0;
	wire [31:0] concat_261_in1;
	wire [63:0] concat_261_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_261(.in0(concat_261_in0), .in1(concat_261_in1), .out(concat_261_out));

	wire [31:0] concat_262_in0;
	wire [31:0] concat_262_in1;
	wire [63:0] concat_262_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_262(.in0(concat_262_in0), .in1(concat_262_in1), .out(concat_262_out));

	wire [0:0] andOp_263_in0;
	wire [0:0] andOp_263_in1;
	wire [0:0] andOp_263_out;
	andOp #(.WIDTH(1)) andOp_263(.in0(andOp_263_in0), .in1(andOp_263_in1), .out(andOp_263_out));

	wire [0:0] andOp_264_in0;
	wire [0:0] andOp_264_in1;
	wire [0:0] andOp_264_out;
	andOp #(.WIDTH(1)) andOp_264(.in0(andOp_264_in0), .in1(andOp_264_in1), .out(andOp_264_out));

	wire [0:0] andOp_265_in0;
	wire [0:0] andOp_265_in1;
	wire [0:0] andOp_265_out;
	andOp #(.WIDTH(1)) andOp_265(.in0(andOp_265_in0), .in1(andOp_265_in1), .out(andOp_265_out));

	wire [0:0] andOp_266_in0;
	wire [0:0] andOp_266_in1;
	wire [0:0] andOp_266_out;
	andOp #(.WIDTH(1)) andOp_266(.in0(andOp_266_in0), .in1(andOp_266_in1), .out(andOp_266_out));

	wire [0:0] andOp_267_in0;
	wire [0:0] andOp_267_in1;
	wire [0:0] andOp_267_out;
	andOp #(.WIDTH(1)) andOp_267(.in0(andOp_267_in0), .in1(andOp_267_in1), .out(andOp_267_out));

	wire [0:0] andOp_268_in0;
	wire [0:0] andOp_268_in1;
	wire [0:0] andOp_268_out;
	andOp #(.WIDTH(1)) andOp_268(.in0(andOp_268_in0), .in1(andOp_268_in1), .out(andOp_268_out));

	wire [0:0] andOp_269_in0;
	wire [0:0] andOp_269_in1;
	wire [0:0] andOp_269_out;
	andOp #(.WIDTH(1)) andOp_269(.in0(andOp_269_in0), .in1(andOp_269_in1), .out(andOp_269_out));

	wire [0:0] andOp_270_in0;
	wire [0:0] andOp_270_in1;
	wire [0:0] andOp_270_out;
	andOp #(.WIDTH(1)) andOp_270(.in0(andOp_270_in0), .in1(andOp_270_in1), .out(andOp_270_out));

	wire [0:0] andOp_271_in0;
	wire [0:0] andOp_271_in1;
	wire [0:0] andOp_271_out;
	andOp #(.WIDTH(1)) andOp_271(.in0(andOp_271_in0), .in1(andOp_271_in1), .out(andOp_271_out));

	wire [0:0] andOp_272_in0;
	wire [0:0] andOp_272_in1;
	wire [0:0] andOp_272_out;
	andOp #(.WIDTH(1)) andOp_272(.in0(andOp_272_in0), .in1(andOp_272_in1), .out(andOp_272_out));

	wire [0:0] andOp_273_in0;
	wire [0:0] andOp_273_in1;
	wire [0:0] andOp_273_out;
	andOp #(.WIDTH(1)) andOp_273(.in0(andOp_273_in0), .in1(andOp_273_in1), .out(andOp_273_out));

	wire [0:0] andOp_274_in0;
	wire [0:0] andOp_274_in1;
	wire [0:0] andOp_274_out;
	andOp #(.WIDTH(1)) andOp_274(.in0(andOp_274_in0), .in1(andOp_274_in1), .out(andOp_274_out));

	wire [0:0] andOp_275_in0;
	wire [0:0] andOp_275_in1;
	wire [0:0] andOp_275_out;
	andOp #(.WIDTH(1)) andOp_275(.in0(andOp_275_in0), .in1(andOp_275_in1), .out(andOp_275_out));

	wire [0:0] andOp_276_in0;
	wire [0:0] andOp_276_in1;
	wire [0:0] andOp_276_out;
	andOp #(.WIDTH(1)) andOp_276(.in0(andOp_276_in0), .in1(andOp_276_in1), .out(andOp_276_out));

	wire [0:0] andOp_277_in0;
	wire [0:0] andOp_277_in1;
	wire [0:0] andOp_277_out;
	andOp #(.WIDTH(1)) andOp_277(.in0(andOp_277_in0), .in1(andOp_277_in1), .out(andOp_277_out));

	wire [0:0] notOp_278_in0;
	wire [0:0] notOp_278_out;
	notOp #(.WIDTH(1)) notOp_278(.in(notOp_278_in0), .out(notOp_278_out));

	wire [0:0] andOp_279_in0;
	wire [0:0] andOp_279_in1;
	wire [0:0] andOp_279_out;
	andOp #(.WIDTH(1)) andOp_279(.in0(andOp_279_in0), .in1(andOp_279_in1), .out(andOp_279_out));

	wire [0:0] notOp_280_in0;
	wire [0:0] notOp_280_out;
	notOp #(.WIDTH(1)) notOp_280(.in(notOp_280_in0), .out(notOp_280_out));

	wire [0:0] andOp_281_in0;
	wire [0:0] andOp_281_in1;
	wire [0:0] andOp_281_out;
	andOp #(.WIDTH(1)) andOp_281(.in0(andOp_281_in0), .in1(andOp_281_in1), .out(andOp_281_out));

	wire [0:0] notOp_282_in0;
	wire [0:0] notOp_282_out;
	notOp #(.WIDTH(1)) notOp_282(.in(notOp_282_in0), .out(notOp_282_out));

	wire [0:0] andOp_283_in0;
	wire [0:0] andOp_283_in1;
	wire [0:0] andOp_283_out;
	andOp #(.WIDTH(1)) andOp_283(.in0(andOp_283_in0), .in1(andOp_283_in1), .out(andOp_283_out));

	wire [0:0] notOp_284_in0;
	wire [0:0] notOp_284_out;
	notOp #(.WIDTH(1)) notOp_284(.in(notOp_284_in0), .out(notOp_284_out));

	wire [0:0] andOp_285_in0;
	wire [0:0] andOp_285_in1;
	wire [0:0] andOp_285_out;
	andOp #(.WIDTH(1)) andOp_285(.in0(andOp_285_in0), .in1(andOp_285_in1), .out(andOp_285_out));

	wire [0:0] notOp_286_in0;
	wire [0:0] notOp_286_out;
	notOp #(.WIDTH(1)) notOp_286(.in(notOp_286_in0), .out(notOp_286_out));

	wire [0:0] andOp_287_in0;
	wire [0:0] andOp_287_in1;
	wire [0:0] andOp_287_out;
	andOp #(.WIDTH(1)) andOp_287(.in0(andOp_287_in0), .in1(andOp_287_in1), .out(andOp_287_out));

	wire [0:0] notOp_288_in0;
	wire [0:0] notOp_288_out;
	notOp #(.WIDTH(1)) notOp_288(.in(notOp_288_in0), .out(notOp_288_out));

	wire [0:0] andOp_289_in0;
	wire [0:0] andOp_289_in1;
	wire [0:0] andOp_289_out;
	andOp #(.WIDTH(1)) andOp_289(.in0(andOp_289_in0), .in1(andOp_289_in1), .out(andOp_289_out));

	wire [0:0] notOp_290_in0;
	wire [0:0] notOp_290_out;
	notOp #(.WIDTH(1)) notOp_290(.in(notOp_290_in0), .out(notOp_290_out));

	wire [0:0] andOp_291_in0;
	wire [0:0] andOp_291_in1;
	wire [0:0] andOp_291_out;
	andOp #(.WIDTH(1)) andOp_291(.in0(andOp_291_in0), .in1(andOp_291_in1), .out(andOp_291_out));

	wire [0:0] notOp_292_in0;
	wire [0:0] notOp_292_out;
	notOp #(.WIDTH(1)) notOp_292(.in(notOp_292_in0), .out(notOp_292_out));

	wire [0:0] andOp_293_in0;
	wire [0:0] andOp_293_in1;
	wire [0:0] andOp_293_out;
	andOp #(.WIDTH(1)) andOp_293(.in0(andOp_293_in0), .in1(andOp_293_in1), .out(andOp_293_out));

	wire [0:0] notOp_294_in0;
	wire [0:0] notOp_294_out;
	notOp #(.WIDTH(1)) notOp_294(.in(notOp_294_in0), .out(notOp_294_out));

	wire [0:0] andOp_295_in0;
	wire [0:0] andOp_295_in1;
	wire [0:0] andOp_295_out;
	andOp #(.WIDTH(1)) andOp_295(.in0(andOp_295_in0), .in1(andOp_295_in1), .out(andOp_295_out));

	wire [0:0] notOp_296_in0;
	wire [0:0] notOp_296_out;
	notOp #(.WIDTH(1)) notOp_296(.in(notOp_296_in0), .out(notOp_296_out));

	wire [0:0] andOp_297_in0;
	wire [0:0] andOp_297_in1;
	wire [0:0] andOp_297_out;
	andOp #(.WIDTH(1)) andOp_297(.in0(andOp_297_in0), .in1(andOp_297_in1), .out(andOp_297_out));

	wire [0:0] notOp_298_in0;
	wire [0:0] notOp_298_out;
	notOp #(.WIDTH(1)) notOp_298(.in(notOp_298_in0), .out(notOp_298_out));

	wire [0:0] andOp_299_in0;
	wire [0:0] andOp_299_in1;
	wire [0:0] andOp_299_out;
	andOp #(.WIDTH(1)) andOp_299(.in0(andOp_299_in0), .in1(andOp_299_in1), .out(andOp_299_out));

	wire [0:0] notOp_300_in0;
	wire [0:0] notOp_300_out;
	notOp #(.WIDTH(1)) notOp_300(.in(notOp_300_in0), .out(notOp_300_out));

	wire [0:0] andOp_301_in0;
	wire [0:0] andOp_301_in1;
	wire [0:0] andOp_301_out;
	andOp #(.WIDTH(1)) andOp_301(.in0(andOp_301_in0), .in1(andOp_301_in1), .out(andOp_301_out));

	wire [0:0] notOp_302_in0;
	wire [0:0] notOp_302_out;
	notOp #(.WIDTH(1)) notOp_302(.in(notOp_302_in0), .out(notOp_302_out));

	wire [0:0] andOp_303_in0;
	wire [0:0] andOp_303_in1;
	wire [0:0] andOp_303_out;
	andOp #(.WIDTH(1)) andOp_303(.in0(andOp_303_in0), .in1(andOp_303_in1), .out(andOp_303_out));

	wire [0:0] notOp_304_in0;
	wire [0:0] notOp_304_out;
	notOp #(.WIDTH(1)) notOp_304(.in(notOp_304_in0), .out(notOp_304_out));

	wire [0:0] andOp_305_in0;
	wire [0:0] andOp_305_in1;
	wire [0:0] andOp_305_out;
	andOp #(.WIDTH(1)) andOp_305(.in0(andOp_305_in0), .in1(andOp_305_in1), .out(andOp_305_out));

	wire [0:0] notOp_306_in0;
	wire [0:0] notOp_306_out;
	notOp #(.WIDTH(1)) notOp_306(.in(notOp_306_in0), .out(notOp_306_out));

	wire [0:0] andOp_307_in0;
	wire [0:0] andOp_307_in1;
	wire [0:0] andOp_307_out;
	andOp #(.WIDTH(1)) andOp_307(.in0(andOp_307_in0), .in1(andOp_307_in1), .out(andOp_307_out));

	wire [0:0] notOp_308_in0;
	wire [0:0] notOp_308_out;
	notOp #(.WIDTH(1)) notOp_308(.in(notOp_308_in0), .out(notOp_308_out));

	wire [0:0] andOp_309_in0;
	wire [0:0] andOp_309_in1;
	wire [0:0] andOp_309_out;
	andOp #(.WIDTH(1)) andOp_309(.in0(andOp_309_in0), .in1(andOp_309_in1), .out(andOp_309_out));

	wire [0:0] notOp_310_in0;
	wire [0:0] notOp_310_out;
	notOp #(.WIDTH(1)) notOp_310(.in(notOp_310_in0), .out(notOp_310_out));

	wire [0:0] andOp_311_in0;
	wire [0:0] andOp_311_in1;
	wire [0:0] andOp_311_out;
	andOp #(.WIDTH(1)) andOp_311(.in0(andOp_311_in0), .in1(andOp_311_in1), .out(andOp_311_out));

	wire [0:0] notOp_312_in0;
	wire [0:0] notOp_312_out;
	notOp #(.WIDTH(1)) notOp_312(.in(notOp_312_in0), .out(notOp_312_out));

	wire [0:0] andOp_313_in0;
	wire [0:0] andOp_313_in1;
	wire [0:0] andOp_313_out;
	andOp #(.WIDTH(1)) andOp_313(.in0(andOp_313_in0), .in1(andOp_313_in1), .out(andOp_313_out));

	wire [0:0] notOp_314_in0;
	wire [0:0] notOp_314_out;
	notOp #(.WIDTH(1)) notOp_314(.in(notOp_314_in0), .out(notOp_314_out));

	wire [0:0] andOp_315_in0;
	wire [0:0] andOp_315_in1;
	wire [0:0] andOp_315_out;
	andOp #(.WIDTH(1)) andOp_315(.in0(andOp_315_in0), .in1(andOp_315_in1), .out(andOp_315_out));

	wire [0:0] notOp_316_in0;
	wire [0:0] notOp_316_out;
	notOp #(.WIDTH(1)) notOp_316(.in(notOp_316_in0), .out(notOp_316_out));

	wire [0:0] andOp_317_in0;
	wire [0:0] andOp_317_in1;
	wire [0:0] andOp_317_out;
	andOp #(.WIDTH(1)) andOp_317(.in0(andOp_317_in0), .in1(andOp_317_in1), .out(andOp_317_out));

	wire [0:0] notOp_318_in0;
	wire [0:0] notOp_318_out;
	notOp #(.WIDTH(1)) notOp_318(.in(notOp_318_in0), .out(notOp_318_out));

	wire [0:0] andOp_319_in0;
	wire [0:0] andOp_319_in1;
	wire [0:0] andOp_319_out;
	andOp #(.WIDTH(1)) andOp_319(.in0(andOp_319_in0), .in1(andOp_319_in1), .out(andOp_319_out));

	wire [31:0] eq_320_in0;
	wire [31:0] eq_320_in1;
	wire [0:0] eq_320_out;
	eq #(.WIDTH(32)) eq_320(.in0(eq_320_in0), .in1(eq_320_in1), .out(eq_320_out));

	wire [31:0] eq_321_in0;
	wire [31:0] eq_321_in1;
	wire [0:0] eq_321_out;
	eq #(.WIDTH(32)) eq_321(.in0(eq_321_in0), .in1(eq_321_in1), .out(eq_321_out));

	wire [31:0] eq_322_in0;
	wire [31:0] eq_322_in1;
	wire [0:0] eq_322_out;
	eq #(.WIDTH(32)) eq_322(.in0(eq_322_in0), .in1(eq_322_in1), .out(eq_322_out));

	wire [31:0] eq_323_in0;
	wire [31:0] eq_323_in1;
	wire [0:0] eq_323_out;
	eq #(.WIDTH(32)) eq_323(.in0(eq_323_in0), .in1(eq_323_in1), .out(eq_323_out));

	wire [0:0] andOp_324_in0;
	wire [0:0] andOp_324_in1;
	wire [0:0] andOp_324_out;
	andOp #(.WIDTH(1)) andOp_324(.in0(andOp_324_in0), .in1(andOp_324_in1), .out(andOp_324_out));

	wire [31:0] eq_325_in0;
	wire [31:0] eq_325_in1;
	wire [0:0] eq_325_out;
	eq #(.WIDTH(32)) eq_325(.in0(eq_325_in0), .in1(eq_325_in1), .out(eq_325_out));

	wire [31:0] eq_326_in0;
	wire [31:0] eq_326_in1;
	wire [0:0] eq_326_out;
	eq #(.WIDTH(32)) eq_326(.in0(eq_326_in0), .in1(eq_326_in1), .out(eq_326_out));

	wire [31:0] eq_327_in0;
	wire [31:0] eq_327_in1;
	wire [0:0] eq_327_out;
	eq #(.WIDTH(32)) eq_327(.in0(eq_327_in0), .in1(eq_327_in1), .out(eq_327_out));

	wire [31:0] eq_328_in0;
	wire [31:0] eq_328_in1;
	wire [0:0] eq_328_out;
	eq #(.WIDTH(32)) eq_328(.in0(eq_328_in0), .in1(eq_328_in1), .out(eq_328_out));

	wire [0:0] andOp_329_in0;
	wire [0:0] andOp_329_in1;
	wire [0:0] andOp_329_out;
	andOp #(.WIDTH(1)) andOp_329(.in0(andOp_329_in0), .in1(andOp_329_in1), .out(andOp_329_out));

	wire [31:0] eq_330_in0;
	wire [31:0] eq_330_in1;
	wire [0:0] eq_330_out;
	eq #(.WIDTH(32)) eq_330(.in0(eq_330_in0), .in1(eq_330_in1), .out(eq_330_out));

	wire [31:0] eq_331_in0;
	wire [31:0] eq_331_in1;
	wire [0:0] eq_331_out;
	eq #(.WIDTH(32)) eq_331(.in0(eq_331_in0), .in1(eq_331_in1), .out(eq_331_out));

	wire [31:0] eq_332_in0;
	wire [31:0] eq_332_in1;
	wire [0:0] eq_332_out;
	eq #(.WIDTH(32)) eq_332(.in0(eq_332_in0), .in1(eq_332_in1), .out(eq_332_out));

	wire [31:0] eq_333_in0;
	wire [31:0] eq_333_in1;
	wire [0:0] eq_333_out;
	eq #(.WIDTH(32)) eq_333(.in0(eq_333_in0), .in1(eq_333_in1), .out(eq_333_out));

	wire [0:0] andOp_334_in0;
	wire [0:0] andOp_334_in1;
	wire [0:0] andOp_334_out;
	andOp #(.WIDTH(1)) andOp_334(.in0(andOp_334_in0), .in1(andOp_334_in1), .out(andOp_334_out));

	wire [31:0] eq_335_in0;
	wire [31:0] eq_335_in1;
	wire [0:0] eq_335_out;
	eq #(.WIDTH(32)) eq_335(.in0(eq_335_in0), .in1(eq_335_in1), .out(eq_335_out));

	wire [31:0] eq_336_in0;
	wire [31:0] eq_336_in1;
	wire [0:0] eq_336_out;
	eq #(.WIDTH(32)) eq_336(.in0(eq_336_in0), .in1(eq_336_in1), .out(eq_336_out));

	wire [0:0] andOp_337_in0;
	wire [0:0] andOp_337_in1;
	wire [0:0] andOp_337_out;
	andOp #(.WIDTH(1)) andOp_337(.in0(andOp_337_in0), .in1(andOp_337_in1), .out(andOp_337_out));

	wire [31:0] eq_338_in0;
	wire [31:0] eq_338_in1;
	wire [0:0] eq_338_out;
	eq #(.WIDTH(32)) eq_338(.in0(eq_338_in0), .in1(eq_338_in1), .out(eq_338_out));

	wire [31:0] eq_339_in0;
	wire [31:0] eq_339_in1;
	wire [0:0] eq_339_out;
	eq #(.WIDTH(32)) eq_339(.in0(eq_339_in0), .in1(eq_339_in1), .out(eq_339_out));

	wire [31:0] eq_340_in0;
	wire [31:0] eq_340_in1;
	wire [0:0] eq_340_out;
	eq #(.WIDTH(32)) eq_340(.in0(eq_340_in0), .in1(eq_340_in1), .out(eq_340_out));

	wire [31:0] eq_341_in0;
	wire [31:0] eq_341_in1;
	wire [0:0] eq_341_out;
	eq #(.WIDTH(32)) eq_341(.in0(eq_341_in0), .in1(eq_341_in1), .out(eq_341_out));

	wire [31:0] eq_342_in0;
	wire [31:0] eq_342_in1;
	wire [0:0] eq_342_out;
	eq #(.WIDTH(32)) eq_342(.in0(eq_342_in0), .in1(eq_342_in1), .out(eq_342_out));

	wire [0:0] andOp_343_in0;
	wire [0:0] andOp_343_in1;
	wire [0:0] andOp_343_out;
	andOp #(.WIDTH(1)) andOp_343(.in0(andOp_343_in0), .in1(andOp_343_in1), .out(andOp_343_out));

	wire [31:0] eq_344_in0;
	wire [31:0] eq_344_in1;
	wire [0:0] eq_344_out;
	eq #(.WIDTH(32)) eq_344(.in0(eq_344_in0), .in1(eq_344_in1), .out(eq_344_out));

	wire [31:0] eq_345_in0;
	wire [31:0] eq_345_in1;
	wire [0:0] eq_345_out;
	eq #(.WIDTH(32)) eq_345(.in0(eq_345_in0), .in1(eq_345_in1), .out(eq_345_out));

	wire [31:0] eq_346_in0;
	wire [31:0] eq_346_in1;
	wire [0:0] eq_346_out;
	eq #(.WIDTH(32)) eq_346(.in0(eq_346_in0), .in1(eq_346_in1), .out(eq_346_out));

	wire [31:0] eq_347_in0;
	wire [31:0] eq_347_in1;
	wire [0:0] eq_347_out;
	eq #(.WIDTH(32)) eq_347(.in0(eq_347_in0), .in1(eq_347_in1), .out(eq_347_out));

	wire [0:0] andOp_348_in0;
	wire [0:0] andOp_348_in1;
	wire [0:0] andOp_348_out;
	andOp #(.WIDTH(1)) andOp_348(.in0(andOp_348_in0), .in1(andOp_348_in1), .out(andOp_348_out));

	wire [31:0] eq_349_in0;
	wire [31:0] eq_349_in1;
	wire [0:0] eq_349_out;
	eq #(.WIDTH(32)) eq_349(.in0(eq_349_in0), .in1(eq_349_in1), .out(eq_349_out));

	wire [31:0] eq_350_in0;
	wire [31:0] eq_350_in1;
	wire [0:0] eq_350_out;
	eq #(.WIDTH(32)) eq_350(.in0(eq_350_in0), .in1(eq_350_in1), .out(eq_350_out));

	wire [0:0] andOp_351_in0;
	wire [0:0] andOp_351_in1;
	wire [0:0] andOp_351_out;
	andOp #(.WIDTH(1)) andOp_351(.in0(andOp_351_in0), .in1(andOp_351_in1), .out(andOp_351_out));

	wire [31:0] eq_352_in0;
	wire [31:0] eq_352_in1;
	wire [0:0] eq_352_out;
	eq #(.WIDTH(32)) eq_352(.in0(eq_352_in0), .in1(eq_352_in1), .out(eq_352_out));

	wire [31:0] eq_353_in0;
	wire [31:0] eq_353_in1;
	wire [0:0] eq_353_out;
	eq #(.WIDTH(32)) eq_353(.in0(eq_353_in0), .in1(eq_353_in1), .out(eq_353_out));

	wire [31:0] eq_354_in0;
	wire [31:0] eq_354_in1;
	wire [0:0] eq_354_out;
	eq #(.WIDTH(32)) eq_354(.in0(eq_354_in0), .in1(eq_354_in1), .out(eq_354_out));

	wire [31:0] eq_355_in0;
	wire [31:0] eq_355_in1;
	wire [0:0] eq_355_out;
	eq #(.WIDTH(32)) eq_355(.in0(eq_355_in0), .in1(eq_355_in1), .out(eq_355_out));

	// End Functional Units

	reg [31:0] data_store_10_53;
	reg [31:0] data_store_10_54;
	reg [31:0] data_store_10_56;
	reg [31:0] data_store_11_58;
	reg [31:0] data_store_11_60;
	reg [31:0] data_store_11_62;
	reg [31:0] data_store_12_64;
	reg [31:0] data_store_12_66;
	reg [31:0] data_store_1_0;
	reg [31:0] data_store_1_2;
	reg [31:0] data_store_1_4;
	reg [31:0] data_store_2_10;
	reg [31:0] data_store_2_6;
	reg [31:0] data_store_2_8;
	reg [31:0] data_store_3_12;
	reg [31:0] data_store_3_14;
	reg [31:0] data_store_3_16;
	reg [31:0] data_store_4_18;
	reg [31:0] data_store_4_20;
	reg [31:0] data_store_4_22;
	reg [31:0] data_store_5_24;
	reg [31:0] data_store_5_25;
	reg [31:0] data_store_5_27;
	reg [31:0] data_store_5_29;
	reg [31:0] data_store_6_31;
	reg [31:0] data_store_6_33;
	reg [31:0] data_store_6_35;
	reg [31:0] data_store_6_37;
	reg [31:0] data_store_7_39;
	reg [31:0] data_store_7_41;
	reg [31:0] data_store_7_43;
	reg [31:0] data_store_8_45;
	reg [31:0] data_store_8_47;
	reg [31:0] data_store_9_49;
	reg [31:0] data_store_9_51;
	reg [31:0] global_state;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_10_entry_BB_reg;
	reg [0:0] state_10_is_active;
	reg [31:0] state_10_last_BB_reg;
	reg [31:0] state_10_last_state;
	reg [31:0] state_11_entry_BB_reg;
	reg [0:0] state_11_is_active;
	reg [31:0] state_11_last_BB_reg;
	reg [31:0] state_11_last_state;
	reg [31:0] state_12_entry_BB_reg;
	reg [0:0] state_12_is_active;
	reg [31:0] state_12_last_BB_reg;
	reg [31:0] state_12_last_state;
	reg [31:0] state_13_entry_BB_reg;
	reg [0:0] state_13_is_active;
	reg [31:0] state_13_last_BB_reg;
	reg [31:0] state_13_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_3_last_state;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;
	reg [31:0] state_4_last_state;
	reg [31:0] state_5_entry_BB_reg;
	reg [0:0] state_5_is_active;
	reg [31:0] state_5_last_BB_reg;
	reg [31:0] state_5_last_state;
	reg [31:0] state_6_entry_BB_reg;
	reg [0:0] state_6_is_active;
	reg [31:0] state_6_last_BB_reg;
	reg [31:0] state_6_last_state;
	reg [31:0] state_7_entry_BB_reg;
	reg [0:0] state_7_is_active;
	reg [31:0] state_7_last_BB_reg;
	reg [31:0] state_7_last_state;
	reg [31:0] state_8_entry_BB_reg;
	reg [0:0] state_8_is_active;
	reg [31:0] state_8_last_BB_reg;
	reg [31:0] state_8_last_state;
	reg [31:0] state_9_entry_BB_reg;
	reg [0:0] state_9_is_active;
	reg [31:0] state_9_last_BB_reg;
	reg [31:0] state_9_last_state;

	// controller for _____dlr_0___eq___alloca___dlr_builtin_fifo_32._____dlr_0___eq___alloca___dlr_builtin_fifo_32_in_data
	always @(*) begin
		if (andOp_243_out) begin 
			_____dlr_0___eq___alloca___dlr_builtin_fifo_32_in_data = data_in_7_42_out_data;
		end else begin
			_____dlr_0___eq___alloca___dlr_builtin_fifo_32_in_data = 0;
		end
	end
	// controller for _____dlr_0___eq___alloca___dlr_builtin_fifo_32._____dlr_0___eq___alloca___dlr_builtin_fifo_32_read_valid
	always @(*) begin
		if (andOp_246_out) begin 
			_____dlr_0___eq___alloca___dlr_builtin_fifo_32_read_valid = -(1'd1);
		end else begin
			_____dlr_0___eq___alloca___dlr_builtin_fifo_32_read_valid = 0;
		end
	end
	// controller for _____dlr_0___eq___alloca___dlr_builtin_fifo_32._____dlr_0___eq___alloca___dlr_builtin_fifo_32_write_valid
	always @(*) begin
		if (andOp_244_out) begin 
			_____dlr_0___eq___alloca___dlr_builtin_fifo_32_write_valid = -(1'd1);
		end else begin
			_____dlr_0___eq___alloca___dlr_builtin_fifo_32_write_valid = 0;
		end
	end
	// controller for add_add22.add_add22_in0
	// controller for add_add22.add_add22_in1
	// Insensitive connections
	assign add_add22_in0 = data_in_6_34_out_data;
	assign add_add22_in1 = data_in_6_32_out_data;
	// controller for add_add32.add_add32_in0
	// controller for add_add32.add_add32_in1
	// Insensitive connections
	assign add_add32_in0 = phi_phi31_out;
	assign add_add32_in1 = 32'd1;
	// controller for add_add7.add_add7_in0
	// controller for add_add7.add_add7_in1
	// Insensitive connections
	assign add_add7_in0 = phi_phi6_out;
	assign add_add7_in1 = 32'd1;
	// controller for andOp_100.andOp_100_in0
	// controller for andOp_100.andOp_100_in1
	// Insensitive connections
	assign andOp_100_in0 = bb_20_active_in_state_6_out_data;
	assign andOp_100_in1 = state_6_is_active;
	// controller for andOp_102.andOp_102_in0
	// controller for andOp_102.andOp_102_in1
	// Insensitive connections
	assign andOp_102_in0 = bb_22_active_in_state_6_out_data;
	assign andOp_102_in1 = state_6_is_active;
	// controller for andOp_104.andOp_104_in0
	// controller for andOp_104.andOp_104_in1
	// Insensitive connections
	assign andOp_104_in0 = andOp_102_out;
	assign andOp_104_in1 = _____dlr_0___eq___alloca___dlr_builtin_fifo_32_write_ready;
	// controller for andOp_106.andOp_106_in0
	// controller for andOp_106.andOp_106_in1
	// Insensitive connections
	assign andOp_106_in0 = andOp_102_out;
	assign andOp_106_in1 = notOp_105_out;
	// controller for andOp_107.andOp_107_in0
	// controller for andOp_107.andOp_107_in1
	// Insensitive connections
	assign andOp_107_in0 = bb_7_active_in_state_7_out_data;
	assign andOp_107_in1 = state_7_is_active;
	// controller for andOp_109.andOp_109_in0
	// controller for andOp_109.andOp_109_in1
	// Insensitive connections
	assign andOp_109_in0 = andOp_107_out;
	assign andOp_109_in1 = icmp_icmp26_out;
	// controller for andOp_111.andOp_111_in0
	// controller for andOp_111.andOp_111_in1
	// Insensitive connections
	assign andOp_111_in0 = andOp_107_out;
	assign andOp_111_in1 = notOp_110_out;
	// controller for andOp_112.andOp_112_in0
	// controller for andOp_112.andOp_112_in1
	// Insensitive connections
	assign andOp_112_in0 = bb_23_active_in_state_7_out_data;
	assign andOp_112_in1 = state_7_is_active;
	// controller for andOp_114.andOp_114_in0
	// controller for andOp_114.andOp_114_in1
	// Insensitive connections
	assign andOp_114_in0 = bb_1_active_in_state_8_out_data;
	assign andOp_114_in1 = state_8_is_active;
	// controller for andOp_116.andOp_116_in0
	// controller for andOp_116.andOp_116_in1
	// Insensitive connections
	assign andOp_116_in0 = bb_9_active_in_state_8_out_data;
	assign andOp_116_in1 = state_8_is_active;
	// controller for andOp_118.andOp_118_in0
	// controller for andOp_118.andOp_118_in1
	// Insensitive connections
	assign andOp_118_in0 = bb_10_active_in_state_8_out_data;
	assign andOp_118_in1 = state_8_is_active;
	// controller for andOp_120.andOp_120_in0
	// controller for andOp_120.andOp_120_in1
	// Insensitive connections
	assign andOp_120_in0 = andOp_118_out;
	assign andOp_120_in1 = _____dlr_0___eq___alloca___dlr_builtin_fifo_32_read_ready;
	// controller for andOp_122.andOp_122_in0
	// controller for andOp_122.andOp_122_in1
	// Insensitive connections
	assign andOp_122_in0 = andOp_118_out;
	assign andOp_122_in1 = notOp_121_out;
	// controller for andOp_123.andOp_123_in0
	// controller for andOp_123.andOp_123_in1
	// Insensitive connections
	assign andOp_123_in0 = bb_11_active_in_state_10_out_data;
	assign andOp_123_in1 = state_10_is_active;
	// controller for andOp_125.andOp_125_in0
	// controller for andOp_125.andOp_125_in1
	// Insensitive connections
	assign andOp_125_in0 = bb_11_active_in_state_10_out_data;
	assign andOp_125_in1 = state_10_is_active;
	// controller for andOp_127.andOp_127_in0
	// controller for andOp_127.andOp_127_in1
	// Insensitive connections
	assign andOp_127_in0 = bb_12_active_in_state_11_out_data;
	assign andOp_127_in1 = state_11_is_active;
	// controller for andOp_129.andOp_129_in0
	// controller for andOp_129.andOp_129_in1
	// Insensitive connections
	assign andOp_129_in0 = bb_13_active_in_state_11_out_data;
	assign andOp_129_in1 = state_11_is_active;
	// controller for andOp_131.andOp_131_in0
	// controller for andOp_131.andOp_131_in1
	// Insensitive connections
	assign andOp_131_in0 = andOp_129_out;
	assign andOp_131_in1 = arg_2_write_ready;
	// controller for andOp_133.andOp_133_in0
	// controller for andOp_133.andOp_133_in1
	// Insensitive connections
	assign andOp_133_in0 = andOp_129_out;
	assign andOp_133_in1 = notOp_132_out;
	// controller for andOp_134.andOp_134_in0
	// controller for andOp_134.andOp_134_in1
	// Insensitive connections
	assign andOp_134_in0 = bb_2_active_in_state_11_out_data;
	assign andOp_134_in1 = state_11_is_active;
	// controller for andOp_136.andOp_136_in0
	// controller for andOp_136.andOp_136_in1
	// Insensitive connections
	assign andOp_136_in0 = bb_3_active_in_state_12_out_data;
	assign andOp_136_in1 = state_12_is_active;
	// controller for andOp_138.andOp_138_in0
	// controller for andOp_138.andOp_138_in1
	// Insensitive connections
	assign andOp_138_in0 = andOp_136_out;
	assign andOp_138_in1 = icmp_icmp45_out;
	// controller for andOp_140.andOp_140_in0
	// controller for andOp_140.andOp_140_in1
	// Insensitive connections
	assign andOp_140_in0 = andOp_136_out;
	assign andOp_140_in1 = notOp_139_out;
	// controller for andOp_141.andOp_141_in0
	// controller for andOp_141.andOp_141_in1
	// Insensitive connections
	assign andOp_141_in0 = bb_14_active_in_state_12_out_data;
	assign andOp_141_in1 = state_12_is_active;
	// controller for andOp_188.andOp_188_in0
	// controller for andOp_188.andOp_188_in1
	// Insensitive connections
	assign andOp_188_in0 = notOp_187_out;
	assign andOp_188_in1 = andOp_75_out;
	// controller for andOp_191.andOp_191_in0
	// controller for andOp_191.andOp_191_in1
	// Insensitive connections
	assign andOp_191_in0 = notOp_190_out;
	assign andOp_191_in1 = andOp_77_out;
	// controller for andOp_196.andOp_196_in0
	// controller for andOp_196.andOp_196_in1
	// Insensitive connections
	assign andOp_196_in0 = notOp_195_out;
	assign andOp_196_in1 = andOp_85_out;
	// controller for andOp_200.andOp_200_in0
	// controller for andOp_200.andOp_200_in1
	// Insensitive connections
	assign andOp_200_in0 = notOp_199_out;
	assign andOp_200_in1 = andOp_79_out;
	// controller for andOp_203.andOp_203_in0
	// controller for andOp_203.andOp_203_in1
	// Insensitive connections
	assign andOp_203_in0 = notOp_202_out;
	assign andOp_203_in1 = andOp_81_out;
	// controller for andOp_208.andOp_208_in0
	// controller for andOp_208.andOp_208_in1
	// Insensitive connections
	assign andOp_208_in0 = notOp_207_out;
	assign andOp_208_in1 = andOp_98_out;
	// controller for andOp_211.andOp_211_in0
	// controller for andOp_211.andOp_211_in1
	// Insensitive connections
	assign andOp_211_in0 = notOp_210_out;
	assign andOp_211_in1 = andOp_92_out;
	// controller for andOp_215.andOp_215_in0
	// controller for andOp_215.andOp_215_in1
	// Insensitive connections
	assign andOp_215_in0 = notOp_214_out;
	assign andOp_215_in1 = andOp_96_out;
	// controller for andOp_218.andOp_218_in0
	// controller for andOp_218.andOp_218_in1
	// Insensitive connections
	assign andOp_218_in0 = notOp_217_out;
	assign andOp_218_in1 = andOp_112_out;
	// controller for andOp_223.andOp_223_in0
	// controller for andOp_223.andOp_223_in1
	// Insensitive connections
	assign andOp_223_in0 = notOp_222_out;
	assign andOp_223_in1 = andOp_114_out;
	// controller for andOp_226.andOp_226_in0
	// controller for andOp_226.andOp_226_in1
	// Insensitive connections
	assign andOp_226_in0 = notOp_225_out;
	assign andOp_226_in1 = andOp_116_out;
	// controller for andOp_231.andOp_231_in0
	// controller for andOp_231.andOp_231_in1
	// Insensitive connections
	assign andOp_231_in0 = notOp_230_out;
	assign andOp_231_in1 = andOp_134_out;
	// controller for andOp_234.andOp_234_in0
	// controller for andOp_234.andOp_234_in1
	// Insensitive connections
	assign andOp_234_in0 = notOp_233_out;
	assign andOp_234_in1 = andOp_127_out;
	// controller for andOp_238.andOp_238_in0
	// controller for andOp_238.andOp_238_in1
	// Insensitive connections
	assign andOp_238_in0 = notOp_237_out;
	assign andOp_238_in1 = andOp_141_out;
	// controller for andOp_241.andOp_241_in0
	// controller for andOp_241.andOp_241_in1
	// Insensitive connections
	assign andOp_241_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_241_in1 = state_0_is_active;
	// controller for andOp_242.andOp_242_in0
	// controller for andOp_242.andOp_242_in1
	// Insensitive connections
	assign andOp_242_in0 = bb_22_active_in_state_6_out_data;
	assign andOp_242_in1 = state_6_is_active;
	// controller for andOp_243.andOp_243_in0
	// controller for andOp_243.andOp_243_in1
	// Insensitive connections
	assign andOp_243_in0 = bb_23_active_in_state_7_out_data;
	assign andOp_243_in1 = state_7_is_active;
	// controller for andOp_244.andOp_244_in0
	// controller for andOp_244.andOp_244_in1
	// Insensitive connections
	assign andOp_244_in0 = bb_23_active_in_state_7_out_data;
	assign andOp_244_in1 = state_7_is_active;
	// controller for andOp_245.andOp_245_in0
	// controller for andOp_245.andOp_245_in1
	// Insensitive connections
	assign andOp_245_in0 = bb_10_active_in_state_8_out_data;
	assign andOp_245_in1 = state_8_is_active;
	// controller for andOp_246.andOp_246_in0
	// controller for andOp_246.andOp_246_in1
	// Insensitive connections
	assign andOp_246_in0 = bb_11_active_in_state_9_out_data;
	assign andOp_246_in1 = state_9_is_active;
	// controller for andOp_247.andOp_247_in0
	// controller for andOp_247.andOp_247_in1
	// Insensitive connections
	assign andOp_247_in0 = bb_11_active_in_state_10_out_data;
	assign andOp_247_in1 = state_10_is_active;
	// controller for andOp_248.andOp_248_in0
	// controller for andOp_248.andOp_248_in1
	// Insensitive connections
	assign andOp_248_in0 = bb_16_active_in_state_1_out_data;
	assign andOp_248_in1 = state_1_is_active;
	// controller for andOp_249.andOp_249_in0
	// controller for andOp_249.andOp_249_in1
	// Insensitive connections
	assign andOp_249_in0 = bb_17_active_in_state_2_out_data;
	assign andOp_249_in1 = state_2_is_active;
	// controller for andOp_250.andOp_250_in0
	// controller for andOp_250.andOp_250_in1
	// Insensitive connections
	assign andOp_250_in0 = bb_17_active_in_state_3_out_data;
	assign andOp_250_in1 = state_3_is_active;
	// controller for andOp_251.andOp_251_in0
	// controller for andOp_251.andOp_251_in1
	// Insensitive connections
	assign andOp_251_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_251_in1 = state_1_is_active;
	// controller for andOp_254.andOp_254_in0
	// controller for andOp_254.andOp_254_in1
	// Insensitive connections
	assign andOp_254_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_254_in1 = state_1_is_active;
	// controller for andOp_255.andOp_255_in0
	// controller for andOp_255.andOp_255_in1
	// Insensitive connections
	assign andOp_255_in0 = bb_19_active_in_state_3_out_data;
	assign andOp_255_in1 = state_3_is_active;
	// controller for andOp_256.andOp_256_in0
	// controller for andOp_256.andOp_256_in1
	// Insensitive connections
	assign andOp_256_in0 = bb_20_active_in_state_4_out_data;
	assign andOp_256_in1 = state_4_is_active;
	// controller for andOp_257.andOp_257_in0
	// controller for andOp_257.andOp_257_in1
	// Insensitive connections
	assign andOp_257_in0 = bb_20_active_in_state_5_out_data;
	assign andOp_257_in1 = state_5_is_active;
	// controller for andOp_258.andOp_258_in0
	// controller for andOp_258.andOp_258_in1
	// Insensitive connections
	assign andOp_258_in0 = bb_6_active_in_state_6_out_data;
	assign andOp_258_in1 = state_6_is_active;
	// controller for andOp_259.andOp_259_in0
	// controller for andOp_259.andOp_259_in1
	// Insensitive connections
	assign andOp_259_in0 = bb_7_active_in_state_7_out_data;
	assign andOp_259_in1 = state_7_is_active;
	// controller for andOp_260.andOp_260_in0
	// controller for andOp_260.andOp_260_in1
	// Insensitive connections
	assign andOp_260_in0 = bb_1_active_in_state_8_out_data;
	assign andOp_260_in1 = state_8_is_active;
	// controller for andOp_263.andOp_263_in0
	// controller for andOp_263.andOp_263_in1
	// Insensitive connections
	assign andOp_263_in0 = bb_1_active_in_state_8_out_data;
	assign andOp_263_in1 = state_8_is_active;
	// controller for andOp_264.andOp_264_in0
	// controller for andOp_264.andOp_264_in1
	// Insensitive connections
	assign andOp_264_in0 = bb_13_active_in_state_11_out_data;
	assign andOp_264_in1 = state_11_is_active;
	// controller for andOp_265.andOp_265_in0
	// controller for andOp_265.andOp_265_in1
	// Insensitive connections
	assign andOp_265_in0 = bb_14_active_in_state_12_out_data;
	assign andOp_265_in1 = state_12_is_active;
	// controller for andOp_266.andOp_266_in0
	// controller for andOp_266.andOp_266_in1
	// Insensitive connections
	assign andOp_266_in0 = bb_14_active_in_state_12_out_data;
	assign andOp_266_in1 = state_12_is_active;
	// controller for andOp_267.andOp_267_in0
	// controller for andOp_267.andOp_267_in1
	// Insensitive connections
	assign andOp_267_in0 = bb_2_active_in_state_11_out_data;
	assign andOp_267_in1 = state_11_is_active;
	// controller for andOp_268.andOp_268_in0
	// controller for andOp_268.andOp_268_in1
	// Insensitive connections
	assign andOp_268_in0 = bb_3_active_in_state_12_out_data;
	assign andOp_268_in1 = state_12_is_active;
	// controller for andOp_269.andOp_269_in0
	// controller for andOp_269.andOp_269_in1
	// Insensitive connections
	assign andOp_269_in0 = bb_8_active_in_state_13_out_data;
	assign andOp_269_in1 = state_13_is_active;
	// controller for andOp_270.andOp_270_in0
	// controller for andOp_270.andOp_270_in1
	// Insensitive connections
	assign andOp_270_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_270_in1 = state_0_is_active;
	// controller for andOp_271.andOp_271_in0
	// controller for andOp_271.andOp_271_in1
	// Insensitive connections
	assign andOp_271_in0 = bb_17_active_in_state_2_out_data;
	assign andOp_271_in1 = state_2_is_active;
	// controller for andOp_272.andOp_272_in0
	// controller for andOp_272.andOp_272_in1
	// Insensitive connections
	assign andOp_272_in0 = bb_20_active_in_state_4_out_data;
	assign andOp_272_in1 = state_4_is_active;
	// controller for andOp_273.andOp_273_in0
	// controller for andOp_273.andOp_273_in1
	// Insensitive connections
	assign andOp_273_in0 = bb_20_active_in_state_5_out_data;
	assign andOp_273_in1 = state_5_is_active;
	// controller for andOp_274.andOp_274_in0
	// controller for andOp_274.andOp_274_in1
	// Insensitive connections
	assign andOp_274_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_274_in1 = state_0_is_active;
	// controller for andOp_275.andOp_275_in0
	// controller for andOp_275.andOp_275_in1
	// Insensitive connections
	assign andOp_275_in0 = bb_11_active_in_state_9_out_data;
	assign andOp_275_in1 = state_9_is_active;
	// controller for andOp_276.andOp_276_in0
	// controller for andOp_276.andOp_276_in1
	// Insensitive connections
	assign andOp_276_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_276_in1 = state_0_is_active;
	// controller for andOp_277.andOp_277_in0
	// controller for andOp_277.andOp_277_in1
	// Insensitive connections
	assign andOp_277_in0 = bb_8_active_in_state_13_out_data;
	assign andOp_277_in1 = state_13_is_active;
	// controller for andOp_279.andOp_279_in0
	// controller for andOp_279.andOp_279_in1
	// Insensitive connections
	assign andOp_279_in0 = notOp_278_out;
	assign andOp_279_in1 = 1'd1;
	// controller for andOp_281.andOp_281_in0
	// controller for andOp_281.andOp_281_in1
	// Insensitive connections
	assign andOp_281_in0 = notOp_280_out;
	assign andOp_281_in1 = andOp_279_out;
	// controller for andOp_283.andOp_283_in0
	// controller for andOp_283.andOp_283_in1
	// Insensitive connections
	assign andOp_283_in0 = notOp_282_out;
	assign andOp_283_in1 = andOp_281_out;
	// controller for andOp_285.andOp_285_in0
	// controller for andOp_285.andOp_285_in1
	// Insensitive connections
	assign andOp_285_in0 = notOp_284_out;
	assign andOp_285_in1 = 1'd1;
	// controller for andOp_287.andOp_287_in0
	// controller for andOp_287.andOp_287_in1
	// Insensitive connections
	assign andOp_287_in0 = notOp_286_out;
	assign andOp_287_in1 = 1'd1;
	// controller for andOp_289.andOp_289_in0
	// controller for andOp_289.andOp_289_in1
	// Insensitive connections
	assign andOp_289_in0 = notOp_288_out;
	assign andOp_289_in1 = andOp_287_out;
	// controller for andOp_291.andOp_291_in0
	// controller for andOp_291.andOp_291_in1
	// Insensitive connections
	assign andOp_291_in0 = notOp_290_out;
	assign andOp_291_in1 = 1'd1;
	// controller for andOp_293.andOp_293_in0
	// controller for andOp_293.andOp_293_in1
	// Insensitive connections
	assign andOp_293_in0 = notOp_292_out;
	assign andOp_293_in1 = 1'd1;
	// controller for andOp_295.andOp_295_in0
	// controller for andOp_295.andOp_295_in1
	// Insensitive connections
	assign andOp_295_in0 = notOp_294_out;
	assign andOp_295_in1 = 1'd1;
	// controller for andOp_297.andOp_297_in0
	// controller for andOp_297.andOp_297_in1
	// Insensitive connections
	assign andOp_297_in0 = notOp_296_out;
	assign andOp_297_in1 = andOp_295_out;
	// controller for andOp_299.andOp_299_in0
	// controller for andOp_299.andOp_299_in1
	// Insensitive connections
	assign andOp_299_in0 = notOp_298_out;
	assign andOp_299_in1 = 1'd1;
	// controller for andOp_301.andOp_301_in0
	// controller for andOp_301.andOp_301_in1
	// Insensitive connections
	assign andOp_301_in0 = notOp_300_out;
	assign andOp_301_in1 = 1'd1;
	// controller for andOp_303.andOp_303_in0
	// controller for andOp_303.andOp_303_in1
	// Insensitive connections
	assign andOp_303_in0 = notOp_302_out;
	assign andOp_303_in1 = andOp_301_out;
	// controller for andOp_305.andOp_305_in0
	// controller for andOp_305.andOp_305_in1
	// Insensitive connections
	assign andOp_305_in0 = notOp_304_out;
	assign andOp_305_in1 = andOp_303_out;
	// controller for andOp_307.andOp_307_in0
	// controller for andOp_307.andOp_307_in1
	// Insensitive connections
	assign andOp_307_in0 = notOp_306_out;
	assign andOp_307_in1 = 1'd1;
	// controller for andOp_309.andOp_309_in0
	// controller for andOp_309.andOp_309_in1
	// Insensitive connections
	assign andOp_309_in0 = notOp_308_out;
	assign andOp_309_in1 = 1'd1;
	// controller for andOp_311.andOp_311_in0
	// controller for andOp_311.andOp_311_in1
	// Insensitive connections
	assign andOp_311_in0 = notOp_310_out;
	assign andOp_311_in1 = 1'd1;
	// controller for andOp_313.andOp_313_in0
	// controller for andOp_313.andOp_313_in1
	// Insensitive connections
	assign andOp_313_in0 = notOp_312_out;
	assign andOp_313_in1 = andOp_311_out;
	// controller for andOp_315.andOp_315_in0
	// controller for andOp_315.andOp_315_in1
	// Insensitive connections
	assign andOp_315_in0 = notOp_314_out;
	assign andOp_315_in1 = 1'd1;
	// controller for andOp_317.andOp_317_in0
	// controller for andOp_317.andOp_317_in1
	// Insensitive connections
	assign andOp_317_in0 = notOp_316_out;
	assign andOp_317_in1 = 1'd1;
	// controller for andOp_319.andOp_319_in0
	// controller for andOp_319.andOp_319_in1
	// Insensitive connections
	assign andOp_319_in0 = notOp_318_out;
	assign andOp_319_in1 = andOp_317_out;
	// controller for andOp_324.andOp_324_in0
	// controller for andOp_324.andOp_324_in1
	// Insensitive connections
	assign andOp_324_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_324_in1 = state_1_is_active;
	// controller for andOp_329.andOp_329_in0
	// controller for andOp_329.andOp_329_in1
	// Insensitive connections
	assign andOp_329_in0 = bb_17_active_in_state_3_out_data;
	assign andOp_329_in1 = state_3_is_active;
	// controller for andOp_334.andOp_334_in0
	// controller for andOp_334.andOp_334_in1
	// Insensitive connections
	assign andOp_334_in0 = bb_20_active_in_state_5_out_data;
	assign andOp_334_in1 = state_5_is_active;
	// controller for andOp_337.andOp_337_in0
	// controller for andOp_337.andOp_337_in1
	// Insensitive connections
	assign andOp_337_in0 = bb_6_active_in_state_6_out_data;
	assign andOp_337_in1 = state_6_is_active;
	// controller for andOp_343.andOp_343_in0
	// controller for andOp_343.andOp_343_in1
	// Insensitive connections
	assign andOp_343_in0 = bb_1_active_in_state_8_out_data;
	assign andOp_343_in1 = state_8_is_active;
	// controller for andOp_348.andOp_348_in0
	// controller for andOp_348.andOp_348_in1
	// Insensitive connections
	assign andOp_348_in0 = bb_11_active_in_state_10_out_data;
	assign andOp_348_in1 = state_10_is_active;
	// controller for andOp_351.andOp_351_in0
	// controller for andOp_351.andOp_351_in1
	// Insensitive connections
	assign andOp_351_in0 = bb_2_active_in_state_11_out_data;
	assign andOp_351_in1 = state_11_is_active;
	// controller for andOp_68.andOp_68_in0
	// controller for andOp_68.andOp_68_in1
	// Insensitive connections
	assign andOp_68_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_68_in1 = state_0_is_active;
	// controller for andOp_70.andOp_70_in0
	// controller for andOp_70.andOp_70_in1
	// Insensitive connections
	assign andOp_70_in0 = bb_16_active_in_state_1_out_data;
	assign andOp_70_in1 = state_1_is_active;
	// controller for andOp_72.andOp_72_in0
	// controller for andOp_72.andOp_72_in1
	// Insensitive connections
	assign andOp_72_in0 = andOp_70_out;
	assign andOp_72_in1 = arg_0_read_ready;
	// controller for andOp_74.andOp_74_in0
	// controller for andOp_74.andOp_74_in1
	// Insensitive connections
	assign andOp_74_in0 = andOp_70_out;
	assign andOp_74_in1 = notOp_73_out;
	// controller for andOp_75.andOp_75_in0
	// controller for andOp_75.andOp_75_in1
	// Insensitive connections
	assign andOp_75_in0 = bb_15_active_in_state_1_out_data;
	assign andOp_75_in1 = state_1_is_active;
	// controller for andOp_77.andOp_77_in0
	// controller for andOp_77.andOp_77_in1
	// Insensitive connections
	assign andOp_77_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_77_in1 = state_1_is_active;
	// controller for andOp_79.andOp_79_in0
	// controller for andOp_79.andOp_79_in1
	// Insensitive connections
	assign andOp_79_in0 = bb_17_active_in_state_3_out_data;
	assign andOp_79_in1 = state_3_is_active;
	// controller for andOp_81.andOp_81_in0
	// controller for andOp_81.andOp_81_in1
	// Insensitive connections
	assign andOp_81_in0 = bb_18_active_in_state_3_out_data;
	assign andOp_81_in1 = state_3_is_active;
	// controller for andOp_83.andOp_83_in0
	// controller for andOp_83.andOp_83_in1
	// Insensitive connections
	assign andOp_83_in0 = bb_17_active_in_state_3_out_data;
	assign andOp_83_in1 = state_3_is_active;
	// controller for andOp_85.andOp_85_in0
	// controller for andOp_85.andOp_85_in1
	// Insensitive connections
	assign andOp_85_in0 = bb_5_active_in_state_3_out_data;
	assign andOp_85_in1 = state_3_is_active;
	// controller for andOp_87.andOp_87_in0
	// controller for andOp_87.andOp_87_in1
	// Insensitive connections
	assign andOp_87_in0 = bb_19_active_in_state_3_out_data;
	assign andOp_87_in1 = state_3_is_active;
	// controller for andOp_89.andOp_89_in0
	// controller for andOp_89.andOp_89_in1
	// Insensitive connections
	assign andOp_89_in0 = andOp_87_out;
	assign andOp_89_in1 = arg_1_read_ready;
	// controller for andOp_91.andOp_91_in0
	// controller for andOp_91.andOp_91_in1
	// Insensitive connections
	assign andOp_91_in0 = andOp_87_out;
	assign andOp_91_in1 = notOp_90_out;
	// controller for andOp_92.andOp_92_in0
	// controller for andOp_92.andOp_92_in1
	// Insensitive connections
	assign andOp_92_in0 = bb_20_active_in_state_6_out_data;
	assign andOp_92_in1 = state_6_is_active;
	// controller for andOp_94.andOp_94_in0
	// controller for andOp_94.andOp_94_in1
	// Insensitive connections
	assign andOp_94_in0 = bb_20_active_in_state_6_out_data;
	assign andOp_94_in1 = state_6_is_active;
	// controller for andOp_96.andOp_96_in0
	// controller for andOp_96.andOp_96_in1
	// Insensitive connections
	assign andOp_96_in0 = bb_21_active_in_state_6_out_data;
	assign andOp_96_in1 = state_6_is_active;
	// controller for andOp_98.andOp_98_in0
	// controller for andOp_98.andOp_98_in1
	// Insensitive connections
	assign andOp_98_in0 = bb_6_active_in_state_6_out_data;
	assign andOp_98_in1 = state_6_is_active;
	// controller for arg_0.arg_0_read_valid_reg
	always @(*) begin
		if (andOp_249_out) begin 
			arg_0_read_valid_reg = -(1'd1);
		end else begin
			arg_0_read_valid_reg = 0;
		end
	end
	// controller for arg_1.arg_1_read_valid_reg
	always @(*) begin
		if (andOp_256_out) begin 
			arg_1_read_valid_reg = -(1'd1);
		end else begin
			arg_1_read_valid_reg = 0;
		end
	end
	// controller for arg_2.arg_2_in_data_reg
	always @(*) begin
		if (andOp_266_out) begin 
			arg_2_in_data_reg = data_in_12_67_out_data;
		end else begin
			arg_2_in_data_reg = 0;
		end
	end
	// controller for arg_2.arg_2_write_valid_reg
	always @(*) begin
		if (andOp_265_out) begin 
			arg_2_write_valid_reg = -(1'd1);
		end else begin
			arg_2_write_valid_reg = 0;
		end
	end
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_143_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_185_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_8.bb_10_active_in_state_8_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_8_in_data = orOp_173_out;
		end else begin
			bb_10_active_in_state_8_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_8.bb_10_predecessor_in_state_8_in_data
	always @(*) begin
		if (andOp_226_out) begin 
			bb_10_predecessor_in_state_8_in_data = 32'd9;
		end else if (eq_224_out) begin 
			bb_10_predecessor_in_state_8_in_data = state_8_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_8_in_data = 0;
		end
	end
	// controller for bb_11_active_in_state_10.bb_11_active_in_state_10_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_11_active_in_state_10_in_data = eq_175_out;
		end else begin
			bb_11_active_in_state_10_in_data = 0;
		end
	end
	// controller for bb_11_active_in_state_9.bb_11_active_in_state_9_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_11_active_in_state_9_in_data = eq_174_out;
		end else begin
			bb_11_active_in_state_9_in_data = 0;
		end
	end
	// controller for bb_11_predecessor_in_state_10.bb_11_predecessor_in_state_10_in_data
	always @(*) begin
		if (eq_228_out) begin 
			bb_11_predecessor_in_state_10_in_data = state_10_last_BB_reg;
		end else begin
			bb_11_predecessor_in_state_10_in_data = 0;
		end
	end
	// controller for bb_11_predecessor_in_state_9.bb_11_predecessor_in_state_9_in_data
	always @(*) begin
		if (eq_227_out) begin 
			bb_11_predecessor_in_state_9_in_data = state_9_last_BB_reg;
		end else begin
			bb_11_predecessor_in_state_9_in_data = 0;
		end
	end
	// controller for bb_12_active_in_state_11.bb_12_active_in_state_11_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_12_active_in_state_11_in_data = orOp_177_out;
		end else begin
			bb_12_active_in_state_11_in_data = 0;
		end
	end
	// controller for bb_12_predecessor_in_state_11.bb_12_predecessor_in_state_11_in_data
	always @(*) begin
		if (andOp_231_out) begin 
			bb_12_predecessor_in_state_11_in_data = 32'd2;
		end else if (eq_229_out) begin 
			bb_12_predecessor_in_state_11_in_data = state_11_last_BB_reg;
		end else begin
			bb_12_predecessor_in_state_11_in_data = 0;
		end
	end
	// controller for bb_13_active_in_state_11.bb_13_active_in_state_11_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_13_active_in_state_11_in_data = orOp_179_out;
		end else begin
			bb_13_active_in_state_11_in_data = 0;
		end
	end
	// controller for bb_13_predecessor_in_state_11.bb_13_predecessor_in_state_11_in_data
	always @(*) begin
		if (andOp_234_out) begin 
			bb_13_predecessor_in_state_11_in_data = 32'd12;
		end else if (eq_232_out) begin 
			bb_13_predecessor_in_state_11_in_data = state_11_last_BB_reg;
		end else begin
			bb_13_predecessor_in_state_11_in_data = 0;
		end
	end
	// controller for bb_14_active_in_state_12.bb_14_active_in_state_12_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_14_active_in_state_12_in_data = eq_183_out;
		end else begin
			bb_14_active_in_state_12_in_data = 0;
		end
	end
	// controller for bb_14_predecessor_in_state_12.bb_14_predecessor_in_state_12_in_data
	always @(*) begin
		if (eq_239_out) begin 
			bb_14_predecessor_in_state_12_in_data = state_12_last_BB_reg;
		end else begin
			bb_14_predecessor_in_state_12_in_data = 0;
		end
	end
	// controller for bb_15_active_in_state_1.bb_15_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_15_active_in_state_1_in_data = orOp_147_out;
		end else begin
			bb_15_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_15_predecessor_in_state_1.bb_15_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_191_out) begin 
			bb_15_predecessor_in_state_1_in_data = 32'd4;
		end else if (eq_189_out) begin 
			bb_15_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_15_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_16_active_in_state_1.bb_16_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_16_active_in_state_1_in_data = orOp_145_out;
		end else begin
			bb_16_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_16_predecessor_in_state_1.bb_16_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_188_out) begin 
			bb_16_predecessor_in_state_1_in_data = 32'd15;
		end else if (eq_186_out) begin 
			bb_16_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_16_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_17_active_in_state_2.bb_17_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_17_active_in_state_2_in_data = eq_149_out;
		end else begin
			bb_17_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_17_active_in_state_3.bb_17_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_17_active_in_state_3_in_data = eq_152_out;
		end else begin
			bb_17_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_17_predecessor_in_state_2.bb_17_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_193_out) begin 
			bb_17_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_17_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_17_predecessor_in_state_3.bb_17_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_197_out) begin 
			bb_17_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_17_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_18_active_in_state_3.bb_18_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_18_active_in_state_3_in_data = orOp_151_out;
		end else begin
			bb_18_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_18_predecessor_in_state_3.bb_18_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_196_out) begin 
			bb_18_predecessor_in_state_3_in_data = 32'd5;
		end else if (eq_194_out) begin 
			bb_18_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_18_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_19_active_in_state_3.bb_19_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_19_active_in_state_3_in_data = orOp_156_out;
		end else begin
			bb_19_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_19_predecessor_in_state_3.bb_19_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_203_out) begin 
			bb_19_predecessor_in_state_3_in_data = 32'd18;
		end else if (eq_201_out) begin 
			bb_19_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_19_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_8.bb_1_active_in_state_8_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_8_in_data = eq_169_out;
		end else begin
			bb_1_active_in_state_8_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_8.bb_1_predecessor_in_state_8_in_data
	always @(*) begin
		if (eq_220_out) begin 
			bb_1_predecessor_in_state_8_in_data = state_8_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_8_in_data = 0;
		end
	end
	// controller for bb_20_active_in_state_4.bb_20_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_20_active_in_state_4_in_data = eq_157_out;
		end else begin
			bb_20_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_20_active_in_state_5.bb_20_active_in_state_5_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_20_active_in_state_5_in_data = eq_158_out;
		end else begin
			bb_20_active_in_state_5_in_data = 0;
		end
	end
	// controller for bb_20_active_in_state_6.bb_20_active_in_state_6_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_20_active_in_state_6_in_data = eq_163_out;
		end else begin
			bb_20_active_in_state_6_in_data = 0;
		end
	end
	// controller for bb_20_predecessor_in_state_4.bb_20_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_204_out) begin 
			bb_20_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_20_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_20_predecessor_in_state_5.bb_20_predecessor_in_state_5_in_data
	always @(*) begin
		if (eq_205_out) begin 
			bb_20_predecessor_in_state_5_in_data = state_5_last_BB_reg;
		end else begin
			bb_20_predecessor_in_state_5_in_data = 0;
		end
	end
	// controller for bb_20_predecessor_in_state_6.bb_20_predecessor_in_state_6_in_data
	always @(*) begin
		if (eq_212_out) begin 
			bb_20_predecessor_in_state_6_in_data = state_6_last_BB_reg;
		end else begin
			bb_20_predecessor_in_state_6_in_data = 0;
		end
	end
	// controller for bb_21_active_in_state_6.bb_21_active_in_state_6_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_21_active_in_state_6_in_data = orOp_160_out;
		end else begin
			bb_21_active_in_state_6_in_data = 0;
		end
	end
	// controller for bb_21_predecessor_in_state_6.bb_21_predecessor_in_state_6_in_data
	always @(*) begin
		if (andOp_208_out) begin 
			bb_21_predecessor_in_state_6_in_data = 32'd6;
		end else if (eq_206_out) begin 
			bb_21_predecessor_in_state_6_in_data = state_6_last_BB_reg;
		end else begin
			bb_21_predecessor_in_state_6_in_data = 0;
		end
	end
	// controller for bb_22_active_in_state_6.bb_22_active_in_state_6_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_22_active_in_state_6_in_data = orOp_165_out;
		end else begin
			bb_22_active_in_state_6_in_data = 0;
		end
	end
	// controller for bb_22_predecessor_in_state_6.bb_22_predecessor_in_state_6_in_data
	always @(*) begin
		if (andOp_215_out) begin 
			bb_22_predecessor_in_state_6_in_data = 32'd21;
		end else if (eq_213_out) begin 
			bb_22_predecessor_in_state_6_in_data = state_6_last_BB_reg;
		end else begin
			bb_22_predecessor_in_state_6_in_data = 0;
		end
	end
	// controller for bb_23_active_in_state_7.bb_23_active_in_state_7_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_23_active_in_state_7_in_data = eq_168_out;
		end else begin
			bb_23_active_in_state_7_in_data = 0;
		end
	end
	// controller for bb_23_predecessor_in_state_7.bb_23_predecessor_in_state_7_in_data
	always @(*) begin
		if (eq_219_out) begin 
			bb_23_predecessor_in_state_7_in_data = state_7_last_BB_reg;
		end else begin
			bb_23_predecessor_in_state_7_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_11.bb_2_active_in_state_11_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_11_in_data = eq_180_out;
		end else begin
			bb_2_active_in_state_11_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_11.bb_2_predecessor_in_state_11_in_data
	always @(*) begin
		if (eq_235_out) begin 
			bb_2_predecessor_in_state_11_in_data = state_11_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_11_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_12.bb_3_active_in_state_12_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_12_in_data = orOp_182_out;
		end else begin
			bb_3_active_in_state_12_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_12.bb_3_predecessor_in_state_12_in_data
	always @(*) begin
		if (andOp_238_out) begin 
			bb_3_predecessor_in_state_12_in_data = 32'd14;
		end else if (eq_236_out) begin 
			bb_3_predecessor_in_state_12_in_data = state_12_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_12_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_1.bb_4_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_1_in_data = eq_148_out;
		end else begin
			bb_4_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_1.bb_4_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_192_out) begin 
			bb_4_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_5_active_in_state_3.bb_5_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_5_active_in_state_3_in_data = orOp_154_out;
		end else begin
			bb_5_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_5_predecessor_in_state_3.bb_5_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_200_out) begin 
			bb_5_predecessor_in_state_3_in_data = 32'd17;
		end else if (eq_198_out) begin 
			bb_5_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_5_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_6_active_in_state_6.bb_6_active_in_state_6_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_6_active_in_state_6_in_data = orOp_162_out;
		end else begin
			bb_6_active_in_state_6_in_data = 0;
		end
	end
	// controller for bb_6_predecessor_in_state_6.bb_6_predecessor_in_state_6_in_data
	always @(*) begin
		if (andOp_211_out) begin 
			bb_6_predecessor_in_state_6_in_data = 32'd20;
		end else if (eq_209_out) begin 
			bb_6_predecessor_in_state_6_in_data = state_6_last_BB_reg;
		end else begin
			bb_6_predecessor_in_state_6_in_data = 0;
		end
	end
	// controller for bb_7_active_in_state_7.bb_7_active_in_state_7_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_7_active_in_state_7_in_data = orOp_167_out;
		end else begin
			bb_7_active_in_state_7_in_data = 0;
		end
	end
	// controller for bb_7_predecessor_in_state_7.bb_7_predecessor_in_state_7_in_data
	always @(*) begin
		if (andOp_218_out) begin 
			bb_7_predecessor_in_state_7_in_data = 32'd23;
		end else if (eq_216_out) begin 
			bb_7_predecessor_in_state_7_in_data = state_7_last_BB_reg;
		end else begin
			bb_7_predecessor_in_state_7_in_data = 0;
		end
	end
	// controller for bb_8_active_in_state_13.bb_8_active_in_state_13_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_state_13_in_data = eq_184_out;
		end else begin
			bb_8_active_in_state_13_in_data = 0;
		end
	end
	// controller for bb_8_predecessor_in_state_13.bb_8_predecessor_in_state_13_in_data
	always @(*) begin
		if (eq_240_out) begin 
			bb_8_predecessor_in_state_13_in_data = state_13_last_BB_reg;
		end else begin
			bb_8_predecessor_in_state_13_in_data = 0;
		end
	end
	// controller for bb_9_active_in_state_8.bb_9_active_in_state_8_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_9_active_in_state_8_in_data = orOp_171_out;
		end else begin
			bb_9_active_in_state_8_in_data = 0;
		end
	end
	// controller for bb_9_predecessor_in_state_8.bb_9_predecessor_in_state_8_in_data
	always @(*) begin
		if (andOp_223_out) begin 
			bb_9_predecessor_in_state_8_in_data = 32'd1;
		end else if (eq_221_out) begin 
			bb_9_predecessor_in_state_8_in_data = state_8_last_BB_reg;
		end else begin
			bb_9_predecessor_in_state_8_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_68_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_69_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_8.br_10_happened_in_state_8_in_data
	always @(*) begin
		if (andOp_118_out) begin 
			br_10_happened_in_state_8_in_data = 1'd1;
		end else if (notOp_119_out) begin 
			br_10_happened_in_state_8_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_8_in_data = 0;
		end
	end
	// controller for br_11_happened_in_state_10.br_11_happened_in_state_10_in_data
	always @(*) begin
		if (andOp_125_out) begin 
			br_11_happened_in_state_10_in_data = 1'd1;
		end else if (notOp_126_out) begin 
			br_11_happened_in_state_10_in_data = 1'd0;
		end else begin
			br_11_happened_in_state_10_in_data = 0;
		end
	end
	// controller for br_11_happened_in_state_9.br_11_happened_in_state_9_in_data
	always @(*) begin
		if (andOp_123_out) begin 
			br_11_happened_in_state_9_in_data = 1'd1;
		end else if (notOp_124_out) begin 
			br_11_happened_in_state_9_in_data = 1'd0;
		end else begin
			br_11_happened_in_state_9_in_data = 0;
		end
	end
	// controller for br_12_happened_in_state_11.br_12_happened_in_state_11_in_data
	always @(*) begin
		if (andOp_127_out) begin 
			br_12_happened_in_state_11_in_data = 1'd1;
		end else if (notOp_128_out) begin 
			br_12_happened_in_state_11_in_data = 1'd0;
		end else begin
			br_12_happened_in_state_11_in_data = 0;
		end
	end
	// controller for br_13_happened_in_state_11.br_13_happened_in_state_11_in_data
	always @(*) begin
		if (andOp_129_out) begin 
			br_13_happened_in_state_11_in_data = 1'd1;
		end else if (notOp_130_out) begin 
			br_13_happened_in_state_11_in_data = 1'd0;
		end else begin
			br_13_happened_in_state_11_in_data = 0;
		end
	end
	// controller for br_14_happened_in_state_12.br_14_happened_in_state_12_in_data
	always @(*) begin
		if (andOp_141_out) begin 
			br_14_happened_in_state_12_in_data = 1'd1;
		end else if (notOp_142_out) begin 
			br_14_happened_in_state_12_in_data = 1'd0;
		end else begin
			br_14_happened_in_state_12_in_data = 0;
		end
	end
	// controller for br_15_happened_in_state_1.br_15_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_75_out) begin 
			br_15_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_76_out) begin 
			br_15_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_15_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_16_happened_in_state_1.br_16_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_70_out) begin 
			br_16_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_71_out) begin 
			br_16_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_16_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_17_happened_in_state_2.br_17_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_79_out) begin 
			br_17_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_80_out) begin 
			br_17_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_17_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_17_happened_in_state_3.br_17_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_83_out) begin 
			br_17_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_84_out) begin 
			br_17_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_17_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_18_happened_in_state_3.br_18_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_81_out) begin 
			br_18_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_82_out) begin 
			br_18_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_18_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_19_happened_in_state_3.br_19_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_87_out) begin 
			br_19_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_88_out) begin 
			br_19_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_19_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_1_happened_in_state_8.br_1_happened_in_state_8_in_data
	always @(*) begin
		if (andOp_114_out) begin 
			br_1_happened_in_state_8_in_data = 1'd1;
		end else if (notOp_115_out) begin 
			br_1_happened_in_state_8_in_data = 1'd0;
		end else begin
			br_1_happened_in_state_8_in_data = 0;
		end
	end
	// controller for br_20_happened_in_state_4.br_20_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_92_out) begin 
			br_20_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_93_out) begin 
			br_20_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_20_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_20_happened_in_state_5.br_20_happened_in_state_5_in_data
	always @(*) begin
		if (andOp_94_out) begin 
			br_20_happened_in_state_5_in_data = 1'd1;
		end else if (notOp_95_out) begin 
			br_20_happened_in_state_5_in_data = 1'd0;
		end else begin
			br_20_happened_in_state_5_in_data = 0;
		end
	end
	// controller for br_20_happened_in_state_6.br_20_happened_in_state_6_in_data
	always @(*) begin
		if (andOp_100_out) begin 
			br_20_happened_in_state_6_in_data = 1'd1;
		end else if (notOp_101_out) begin 
			br_20_happened_in_state_6_in_data = 1'd0;
		end else begin
			br_20_happened_in_state_6_in_data = 0;
		end
	end
	// controller for br_21_happened_in_state_6.br_21_happened_in_state_6_in_data
	always @(*) begin
		if (andOp_96_out) begin 
			br_21_happened_in_state_6_in_data = 1'd1;
		end else if (notOp_97_out) begin 
			br_21_happened_in_state_6_in_data = 1'd0;
		end else begin
			br_21_happened_in_state_6_in_data = 0;
		end
	end
	// controller for br_22_happened_in_state_6.br_22_happened_in_state_6_in_data
	always @(*) begin
		if (andOp_102_out) begin 
			br_22_happened_in_state_6_in_data = 1'd1;
		end else if (notOp_103_out) begin 
			br_22_happened_in_state_6_in_data = 1'd0;
		end else begin
			br_22_happened_in_state_6_in_data = 0;
		end
	end
	// controller for br_23_happened_in_state_7.br_23_happened_in_state_7_in_data
	always @(*) begin
		if (andOp_112_out) begin 
			br_23_happened_in_state_7_in_data = 1'd1;
		end else if (notOp_113_out) begin 
			br_23_happened_in_state_7_in_data = 1'd0;
		end else begin
			br_23_happened_in_state_7_in_data = 0;
		end
	end
	// controller for br_2_happened_in_state_11.br_2_happened_in_state_11_in_data
	always @(*) begin
		if (andOp_134_out) begin 
			br_2_happened_in_state_11_in_data = 1'd1;
		end else if (notOp_135_out) begin 
			br_2_happened_in_state_11_in_data = 1'd0;
		end else begin
			br_2_happened_in_state_11_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_12.br_3_happened_in_state_12_in_data
	always @(*) begin
		if (andOp_136_out) begin 
			br_3_happened_in_state_12_in_data = 1'd1;
		end else if (notOp_137_out) begin 
			br_3_happened_in_state_12_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_12_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_1.br_4_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_77_out) begin 
			br_4_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_78_out) begin 
			br_4_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_5_happened_in_state_3.br_5_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_85_out) begin 
			br_5_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_86_out) begin 
			br_5_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_5_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_6_happened_in_state_6.br_6_happened_in_state_6_in_data
	always @(*) begin
		if (andOp_98_out) begin 
			br_6_happened_in_state_6_in_data = 1'd1;
		end else if (notOp_99_out) begin 
			br_6_happened_in_state_6_in_data = 1'd0;
		end else begin
			br_6_happened_in_state_6_in_data = 0;
		end
	end
	// controller for br_7_happened_in_state_7.br_7_happened_in_state_7_in_data
	always @(*) begin
		if (andOp_107_out) begin 
			br_7_happened_in_state_7_in_data = 1'd1;
		end else if (notOp_108_out) begin 
			br_7_happened_in_state_7_in_data = 1'd0;
		end else begin
			br_7_happened_in_state_7_in_data = 0;
		end
	end
	// controller for br_9_happened_in_state_8.br_9_happened_in_state_8_in_data
	always @(*) begin
		if (andOp_116_out) begin 
			br_9_happened_in_state_8_in_data = 1'd1;
		end else if (notOp_117_out) begin 
			br_9_happened_in_state_8_in_data = 1'd0;
		end else begin
			br_9_happened_in_state_8_in_data = 0;
		end
	end
	// controller for concat_252.concat_252_in0
	// controller for concat_252.concat_252_in1
	// Insensitive connections
	assign concat_252_in0 = data_in_1_5_out_data;
	assign concat_252_in1 = 32'd0;
	// controller for concat_253.concat_253_in0
	// controller for concat_253.concat_253_in1
	// Insensitive connections
	assign concat_253_in0 = 32'd7;
	assign concat_253_in1 = 32'd0;
	// controller for concat_261.concat_261_in0
	// controller for concat_261.concat_261_in1
	// Insensitive connections
	assign concat_261_in0 = data_in_8_46_out_data;
	assign concat_261_in1 = 32'd0;
	// controller for concat_262.concat_262_in0
	// controller for concat_262.concat_262_in1
	// Insensitive connections
	assign concat_262_in0 = 32'd3;
	assign concat_262_in1 = 32'd7;
	// controller for data_in_10_55.data_in_10_55_in_data
	always @(*) begin
		if (eq_346_out) begin 
			data_in_10_55_in_data = data_store_9_49;
		end else if (eq_347_out) begin 
			data_in_10_55_in_data = data_store_10_54;
		end else begin
			data_in_10_55_in_data = 0;
		end
	end
	// controller for data_in_10_57.data_in_10_57_in_data
	always @(*) begin
		if (eq_346_out) begin 
			data_in_10_57_in_data = data_store_9_51;
		end else if (eq_347_out) begin 
			data_in_10_57_in_data = data_store_10_56;
		end else begin
			data_in_10_57_in_data = 0;
		end
	end
	// controller for data_in_11_59.data_in_11_59_in_data
	always @(*) begin
		if (eq_349_out) begin 
			data_in_11_59_in_data = data_store_10_53;
		end else if (eq_350_out) begin 
			data_in_11_59_in_data = data_store_11_58;
		end else begin
			data_in_11_59_in_data = 0;
		end
	end
	// controller for data_in_11_61.data_in_11_61_in_data
	always @(*) begin
		if (eq_349_out) begin 
			data_in_11_61_in_data = data_store_10_54;
		end else if (eq_350_out) begin 
			data_in_11_61_in_data = data_store_11_60;
		end else begin
			data_in_11_61_in_data = 0;
		end
	end
	// controller for data_in_11_63.data_in_11_63_in_data
	always @(*) begin
		if (eq_349_out) begin 
			data_in_11_63_in_data = data_store_10_56;
		end else if (eq_350_out) begin 
			data_in_11_63_in_data = data_store_11_62;
		end else begin
			data_in_11_63_in_data = 0;
		end
	end
	// controller for data_in_12_65.data_in_12_65_in_data
	always @(*) begin
		if (eq_352_out) begin 
			data_in_12_65_in_data = data_store_11_60;
		end else if (eq_353_out) begin 
			data_in_12_65_in_data = data_store_12_64;
		end else begin
			data_in_12_65_in_data = 0;
		end
	end
	// controller for data_in_12_67.data_in_12_67_in_data
	always @(*) begin
		if (eq_352_out) begin 
			data_in_12_67_in_data = data_store_11_62;
		end else if (eq_353_out) begin 
			data_in_12_67_in_data = data_store_12_66;
		end else begin
			data_in_12_67_in_data = 0;
		end
	end
	// controller for data_in_1_1.data_in_1_1_in_data
	always @(*) begin
		if (eq_321_out) begin 
			data_in_1_1_in_data = 32'd0;
		end else if (eq_322_out) begin 
			data_in_1_1_in_data = data_store_1_0;
		end else if (eq_323_out) begin 
			data_in_1_1_in_data = data_store_7_39;
		end else begin
			data_in_1_1_in_data = 0;
		end
	end
	// controller for data_in_1_3.data_in_1_3_in_data
	always @(*) begin
		if (eq_321_out) begin 
			data_in_1_3_in_data = 32'd0;
		end else if (eq_322_out) begin 
			data_in_1_3_in_data = data_store_1_2;
		end else if (eq_323_out) begin 
			data_in_1_3_in_data = data_store_7_41;
		end else begin
			data_in_1_3_in_data = 0;
		end
	end
	// controller for data_in_1_5.data_in_1_5_in_data
	always @(*) begin
		if (eq_321_out) begin 
			data_in_1_5_in_data = 32'd0;
		end else if (eq_322_out) begin 
			data_in_1_5_in_data = data_store_1_4;
		end else if (eq_323_out) begin 
			data_in_1_5_in_data = data_store_7_43;
		end else begin
			data_in_1_5_in_data = 0;
		end
	end
	// controller for data_in_2_11.data_in_2_11_in_data
	always @(*) begin
		if (eq_325_out) begin 
			data_in_2_11_in_data = data_store_1_4;
		end else if (eq_326_out) begin 
			data_in_2_11_in_data = data_store_2_10;
		end else begin
			data_in_2_11_in_data = 0;
		end
	end
	// controller for data_in_2_7.data_in_2_7_in_data
	always @(*) begin
		if (eq_325_out) begin 
			data_in_2_7_in_data = data_store_1_0;
		end else if (eq_326_out) begin 
			data_in_2_7_in_data = data_store_2_6;
		end else begin
			data_in_2_7_in_data = 0;
		end
	end
	// controller for data_in_2_9.data_in_2_9_in_data
	always @(*) begin
		if (eq_325_out) begin 
			data_in_2_9_in_data = data_store_1_2;
		end else if (eq_326_out) begin 
			data_in_2_9_in_data = data_store_2_8;
		end else begin
			data_in_2_9_in_data = 0;
		end
	end
	// controller for data_in_3_13.data_in_3_13_in_data
	always @(*) begin
		if (eq_327_out) begin 
			data_in_3_13_in_data = data_store_2_6;
		end else if (eq_328_out) begin 
			data_in_3_13_in_data = data_store_3_12;
		end else begin
			data_in_3_13_in_data = 0;
		end
	end
	// controller for data_in_3_15.data_in_3_15_in_data
	always @(*) begin
		if (eq_327_out) begin 
			data_in_3_15_in_data = data_store_2_8;
		end else if (eq_328_out) begin 
			data_in_3_15_in_data = data_store_3_14;
		end else begin
			data_in_3_15_in_data = 0;
		end
	end
	// controller for data_in_3_17.data_in_3_17_in_data
	always @(*) begin
		if (eq_327_out) begin 
			data_in_3_17_in_data = data_store_2_10;
		end else if (eq_328_out) begin 
			data_in_3_17_in_data = data_store_3_16;
		end else begin
			data_in_3_17_in_data = 0;
		end
	end
	// controller for data_in_4_19.data_in_4_19_in_data
	always @(*) begin
		if (eq_330_out) begin 
			data_in_4_19_in_data = data_store_3_12;
		end else if (eq_331_out) begin 
			data_in_4_19_in_data = data_store_4_18;
		end else begin
			data_in_4_19_in_data = 0;
		end
	end
	// controller for data_in_4_21.data_in_4_21_in_data
	always @(*) begin
		if (eq_330_out) begin 
			data_in_4_21_in_data = data_store_3_14;
		end else if (eq_331_out) begin 
			data_in_4_21_in_data = data_store_4_20;
		end else begin
			data_in_4_21_in_data = 0;
		end
	end
	// controller for data_in_4_23.data_in_4_23_in_data
	always @(*) begin
		if (eq_330_out) begin 
			data_in_4_23_in_data = data_store_3_16;
		end else if (eq_331_out) begin 
			data_in_4_23_in_data = data_store_4_22;
		end else begin
			data_in_4_23_in_data = 0;
		end
	end
	// controller for data_in_5_26.data_in_5_26_in_data
	always @(*) begin
		if (eq_332_out) begin 
			data_in_5_26_in_data = data_store_4_18;
		end else if (eq_333_out) begin 
			data_in_5_26_in_data = data_store_5_25;
		end else begin
			data_in_5_26_in_data = 0;
		end
	end
	// controller for data_in_5_28.data_in_5_28_in_data
	always @(*) begin
		if (eq_332_out) begin 
			data_in_5_28_in_data = data_store_4_20;
		end else if (eq_333_out) begin 
			data_in_5_28_in_data = data_store_5_27;
		end else begin
			data_in_5_28_in_data = 0;
		end
	end
	// controller for data_in_5_30.data_in_5_30_in_data
	always @(*) begin
		if (eq_332_out) begin 
			data_in_5_30_in_data = data_store_4_22;
		end else if (eq_333_out) begin 
			data_in_5_30_in_data = data_store_5_29;
		end else begin
			data_in_5_30_in_data = 0;
		end
	end
	// controller for data_in_6_32.data_in_6_32_in_data
	always @(*) begin
		if (eq_335_out) begin 
			data_in_6_32_in_data = data_store_5_24;
		end else if (eq_336_out) begin 
			data_in_6_32_in_data = data_store_6_31;
		end else begin
			data_in_6_32_in_data = 0;
		end
	end
	// controller for data_in_6_34.data_in_6_34_in_data
	always @(*) begin
		if (eq_335_out) begin 
			data_in_6_34_in_data = data_store_5_25;
		end else if (eq_336_out) begin 
			data_in_6_34_in_data = data_store_6_33;
		end else begin
			data_in_6_34_in_data = 0;
		end
	end
	// controller for data_in_6_36.data_in_6_36_in_data
	always @(*) begin
		if (eq_335_out) begin 
			data_in_6_36_in_data = data_store_5_27;
		end else if (eq_336_out) begin 
			data_in_6_36_in_data = data_store_6_35;
		end else begin
			data_in_6_36_in_data = 0;
		end
	end
	// controller for data_in_6_38.data_in_6_38_in_data
	always @(*) begin
		if (eq_335_out) begin 
			data_in_6_38_in_data = data_store_5_29;
		end else if (eq_336_out) begin 
			data_in_6_38_in_data = data_store_6_37;
		end else begin
			data_in_6_38_in_data = 0;
		end
	end
	// controller for data_in_7_40.data_in_7_40_in_data
	always @(*) begin
		if (eq_338_out) begin 
			data_in_7_40_in_data = data_store_6_33;
		end else if (eq_339_out) begin 
			data_in_7_40_in_data = data_store_7_39;
		end else begin
			data_in_7_40_in_data = 0;
		end
	end
	// controller for data_in_7_42.data_in_7_42_in_data
	always @(*) begin
		if (eq_338_out) begin 
			data_in_7_42_in_data = data_store_6_35;
		end else if (eq_339_out) begin 
			data_in_7_42_in_data = data_store_7_41;
		end else begin
			data_in_7_42_in_data = 0;
		end
	end
	// controller for data_in_7_44.data_in_7_44_in_data
	always @(*) begin
		if (eq_338_out) begin 
			data_in_7_44_in_data = data_store_6_37;
		end else if (eq_339_out) begin 
			data_in_7_44_in_data = data_store_7_43;
		end else begin
			data_in_7_44_in_data = 0;
		end
	end
	// controller for data_in_8_46.data_in_8_46_in_data
	always @(*) begin
		if (eq_340_out) begin 
			data_in_8_46_in_data = 32'd0;
		end else if (eq_341_out) begin 
			data_in_8_46_in_data = data_store_8_45;
		end else if (eq_342_out) begin 
			data_in_8_46_in_data = data_store_12_64;
		end else begin
			data_in_8_46_in_data = 0;
		end
	end
	// controller for data_in_8_48.data_in_8_48_in_data
	always @(*) begin
		if (eq_340_out) begin 
			data_in_8_48_in_data = 32'd0;
		end else if (eq_341_out) begin 
			data_in_8_48_in_data = data_store_8_47;
		end else if (eq_342_out) begin 
			data_in_8_48_in_data = data_store_12_66;
		end else begin
			data_in_8_48_in_data = 0;
		end
	end
	// controller for data_in_9_50.data_in_9_50_in_data
	always @(*) begin
		if (eq_344_out) begin 
			data_in_9_50_in_data = data_store_8_45;
		end else if (eq_345_out) begin 
			data_in_9_50_in_data = data_store_9_49;
		end else begin
			data_in_9_50_in_data = 0;
		end
	end
	// controller for data_in_9_52.data_in_9_52_in_data
	always @(*) begin
		if (eq_344_out) begin 
			data_in_9_52_in_data = data_store_8_47;
		end else if (eq_345_out) begin 
			data_in_9_52_in_data = data_store_9_51;
		end else begin
			data_in_9_52_in_data = 0;
		end
	end
	// controller for eq_143.eq_143_in0
	// controller for eq_143.eq_143_in1
	// Insensitive connections
	assign eq_143_in0 = 32'd0;
	assign eq_143_in1 = state_0_entry_BB_reg;
	// controller for eq_144.eq_144_in0
	// controller for eq_144.eq_144_in1
	// Insensitive connections
	assign eq_144_in0 = 32'd16;
	assign eq_144_in1 = state_1_entry_BB_reg;
	// controller for eq_146.eq_146_in0
	// controller for eq_146.eq_146_in1
	// Insensitive connections
	assign eq_146_in0 = 32'd15;
	assign eq_146_in1 = state_1_entry_BB_reg;
	// controller for eq_148.eq_148_in0
	// controller for eq_148.eq_148_in1
	// Insensitive connections
	assign eq_148_in0 = 32'd4;
	assign eq_148_in1 = state_1_entry_BB_reg;
	// controller for eq_149.eq_149_in0
	// controller for eq_149.eq_149_in1
	// Insensitive connections
	assign eq_149_in0 = 32'd17;
	assign eq_149_in1 = state_2_entry_BB_reg;
	// controller for eq_150.eq_150_in0
	// controller for eq_150.eq_150_in1
	// Insensitive connections
	assign eq_150_in0 = 32'd18;
	assign eq_150_in1 = state_3_entry_BB_reg;
	// controller for eq_152.eq_152_in0
	// controller for eq_152.eq_152_in1
	// Insensitive connections
	assign eq_152_in0 = 32'd17;
	assign eq_152_in1 = state_3_entry_BB_reg;
	// controller for eq_153.eq_153_in0
	// controller for eq_153.eq_153_in1
	// Insensitive connections
	assign eq_153_in0 = 32'd5;
	assign eq_153_in1 = state_3_entry_BB_reg;
	// controller for eq_155.eq_155_in0
	// controller for eq_155.eq_155_in1
	// Insensitive connections
	assign eq_155_in0 = 32'd19;
	assign eq_155_in1 = state_3_entry_BB_reg;
	// controller for eq_157.eq_157_in0
	// controller for eq_157.eq_157_in1
	// Insensitive connections
	assign eq_157_in0 = 32'd20;
	assign eq_157_in1 = state_4_entry_BB_reg;
	// controller for eq_158.eq_158_in0
	// controller for eq_158.eq_158_in1
	// Insensitive connections
	assign eq_158_in0 = 32'd20;
	assign eq_158_in1 = state_5_entry_BB_reg;
	// controller for eq_159.eq_159_in0
	// controller for eq_159.eq_159_in1
	// Insensitive connections
	assign eq_159_in0 = 32'd21;
	assign eq_159_in1 = state_6_entry_BB_reg;
	// controller for eq_161.eq_161_in0
	// controller for eq_161.eq_161_in1
	// Insensitive connections
	assign eq_161_in0 = 32'd6;
	assign eq_161_in1 = state_6_entry_BB_reg;
	// controller for eq_163.eq_163_in0
	// controller for eq_163.eq_163_in1
	// Insensitive connections
	assign eq_163_in0 = 32'd20;
	assign eq_163_in1 = state_6_entry_BB_reg;
	// controller for eq_164.eq_164_in0
	// controller for eq_164.eq_164_in1
	// Insensitive connections
	assign eq_164_in0 = 32'd22;
	assign eq_164_in1 = state_6_entry_BB_reg;
	// controller for eq_166.eq_166_in0
	// controller for eq_166.eq_166_in1
	// Insensitive connections
	assign eq_166_in0 = 32'd7;
	assign eq_166_in1 = state_7_entry_BB_reg;
	// controller for eq_168.eq_168_in0
	// controller for eq_168.eq_168_in1
	// Insensitive connections
	assign eq_168_in0 = 32'd23;
	assign eq_168_in1 = state_7_entry_BB_reg;
	// controller for eq_169.eq_169_in0
	// controller for eq_169.eq_169_in1
	// Insensitive connections
	assign eq_169_in0 = 32'd1;
	assign eq_169_in1 = state_8_entry_BB_reg;
	// controller for eq_170.eq_170_in0
	// controller for eq_170.eq_170_in1
	// Insensitive connections
	assign eq_170_in0 = 32'd9;
	assign eq_170_in1 = state_8_entry_BB_reg;
	// controller for eq_172.eq_172_in0
	// controller for eq_172.eq_172_in1
	// Insensitive connections
	assign eq_172_in0 = 32'd10;
	assign eq_172_in1 = state_8_entry_BB_reg;
	// controller for eq_174.eq_174_in0
	// controller for eq_174.eq_174_in1
	// Insensitive connections
	assign eq_174_in0 = 32'd11;
	assign eq_174_in1 = state_9_entry_BB_reg;
	// controller for eq_175.eq_175_in0
	// controller for eq_175.eq_175_in1
	// Insensitive connections
	assign eq_175_in0 = 32'd11;
	assign eq_175_in1 = state_10_entry_BB_reg;
	// controller for eq_176.eq_176_in0
	// controller for eq_176.eq_176_in1
	// Insensitive connections
	assign eq_176_in0 = 32'd12;
	assign eq_176_in1 = state_11_entry_BB_reg;
	// controller for eq_178.eq_178_in0
	// controller for eq_178.eq_178_in1
	// Insensitive connections
	assign eq_178_in0 = 32'd13;
	assign eq_178_in1 = state_11_entry_BB_reg;
	// controller for eq_180.eq_180_in0
	// controller for eq_180.eq_180_in1
	// Insensitive connections
	assign eq_180_in0 = 32'd2;
	assign eq_180_in1 = state_11_entry_BB_reg;
	// controller for eq_181.eq_181_in0
	// controller for eq_181.eq_181_in1
	// Insensitive connections
	assign eq_181_in0 = 32'd3;
	assign eq_181_in1 = state_12_entry_BB_reg;
	// controller for eq_183.eq_183_in0
	// controller for eq_183.eq_183_in1
	// Insensitive connections
	assign eq_183_in0 = 32'd14;
	assign eq_183_in1 = state_12_entry_BB_reg;
	// controller for eq_184.eq_184_in0
	// controller for eq_184.eq_184_in1
	// Insensitive connections
	assign eq_184_in0 = 32'd8;
	assign eq_184_in1 = state_13_entry_BB_reg;
	// controller for eq_185.eq_185_in0
	// controller for eq_185.eq_185_in1
	// Insensitive connections
	assign eq_185_in0 = 32'd0;
	assign eq_185_in1 = state_0_entry_BB_reg;
	// controller for eq_186.eq_186_in0
	// controller for eq_186.eq_186_in1
	// Insensitive connections
	assign eq_186_in0 = 32'd16;
	assign eq_186_in1 = state_1_entry_BB_reg;
	// controller for eq_189.eq_189_in0
	// controller for eq_189.eq_189_in1
	// Insensitive connections
	assign eq_189_in0 = 32'd15;
	assign eq_189_in1 = state_1_entry_BB_reg;
	// controller for eq_192.eq_192_in0
	// controller for eq_192.eq_192_in1
	// Insensitive connections
	assign eq_192_in0 = 32'd4;
	assign eq_192_in1 = state_1_entry_BB_reg;
	// controller for eq_193.eq_193_in0
	// controller for eq_193.eq_193_in1
	// Insensitive connections
	assign eq_193_in0 = 32'd17;
	assign eq_193_in1 = state_2_entry_BB_reg;
	// controller for eq_194.eq_194_in0
	// controller for eq_194.eq_194_in1
	// Insensitive connections
	assign eq_194_in0 = 32'd18;
	assign eq_194_in1 = state_3_entry_BB_reg;
	// controller for eq_197.eq_197_in0
	// controller for eq_197.eq_197_in1
	// Insensitive connections
	assign eq_197_in0 = 32'd17;
	assign eq_197_in1 = state_3_entry_BB_reg;
	// controller for eq_198.eq_198_in0
	// controller for eq_198.eq_198_in1
	// Insensitive connections
	assign eq_198_in0 = 32'd5;
	assign eq_198_in1 = state_3_entry_BB_reg;
	// controller for eq_201.eq_201_in0
	// controller for eq_201.eq_201_in1
	// Insensitive connections
	assign eq_201_in0 = 32'd19;
	assign eq_201_in1 = state_3_entry_BB_reg;
	// controller for eq_204.eq_204_in0
	// controller for eq_204.eq_204_in1
	// Insensitive connections
	assign eq_204_in0 = 32'd20;
	assign eq_204_in1 = state_4_entry_BB_reg;
	// controller for eq_205.eq_205_in0
	// controller for eq_205.eq_205_in1
	// Insensitive connections
	assign eq_205_in0 = 32'd20;
	assign eq_205_in1 = state_5_entry_BB_reg;
	// controller for eq_206.eq_206_in0
	// controller for eq_206.eq_206_in1
	// Insensitive connections
	assign eq_206_in0 = 32'd21;
	assign eq_206_in1 = state_6_entry_BB_reg;
	// controller for eq_209.eq_209_in0
	// controller for eq_209.eq_209_in1
	// Insensitive connections
	assign eq_209_in0 = 32'd6;
	assign eq_209_in1 = state_6_entry_BB_reg;
	// controller for eq_212.eq_212_in0
	// controller for eq_212.eq_212_in1
	// Insensitive connections
	assign eq_212_in0 = 32'd20;
	assign eq_212_in1 = state_6_entry_BB_reg;
	// controller for eq_213.eq_213_in0
	// controller for eq_213.eq_213_in1
	// Insensitive connections
	assign eq_213_in0 = 32'd22;
	assign eq_213_in1 = state_6_entry_BB_reg;
	// controller for eq_216.eq_216_in0
	// controller for eq_216.eq_216_in1
	// Insensitive connections
	assign eq_216_in0 = 32'd7;
	assign eq_216_in1 = state_7_entry_BB_reg;
	// controller for eq_219.eq_219_in0
	// controller for eq_219.eq_219_in1
	// Insensitive connections
	assign eq_219_in0 = 32'd23;
	assign eq_219_in1 = state_7_entry_BB_reg;
	// controller for eq_220.eq_220_in0
	// controller for eq_220.eq_220_in1
	// Insensitive connections
	assign eq_220_in0 = 32'd1;
	assign eq_220_in1 = state_8_entry_BB_reg;
	// controller for eq_221.eq_221_in0
	// controller for eq_221.eq_221_in1
	// Insensitive connections
	assign eq_221_in0 = 32'd9;
	assign eq_221_in1 = state_8_entry_BB_reg;
	// controller for eq_224.eq_224_in0
	// controller for eq_224.eq_224_in1
	// Insensitive connections
	assign eq_224_in0 = 32'd10;
	assign eq_224_in1 = state_8_entry_BB_reg;
	// controller for eq_227.eq_227_in0
	// controller for eq_227.eq_227_in1
	// Insensitive connections
	assign eq_227_in0 = 32'd11;
	assign eq_227_in1 = state_9_entry_BB_reg;
	// controller for eq_228.eq_228_in0
	// controller for eq_228.eq_228_in1
	// Insensitive connections
	assign eq_228_in0 = 32'd11;
	assign eq_228_in1 = state_10_entry_BB_reg;
	// controller for eq_229.eq_229_in0
	// controller for eq_229.eq_229_in1
	// Insensitive connections
	assign eq_229_in0 = 32'd12;
	assign eq_229_in1 = state_11_entry_BB_reg;
	// controller for eq_232.eq_232_in0
	// controller for eq_232.eq_232_in1
	// Insensitive connections
	assign eq_232_in0 = 32'd13;
	assign eq_232_in1 = state_11_entry_BB_reg;
	// controller for eq_235.eq_235_in0
	// controller for eq_235.eq_235_in1
	// Insensitive connections
	assign eq_235_in0 = 32'd2;
	assign eq_235_in1 = state_11_entry_BB_reg;
	// controller for eq_236.eq_236_in0
	// controller for eq_236.eq_236_in1
	// Insensitive connections
	assign eq_236_in0 = 32'd3;
	assign eq_236_in1 = state_12_entry_BB_reg;
	// controller for eq_239.eq_239_in0
	// controller for eq_239.eq_239_in1
	// Insensitive connections
	assign eq_239_in0 = 32'd14;
	assign eq_239_in1 = state_12_entry_BB_reg;
	// controller for eq_240.eq_240_in0
	// controller for eq_240.eq_240_in1
	// Insensitive connections
	assign eq_240_in0 = 32'd8;
	assign eq_240_in1 = state_13_entry_BB_reg;
	// controller for eq_320.eq_320_in0
	// controller for eq_320.eq_320_in1
	// Insensitive connections
	assign eq_320_in0 = 32'd0;
	assign eq_320_in1 = state_0_last_state;
	// controller for eq_321.eq_321_in0
	// controller for eq_321.eq_321_in1
	// Insensitive connections
	assign eq_321_in0 = 32'd0;
	assign eq_321_in1 = state_1_last_state;
	// controller for eq_322.eq_322_in0
	// controller for eq_322.eq_322_in1
	// Insensitive connections
	assign eq_322_in0 = 32'd1;
	assign eq_322_in1 = state_1_last_state;
	// controller for eq_323.eq_323_in0
	// controller for eq_323.eq_323_in1
	// Insensitive connections
	assign eq_323_in0 = 32'd7;
	assign eq_323_in1 = state_1_last_state;
	// controller for eq_325.eq_325_in0
	// controller for eq_325.eq_325_in1
	// Insensitive connections
	assign eq_325_in0 = 32'd1;
	assign eq_325_in1 = state_2_last_state;
	// controller for eq_326.eq_326_in0
	// controller for eq_326.eq_326_in1
	// Insensitive connections
	assign eq_326_in0 = 32'd2;
	assign eq_326_in1 = state_2_last_state;
	// controller for eq_327.eq_327_in0
	// controller for eq_327.eq_327_in1
	// Insensitive connections
	assign eq_327_in0 = 32'd2;
	assign eq_327_in1 = state_3_last_state;
	// controller for eq_328.eq_328_in0
	// controller for eq_328.eq_328_in1
	// Insensitive connections
	assign eq_328_in0 = 32'd3;
	assign eq_328_in1 = state_3_last_state;
	// controller for eq_330.eq_330_in0
	// controller for eq_330.eq_330_in1
	// Insensitive connections
	assign eq_330_in0 = 32'd3;
	assign eq_330_in1 = state_4_last_state;
	// controller for eq_331.eq_331_in0
	// controller for eq_331.eq_331_in1
	// Insensitive connections
	assign eq_331_in0 = 32'd4;
	assign eq_331_in1 = state_4_last_state;
	// controller for eq_332.eq_332_in0
	// controller for eq_332.eq_332_in1
	// Insensitive connections
	assign eq_332_in0 = 32'd4;
	assign eq_332_in1 = state_5_last_state;
	// controller for eq_333.eq_333_in0
	// controller for eq_333.eq_333_in1
	// Insensitive connections
	assign eq_333_in0 = 32'd5;
	assign eq_333_in1 = state_5_last_state;
	// controller for eq_335.eq_335_in0
	// controller for eq_335.eq_335_in1
	// Insensitive connections
	assign eq_335_in0 = 32'd5;
	assign eq_335_in1 = state_6_last_state;
	// controller for eq_336.eq_336_in0
	// controller for eq_336.eq_336_in1
	// Insensitive connections
	assign eq_336_in0 = 32'd6;
	assign eq_336_in1 = state_6_last_state;
	// controller for eq_338.eq_338_in0
	// controller for eq_338.eq_338_in1
	// Insensitive connections
	assign eq_338_in0 = 32'd6;
	assign eq_338_in1 = state_7_last_state;
	// controller for eq_339.eq_339_in0
	// controller for eq_339.eq_339_in1
	// Insensitive connections
	assign eq_339_in0 = 32'd7;
	assign eq_339_in1 = state_7_last_state;
	// controller for eq_340.eq_340_in0
	// controller for eq_340.eq_340_in1
	// Insensitive connections
	assign eq_340_in0 = 32'd7;
	assign eq_340_in1 = state_8_last_state;
	// controller for eq_341.eq_341_in0
	// controller for eq_341.eq_341_in1
	// Insensitive connections
	assign eq_341_in0 = 32'd8;
	assign eq_341_in1 = state_8_last_state;
	// controller for eq_342.eq_342_in0
	// controller for eq_342.eq_342_in1
	// Insensitive connections
	assign eq_342_in0 = 32'd12;
	assign eq_342_in1 = state_8_last_state;
	// controller for eq_344.eq_344_in0
	// controller for eq_344.eq_344_in1
	// Insensitive connections
	assign eq_344_in0 = 32'd8;
	assign eq_344_in1 = state_9_last_state;
	// controller for eq_345.eq_345_in0
	// controller for eq_345.eq_345_in1
	// Insensitive connections
	assign eq_345_in0 = 32'd9;
	assign eq_345_in1 = state_9_last_state;
	// controller for eq_346.eq_346_in0
	// controller for eq_346.eq_346_in1
	// Insensitive connections
	assign eq_346_in0 = 32'd9;
	assign eq_346_in1 = state_10_last_state;
	// controller for eq_347.eq_347_in0
	// controller for eq_347.eq_347_in1
	// Insensitive connections
	assign eq_347_in0 = 32'd10;
	assign eq_347_in1 = state_10_last_state;
	// controller for eq_349.eq_349_in0
	// controller for eq_349.eq_349_in1
	// Insensitive connections
	assign eq_349_in0 = 32'd10;
	assign eq_349_in1 = state_11_last_state;
	// controller for eq_350.eq_350_in0
	// controller for eq_350.eq_350_in1
	// Insensitive connections
	assign eq_350_in0 = 32'd11;
	assign eq_350_in1 = state_11_last_state;
	// controller for eq_352.eq_352_in0
	// controller for eq_352.eq_352_in1
	// Insensitive connections
	assign eq_352_in0 = 32'd11;
	assign eq_352_in1 = state_12_last_state;
	// controller for eq_353.eq_353_in0
	// controller for eq_353.eq_353_in1
	// Insensitive connections
	assign eq_353_in0 = 32'd12;
	assign eq_353_in1 = state_12_last_state;
	// controller for eq_354.eq_354_in0
	// controller for eq_354.eq_354_in1
	// Insensitive connections
	assign eq_354_in0 = 32'd12;
	assign eq_354_in1 = state_13_last_state;
	// controller for eq_355.eq_355_in0
	// controller for eq_355.eq_355_in1
	// Insensitive connections
	assign eq_355_in0 = 32'd13;
	assign eq_355_in1 = state_13_last_state;
	// controller for icmp_icmp26.icmp_icmp26_in0
	// controller for icmp_icmp26.icmp_icmp26_in1
	// Insensitive connections
	assign icmp_icmp26_in0 = data_in_7_44_out_data;
	assign icmp_icmp26_in1 = 32'd15;
	// controller for icmp_icmp45.icmp_icmp45_in0
	// controller for icmp_icmp45.icmp_icmp45_in1
	// Insensitive connections
	assign icmp_icmp45_in0 = data_in_12_65_out_data;
	assign icmp_icmp45_in1 = 32'd15;
	// controller for mul_mul41.mul_mul41_in0
	// controller for mul_mul41.mul_mul41_in1
	// Insensitive connections
	assign mul_mul41_in0 = 32'd2;
	assign mul_mul41_in1 = data_in_11_59_out_data;
	// controller for notOp_101.notOp_101_in0
	// Insensitive connections
	assign notOp_101_in0 = andOp_100_out;
	// controller for notOp_103.notOp_103_in0
	// Insensitive connections
	assign notOp_103_in0 = andOp_102_out;
	// controller for notOp_105.notOp_105_in0
	// Insensitive connections
	assign notOp_105_in0 = _____dlr_0___eq___alloca___dlr_builtin_fifo_32_write_ready;
	// controller for notOp_108.notOp_108_in0
	// Insensitive connections
	assign notOp_108_in0 = andOp_107_out;
	// controller for notOp_110.notOp_110_in0
	// Insensitive connections
	assign notOp_110_in0 = icmp_icmp26_out;
	// controller for notOp_113.notOp_113_in0
	// Insensitive connections
	assign notOp_113_in0 = andOp_112_out;
	// controller for notOp_115.notOp_115_in0
	// Insensitive connections
	assign notOp_115_in0 = andOp_114_out;
	// controller for notOp_117.notOp_117_in0
	// Insensitive connections
	assign notOp_117_in0 = andOp_116_out;
	// controller for notOp_119.notOp_119_in0
	// Insensitive connections
	assign notOp_119_in0 = andOp_118_out;
	// controller for notOp_121.notOp_121_in0
	// Insensitive connections
	assign notOp_121_in0 = _____dlr_0___eq___alloca___dlr_builtin_fifo_32_read_ready;
	// controller for notOp_124.notOp_124_in0
	// Insensitive connections
	assign notOp_124_in0 = andOp_123_out;
	// controller for notOp_126.notOp_126_in0
	// Insensitive connections
	assign notOp_126_in0 = andOp_125_out;
	// controller for notOp_128.notOp_128_in0
	// Insensitive connections
	assign notOp_128_in0 = andOp_127_out;
	// controller for notOp_130.notOp_130_in0
	// Insensitive connections
	assign notOp_130_in0 = andOp_129_out;
	// controller for notOp_132.notOp_132_in0
	// Insensitive connections
	assign notOp_132_in0 = arg_2_write_ready;
	// controller for notOp_135.notOp_135_in0
	// Insensitive connections
	assign notOp_135_in0 = andOp_134_out;
	// controller for notOp_137.notOp_137_in0
	// Insensitive connections
	assign notOp_137_in0 = andOp_136_out;
	// controller for notOp_139.notOp_139_in0
	// Insensitive connections
	assign notOp_139_in0 = icmp_icmp45_out;
	// controller for notOp_142.notOp_142_in0
	// Insensitive connections
	assign notOp_142_in0 = andOp_141_out;
	// controller for notOp_187.notOp_187_in0
	// Insensitive connections
	assign notOp_187_in0 = eq_186_out;
	// controller for notOp_190.notOp_190_in0
	// Insensitive connections
	assign notOp_190_in0 = eq_189_out;
	// controller for notOp_195.notOp_195_in0
	// Insensitive connections
	assign notOp_195_in0 = eq_194_out;
	// controller for notOp_199.notOp_199_in0
	// Insensitive connections
	assign notOp_199_in0 = eq_198_out;
	// controller for notOp_202.notOp_202_in0
	// Insensitive connections
	assign notOp_202_in0 = eq_201_out;
	// controller for notOp_207.notOp_207_in0
	// Insensitive connections
	assign notOp_207_in0 = eq_206_out;
	// controller for notOp_210.notOp_210_in0
	// Insensitive connections
	assign notOp_210_in0 = eq_209_out;
	// controller for notOp_214.notOp_214_in0
	// Insensitive connections
	assign notOp_214_in0 = eq_213_out;
	// controller for notOp_217.notOp_217_in0
	// Insensitive connections
	assign notOp_217_in0 = eq_216_out;
	// controller for notOp_222.notOp_222_in0
	// Insensitive connections
	assign notOp_222_in0 = eq_221_out;
	// controller for notOp_225.notOp_225_in0
	// Insensitive connections
	assign notOp_225_in0 = eq_224_out;
	// controller for notOp_230.notOp_230_in0
	// Insensitive connections
	assign notOp_230_in0 = eq_229_out;
	// controller for notOp_233.notOp_233_in0
	// Insensitive connections
	assign notOp_233_in0 = eq_232_out;
	// controller for notOp_237.notOp_237_in0
	// Insensitive connections
	assign notOp_237_in0 = eq_236_out;
	// controller for notOp_278.notOp_278_in0
	// Insensitive connections
	assign notOp_278_in0 = andOp_109_out;
	// controller for notOp_280.notOp_280_in0
	// Insensitive connections
	assign notOp_280_in0 = andOp_270_out;
	// controller for notOp_282.notOp_282_in0
	// Insensitive connections
	assign notOp_282_in0 = andOp_74_out;
	// controller for notOp_284.notOp_284_in0
	// Insensitive connections
	assign notOp_284_in0 = andOp_72_out;
	// controller for notOp_286.notOp_286_in0
	// Insensitive connections
	assign notOp_286_in0 = andOp_271_out;
	// controller for notOp_288.notOp_288_in0
	// Insensitive connections
	assign notOp_288_in0 = andOp_91_out;
	// controller for notOp_290.notOp_290_in0
	// Insensitive connections
	assign notOp_290_in0 = andOp_89_out;
	// controller for notOp_292.notOp_292_in0
	// Insensitive connections
	assign notOp_292_in0 = andOp_272_out;
	// controller for notOp_294.notOp_294_in0
	// Insensitive connections
	assign notOp_294_in0 = andOp_106_out;
	// controller for notOp_296.notOp_296_in0
	// Insensitive connections
	assign notOp_296_in0 = andOp_273_out;
	// controller for notOp_298.notOp_298_in0
	// Insensitive connections
	assign notOp_298_in0 = andOp_104_out;
	// controller for notOp_300.notOp_300_in0
	// Insensitive connections
	assign notOp_300_in0 = andOp_122_out;
	// controller for notOp_302.notOp_302_in0
	// Insensitive connections
	assign notOp_302_in0 = andOp_138_out;
	// controller for notOp_304.notOp_304_in0
	// Insensitive connections
	assign notOp_304_in0 = andOp_274_out;
	// controller for notOp_306.notOp_306_in0
	// Insensitive connections
	assign notOp_306_in0 = andOp_120_out;
	// controller for notOp_308.notOp_308_in0
	// Insensitive connections
	assign notOp_308_in0 = andOp_275_out;
	// controller for notOp_310.notOp_310_in0
	// Insensitive connections
	assign notOp_310_in0 = andOp_123_out;
	// controller for notOp_312.notOp_312_in0
	// Insensitive connections
	assign notOp_312_in0 = andOp_133_out;
	// controller for notOp_314.notOp_314_in0
	// Insensitive connections
	assign notOp_314_in0 = andOp_131_out;
	// controller for notOp_316.notOp_316_in0
	// Insensitive connections
	assign notOp_316_in0 = andOp_276_out;
	// controller for notOp_318.notOp_318_in0
	// Insensitive connections
	assign notOp_318_in0 = andOp_277_out;
	// controller for notOp_69.notOp_69_in0
	// Insensitive connections
	assign notOp_69_in0 = andOp_68_out;
	// controller for notOp_71.notOp_71_in0
	// Insensitive connections
	assign notOp_71_in0 = andOp_70_out;
	// controller for notOp_73.notOp_73_in0
	// Insensitive connections
	assign notOp_73_in0 = arg_0_read_ready;
	// controller for notOp_76.notOp_76_in0
	// Insensitive connections
	assign notOp_76_in0 = andOp_75_out;
	// controller for notOp_78.notOp_78_in0
	// Insensitive connections
	assign notOp_78_in0 = andOp_77_out;
	// controller for notOp_80.notOp_80_in0
	// Insensitive connections
	assign notOp_80_in0 = andOp_79_out;
	// controller for notOp_82.notOp_82_in0
	// Insensitive connections
	assign notOp_82_in0 = andOp_81_out;
	// controller for notOp_84.notOp_84_in0
	// Insensitive connections
	assign notOp_84_in0 = andOp_83_out;
	// controller for notOp_86.notOp_86_in0
	// Insensitive connections
	assign notOp_86_in0 = andOp_85_out;
	// controller for notOp_88.notOp_88_in0
	// Insensitive connections
	assign notOp_88_in0 = andOp_87_out;
	// controller for notOp_90.notOp_90_in0
	// Insensitive connections
	assign notOp_90_in0 = arg_1_read_ready;
	// controller for notOp_93.notOp_93_in0
	// Insensitive connections
	assign notOp_93_in0 = andOp_92_out;
	// controller for notOp_95.notOp_95_in0
	// Insensitive connections
	assign notOp_95_in0 = andOp_94_out;
	// controller for notOp_97.notOp_97_in0
	// Insensitive connections
	assign notOp_97_in0 = andOp_96_out;
	// controller for notOp_99.notOp_99_in0
	// Insensitive connections
	assign notOp_99_in0 = andOp_98_out;
	// controller for orOp_145.orOp_145_in0
	// controller for orOp_145.orOp_145_in1
	// Insensitive connections
	assign orOp_145_in0 = eq_144_out;
	assign orOp_145_in1 = andOp_75_out;
	// controller for orOp_147.orOp_147_in0
	// controller for orOp_147.orOp_147_in1
	// Insensitive connections
	assign orOp_147_in0 = eq_146_out;
	assign orOp_147_in1 = andOp_77_out;
	// controller for orOp_151.orOp_151_in0
	// controller for orOp_151.orOp_151_in1
	// Insensitive connections
	assign orOp_151_in0 = eq_150_out;
	assign orOp_151_in1 = andOp_85_out;
	// controller for orOp_154.orOp_154_in0
	// controller for orOp_154.orOp_154_in1
	// Insensitive connections
	assign orOp_154_in0 = eq_153_out;
	assign orOp_154_in1 = andOp_79_out;
	// controller for orOp_156.orOp_156_in0
	// controller for orOp_156.orOp_156_in1
	// Insensitive connections
	assign orOp_156_in0 = eq_155_out;
	assign orOp_156_in1 = andOp_81_out;
	// controller for orOp_160.orOp_160_in0
	// controller for orOp_160.orOp_160_in1
	// Insensitive connections
	assign orOp_160_in0 = eq_159_out;
	assign orOp_160_in1 = andOp_98_out;
	// controller for orOp_162.orOp_162_in0
	// controller for orOp_162.orOp_162_in1
	// Insensitive connections
	assign orOp_162_in0 = eq_161_out;
	assign orOp_162_in1 = andOp_92_out;
	// controller for orOp_165.orOp_165_in0
	// controller for orOp_165.orOp_165_in1
	// Insensitive connections
	assign orOp_165_in0 = eq_164_out;
	assign orOp_165_in1 = andOp_96_out;
	// controller for orOp_167.orOp_167_in0
	// controller for orOp_167.orOp_167_in1
	// Insensitive connections
	assign orOp_167_in0 = eq_166_out;
	assign orOp_167_in1 = andOp_112_out;
	// controller for orOp_171.orOp_171_in0
	// controller for orOp_171.orOp_171_in1
	// Insensitive connections
	assign orOp_171_in0 = eq_170_out;
	assign orOp_171_in1 = andOp_114_out;
	// controller for orOp_173.orOp_173_in0
	// controller for orOp_173.orOp_173_in1
	// Insensitive connections
	assign orOp_173_in0 = eq_172_out;
	assign orOp_173_in1 = andOp_116_out;
	// controller for orOp_177.orOp_177_in0
	// controller for orOp_177.orOp_177_in1
	// Insensitive connections
	assign orOp_177_in0 = eq_176_out;
	assign orOp_177_in1 = andOp_134_out;
	// controller for orOp_179.orOp_179_in0
	// controller for orOp_179.orOp_179_in1
	// Insensitive connections
	assign orOp_179_in0 = eq_178_out;
	assign orOp_179_in1 = andOp_127_out;
	// controller for orOp_182.orOp_182_in0
	// controller for orOp_182.orOp_182_in1
	// Insensitive connections
	assign orOp_182_in0 = eq_181_out;
	assign orOp_182_in1 = andOp_141_out;
	// controller for phi_phi31.phi_phi31_in
	// controller for phi_phi31.phi_phi31_last_block
	// controller for phi_phi31.phi_phi31_s
	// Insensitive connections
	assign phi_phi31_in = concat_261_out;
	assign phi_phi31_last_block = bb_1_predecessor_in_state_8_out_data;
	assign phi_phi31_s = concat_262_out;
	// controller for phi_phi6.phi_phi6_in
	// controller for phi_phi6.phi_phi6_last_block
	// controller for phi_phi6.phi_phi6_s
	// Insensitive connections
	assign phi_phi6_in = concat_252_out;
	assign phi_phi6_last_block = bb_4_predecessor_in_state_1_out_data;
	assign phi_phi6_s = concat_253_out;
	// controller for ret47.valid_reg
	always @(*) begin
		if (andOp_269_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			data_store_10_53 <= 0;
		end else begin
			if (andOp_348_out) begin
				data_store_10_53 <= _____dlr_0___eq___alloca___dlr_builtin_fifo_32_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_10_54 <= 0;
		end else begin
			if (state_10_is_active) begin
				data_store_10_54 <= data_in_10_55_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_10_56 <= 0;
		end else begin
			if (state_10_is_active) begin
				data_store_10_56 <= data_in_10_57_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_11_58 <= 0;
		end else begin
			if (state_11_is_active) begin
				data_store_11_58 <= data_in_11_59_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_11_60 <= 0;
		end else begin
			if (state_11_is_active) begin
				data_store_11_60 <= data_in_11_61_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_11_62 <= 0;
		end else begin
			if (andOp_351_out) begin
				data_store_11_62 <= mul_mul41_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_12_64 <= 0;
		end else begin
			if (state_12_is_active) begin
				data_store_12_64 <= data_in_12_65_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_12_66 <= 0;
		end else begin
			if (state_12_is_active) begin
				data_store_12_66 <= data_in_12_67_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_0 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_0 <= data_in_1_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_2 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_2 <= data_in_1_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_4 <= 0;
		end else begin
			if (andOp_324_out) begin
				data_store_1_4 <= add_add7_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_10 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_10 <= data_in_2_11_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_6 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_6 <= data_in_2_7_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_8 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_8 <= data_in_2_9_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_12 <= 0;
		end else begin
			if (andOp_329_out) begin
				data_store_3_12 <= arg_0_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_14 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_14 <= data_in_3_15_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_16 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_16 <= data_in_3_17_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_18 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_18 <= data_in_4_19_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_20 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_20 <= data_in_4_21_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_22 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_22 <= data_in_4_23_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_24 <= 0;
		end else begin
			if (andOp_334_out) begin
				data_store_5_24 <= arg_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_25 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_25 <= data_in_5_26_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_27 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_27 <= data_in_5_28_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_29 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_29 <= data_in_5_30_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_31 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_31 <= data_in_6_32_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_33 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_33 <= data_in_6_34_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_35 <= 0;
		end else begin
			if (andOp_337_out) begin
				data_store_6_35 <= add_add22_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_37 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_37 <= data_in_6_38_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_7_39 <= 0;
		end else begin
			if (state_7_is_active) begin
				data_store_7_39 <= data_in_7_40_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_7_41 <= 0;
		end else begin
			if (state_7_is_active) begin
				data_store_7_41 <= data_in_7_42_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_7_43 <= 0;
		end else begin
			if (state_7_is_active) begin
				data_store_7_43 <= data_in_7_44_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_8_45 <= 0;
		end else begin
			if (andOp_343_out) begin
				data_store_8_45 <= add_add32_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_8_47 <= 0;
		end else begin
			if (state_8_is_active) begin
				data_store_8_47 <= data_in_8_48_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_9_49 <= 0;
		end else begin
			if (state_9_is_active) begin
				data_store_9_49 <= data_in_9_50_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_9_51 <= 0;
		end else begin
			if (state_9_is_active) begin
				data_store_9_51 <= data_in_9_52_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_104_out) begin
				global_state <= 32'd7;
			end
			if (andOp_106_out) begin
				global_state <= 32'd6;
			end
			if (andOp_109_out) begin
				global_state <= 32'd1;
			end
			if (andOp_120_out) begin
				global_state <= 32'd9;
			end
			if (andOp_122_out) begin
				global_state <= 32'd8;
			end
			if (andOp_123_out) begin
				global_state <= 32'd11;
			end
			if (andOp_131_out) begin
				global_state <= 32'd12;
			end
			if (andOp_133_out) begin
				global_state <= 32'd11;
			end
			if (andOp_138_out) begin
				global_state <= 32'd8;
			end
			if (andOp_270_out) begin
				global_state <= 32'd1;
			end
			if (andOp_271_out) begin
				global_state <= 32'd3;
			end
			if (andOp_272_out) begin
				global_state <= 32'd5;
			end
			if (andOp_273_out) begin
				global_state <= 32'd6;
			end
			if (andOp_274_out) begin
				global_state <= 32'd8;
			end
			if (andOp_275_out) begin
				global_state <= 32'd10;
			end
			if (andOp_276_out) begin
				global_state <= 32'd13;
			end
			if (andOp_277_out) begin
				global_state <= 32'd13;
			end
			if (andOp_72_out) begin
				global_state <= 32'd2;
			end
			if (andOp_74_out) begin
				global_state <= 32'd1;
			end
			if (andOp_89_out) begin
				global_state <= 32'd4;
			end
			if (andOp_91_out) begin
				global_state <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (1'd1) begin
				state_0_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_10_entry_BB_reg <= 0;
		end else begin
			if (andOp_275_out) begin
				state_10_entry_BB_reg <= 32'd11;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_10_is_active <= 0;
		end else begin
			if (andOp_275_out) begin
				state_10_is_active <= 1'd1;
			end
			if (andOp_309_out) begin
				state_10_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_10_last_BB_reg <= 0;
		end else begin
			if (andOp_275_out) begin
				state_10_last_BB_reg <= bb_11_predecessor_in_state_9_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_10_last_state <= 0;
		end else begin
			if (andOp_275_out) begin
				state_10_last_state <= 32'd9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_11_entry_BB_reg <= 0;
		end else begin
			if (andOp_123_out) begin
				state_11_entry_BB_reg <= 32'd2;
			end
			if (andOp_133_out) begin
				state_11_entry_BB_reg <= 32'd13;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_11_is_active <= 0;
		end else begin
			if (andOp_123_out) begin
				state_11_is_active <= 1'd1;
			end
			if (andOp_133_out) begin
				state_11_is_active <= 1'd1;
			end
			if (andOp_313_out) begin
				state_11_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_11_last_BB_reg <= 0;
		end else begin
			if (andOp_123_out) begin
				state_11_last_BB_reg <= 32'd11;
			end
			if (andOp_133_out) begin
				state_11_last_BB_reg <= 32'd13;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_11_last_state <= 0;
		end else begin
			if (andOp_123_out) begin
				state_11_last_state <= 32'd10;
			end
			if (andOp_133_out) begin
				state_11_last_state <= 32'd11;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_12_entry_BB_reg <= 0;
		end else begin
			if (andOp_131_out) begin
				state_12_entry_BB_reg <= 32'd14;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_12_is_active <= 0;
		end else begin
			if (andOp_131_out) begin
				state_12_is_active <= 1'd1;
			end
			if (andOp_315_out) begin
				state_12_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_12_last_BB_reg <= 0;
		end else begin
			if (andOp_131_out) begin
				state_12_last_BB_reg <= 32'd13;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_12_last_state <= 0;
		end else begin
			if (andOp_131_out) begin
				state_12_last_state <= 32'd11;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_13_entry_BB_reg <= 0;
		end else begin
			if (andOp_276_out) begin
				state_13_entry_BB_reg <= 32'd8;
			end
			if (andOp_277_out) begin
				state_13_entry_BB_reg <= 32'd8;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_13_is_active <= 1;
		end else begin
			if (andOp_276_out) begin
				state_13_is_active <= 1'd1;
			end
			if (andOp_277_out) begin
				state_13_is_active <= 1'd1;
			end
			if (andOp_319_out) begin
				state_13_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_13_last_BB_reg <= 0;
		end else begin
			if (andOp_276_out) begin
				state_13_last_BB_reg <= 32'd3;
			end
			if (andOp_277_out) begin
				state_13_last_BB_reg <= bb_8_predecessor_in_state_13_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_13_last_state <= 0;
		end else begin
			if (andOp_276_out) begin
				state_13_last_state <= 32'd12;
			end
			if (andOp_277_out) begin
				state_13_last_state <= 32'd13;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_109_out) begin
				state_1_entry_BB_reg <= 32'd4;
			end
			if (andOp_270_out) begin
				state_1_entry_BB_reg <= 32'd4;
			end
			if (andOp_74_out) begin
				state_1_entry_BB_reg <= 32'd16;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 1;
		end else begin
			if (andOp_109_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_270_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_283_out) begin
				state_1_is_active <= 1'd0;
			end
			if (andOp_74_out) begin
				state_1_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_109_out) begin
				state_1_last_BB_reg <= 32'd7;
			end
			if (andOp_270_out) begin
				state_1_last_BB_reg <= 32'd0;
			end
			if (andOp_74_out) begin
				state_1_last_BB_reg <= 32'd16;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_109_out) begin
				state_1_last_state <= 32'd7;
			end
			if (andOp_270_out) begin
				state_1_last_state <= 32'd0;
			end
			if (andOp_74_out) begin
				state_1_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_72_out) begin
				state_2_entry_BB_reg <= 32'd17;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_285_out) begin
				state_2_is_active <= 1'd0;
			end
			if (andOp_72_out) begin
				state_2_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_72_out) begin
				state_2_last_BB_reg <= 32'd16;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_72_out) begin
				state_2_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_271_out) begin
				state_3_entry_BB_reg <= 32'd17;
			end
			if (andOp_91_out) begin
				state_3_entry_BB_reg <= 32'd19;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_271_out) begin
				state_3_is_active <= 1'd1;
			end
			if (andOp_289_out) begin
				state_3_is_active <= 1'd0;
			end
			if (andOp_91_out) begin
				state_3_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_271_out) begin
				state_3_last_BB_reg <= bb_17_predecessor_in_state_2_out_data;
			end
			if (andOp_91_out) begin
				state_3_last_BB_reg <= 32'd19;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_state <= 0;
		end else begin
			if (andOp_271_out) begin
				state_3_last_state <= 32'd2;
			end
			if (andOp_91_out) begin
				state_3_last_state <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_89_out) begin
				state_4_entry_BB_reg <= 32'd20;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_291_out) begin
				state_4_is_active <= 1'd0;
			end
			if (andOp_89_out) begin
				state_4_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_89_out) begin
				state_4_last_BB_reg <= 32'd19;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_state <= 0;
		end else begin
			if (andOp_89_out) begin
				state_4_last_state <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_entry_BB_reg <= 0;
		end else begin
			if (andOp_272_out) begin
				state_5_entry_BB_reg <= 32'd20;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_is_active <= 0;
		end else begin
			if (andOp_272_out) begin
				state_5_is_active <= 1'd1;
			end
			if (andOp_293_out) begin
				state_5_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_last_BB_reg <= 0;
		end else begin
			if (andOp_272_out) begin
				state_5_last_BB_reg <= bb_20_predecessor_in_state_4_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_last_state <= 0;
		end else begin
			if (andOp_272_out) begin
				state_5_last_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_entry_BB_reg <= 0;
		end else begin
			if (andOp_106_out) begin
				state_6_entry_BB_reg <= 32'd22;
			end
			if (andOp_273_out) begin
				state_6_entry_BB_reg <= 32'd20;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_is_active <= 0;
		end else begin
			if (andOp_106_out) begin
				state_6_is_active <= 1'd1;
			end
			if (andOp_273_out) begin
				state_6_is_active <= 1'd1;
			end
			if (andOp_297_out) begin
				state_6_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_last_BB_reg <= 0;
		end else begin
			if (andOp_106_out) begin
				state_6_last_BB_reg <= 32'd22;
			end
			if (andOp_273_out) begin
				state_6_last_BB_reg <= bb_20_predecessor_in_state_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_last_state <= 0;
		end else begin
			if (andOp_106_out) begin
				state_6_last_state <= 32'd6;
			end
			if (andOp_273_out) begin
				state_6_last_state <= 32'd5;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_entry_BB_reg <= 0;
		end else begin
			if (andOp_104_out) begin
				state_7_entry_BB_reg <= 32'd23;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_is_active <= 0;
		end else begin
			if (andOp_104_out) begin
				state_7_is_active <= 1'd1;
			end
			if (andOp_299_out) begin
				state_7_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_last_BB_reg <= 0;
		end else begin
			if (andOp_104_out) begin
				state_7_last_BB_reg <= 32'd22;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_last_state <= 0;
		end else begin
			if (andOp_104_out) begin
				state_7_last_state <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_8_entry_BB_reg <= 0;
		end else begin
			if (andOp_122_out) begin
				state_8_entry_BB_reg <= 32'd10;
			end
			if (andOp_138_out) begin
				state_8_entry_BB_reg <= 32'd1;
			end
			if (andOp_274_out) begin
				state_8_entry_BB_reg <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_8_is_active <= 1;
		end else begin
			if (andOp_122_out) begin
				state_8_is_active <= 1'd1;
			end
			if (andOp_138_out) begin
				state_8_is_active <= 1'd1;
			end
			if (andOp_274_out) begin
				state_8_is_active <= 1'd1;
			end
			if (andOp_305_out) begin
				state_8_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_8_last_BB_reg <= 0;
		end else begin
			if (andOp_122_out) begin
				state_8_last_BB_reg <= 32'd10;
			end
			if (andOp_138_out) begin
				state_8_last_BB_reg <= 32'd3;
			end
			if (andOp_274_out) begin
				state_8_last_BB_reg <= 32'd7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_8_last_state <= 0;
		end else begin
			if (andOp_122_out) begin
				state_8_last_state <= 32'd8;
			end
			if (andOp_138_out) begin
				state_8_last_state <= 32'd12;
			end
			if (andOp_274_out) begin
				state_8_last_state <= 32'd7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_9_entry_BB_reg <= 0;
		end else begin
			if (andOp_120_out) begin
				state_9_entry_BB_reg <= 32'd11;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_9_is_active <= 0;
		end else begin
			if (andOp_120_out) begin
				state_9_is_active <= 1'd1;
			end
			if (andOp_307_out) begin
				state_9_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_9_last_BB_reg <= 0;
		end else begin
			if (andOp_120_out) begin
				state_9_last_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_9_last_state <= 0;
		end else begin
			if (andOp_120_out) begin
				state_9_last_state <= 32'd8;
			end
		end
	end

endmodule

