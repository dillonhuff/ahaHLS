module axi_wb(input [0:0] clk, input [0:0] rst, output [0:0] valid, output [31:0] arg_0_in_data, input [31:0] arg_0_out_data, input [0:0] arg_0_read_ready, output [0:0] arg_0_read_valid, input [0:0] arg_0_write_ready, output [0:0] arg_0_write_valid, output [7:0] arg_1_raddr, input [7:0] arg_1_rdata, output [7:0] arg_1_waddr, output [7:0] arg_1_wdata, output [0:0] arg_1_wen, output [15:0] arg_2_raddr, input [15:0] arg_2_rdata, output [15:0] arg_2_waddr, output [15:0] arg_2_wdata, output [0:0] arg_2_wen, output [15:0] arg_3_s_axi_araddr, output [1:0] arg_3_s_axi_arburst, output [7:0] arg_3_s_axi_arlen, input [0:0] arg_3_s_axi_arready, output [2:0] arg_3_s_axi_arsize, output [0:0] arg_3_s_axi_arvalid, output [15:0] arg_3_s_axi_awaddr, output [1:0] arg_3_s_axi_awburst, output [7:0] arg_3_s_axi_awlen, input [0:0] arg_3_s_axi_awready, output [2:0] arg_3_s_axi_awsize, output [0:0] arg_3_s_axi_awvalid, output [0:0] arg_3_s_axi_bready, input [0:0] arg_3_s_axi_bvalid, input [31:0] arg_3_s_axi_rdata, output [0:0] arg_3_s_axi_rready, input [0:0] arg_3_s_axi_rvalid, output [31:0] arg_3_s_axi_wdata, input [0:0] arg_3_s_axi_wready, output [3:0] arg_3_s_axi_wstrb, output [0:0] arg_3_s_axi_wvalid);

	reg [0:0] valid_reg;
	reg [31:0] arg_0_in_data_reg;
	reg [0:0] arg_0_read_valid_reg;
	reg [0:0] arg_0_write_valid_reg;
	reg [7:0] arg_1_raddr_reg;
	reg [7:0] arg_1_waddr_reg;
	reg [7:0] arg_1_wdata_reg;
	reg [0:0] arg_1_wen_reg;
	reg [15:0] arg_2_raddr_reg;
	reg [15:0] arg_2_waddr_reg;
	reg [15:0] arg_2_wdata_reg;
	reg [0:0] arg_2_wen_reg;
	reg [15:0] arg_3_s_axi_araddr_reg;
	reg [1:0] arg_3_s_axi_arburst_reg;
	reg [7:0] arg_3_s_axi_arlen_reg;
	reg [2:0] arg_3_s_axi_arsize_reg;
	reg [0:0] arg_3_s_axi_arvalid_reg;
	reg [15:0] arg_3_s_axi_awaddr_reg;
	reg [1:0] arg_3_s_axi_awburst_reg;
	reg [7:0] arg_3_s_axi_awlen_reg;
	reg [2:0] arg_3_s_axi_awsize_reg;
	reg [0:0] arg_3_s_axi_awvalid_reg;
	reg [0:0] arg_3_s_axi_bready_reg;
	reg [0:0] arg_3_s_axi_rready_reg;
	reg [31:0] arg_3_s_axi_wdata_reg;
	reg [3:0] arg_3_s_axi_wstrb_reg;
	reg [0:0] arg_3_s_axi_wvalid_reg;

	assign valid = valid_reg;
	assign arg_0_in_data = arg_0_in_data_reg;
	assign arg_0_read_valid = arg_0_read_valid_reg;
	assign arg_0_write_valid = arg_0_write_valid_reg;
	assign arg_1_raddr = arg_1_raddr_reg;
	assign arg_1_waddr = arg_1_waddr_reg;
	assign arg_1_wdata = arg_1_wdata_reg;
	assign arg_1_wen = arg_1_wen_reg;
	assign arg_2_raddr = arg_2_raddr_reg;
	assign arg_2_waddr = arg_2_waddr_reg;
	assign arg_2_wdata = arg_2_wdata_reg;
	assign arg_2_wen = arg_2_wen_reg;
	assign arg_3_s_axi_araddr = arg_3_s_axi_araddr_reg;
	assign arg_3_s_axi_arburst = arg_3_s_axi_arburst_reg;
	assign arg_3_s_axi_arlen = arg_3_s_axi_arlen_reg;
	assign arg_3_s_axi_arsize = arg_3_s_axi_arsize_reg;
	assign arg_3_s_axi_arvalid = arg_3_s_axi_arvalid_reg;
	assign arg_3_s_axi_awaddr = arg_3_s_axi_awaddr_reg;
	assign arg_3_s_axi_awburst = arg_3_s_axi_awburst_reg;
	assign arg_3_s_axi_awlen = arg_3_s_axi_awlen_reg;
	assign arg_3_s_axi_awsize = arg_3_s_axi_awsize_reg;
	assign arg_3_s_axi_awvalid = arg_3_s_axi_awvalid_reg;
	assign arg_3_s_axi_bready = arg_3_s_axi_bready_reg;
	assign arg_3_s_axi_rready = arg_3_s_axi_rready_reg;
	assign arg_3_s_axi_wdata = arg_3_s_axi_wdata_reg;
	assign arg_3_s_axi_wstrb = arg_3_s_axi_wstrb_reg;
	assign arg_3_s_axi_wvalid = arg_3_s_axi_wvalid_reg;

	// Start debug wires and ports

	initial begin
	end





	// End debug wires and ports

	// Start Functional Units
	wire [31:0] sext_sext0_in;
	wire [63:0] sext_sext0_out;
	sext sext_sext0(.in(sext_sext0_in), .out(sext_sext0_out));

	br_dummy br_unit();

	wire [31:0] sext_sext8_in;
	wire [63:0] sext_sext8_out;
	sext sext_sext8(.in(sext_sext8_in), .out(sext_sext8_out));

	wire [31:0] icmp_icmp9_in0;
	wire [31:0] icmp_icmp9_in1;
	wire [0:0] icmp_icmp9_out;
	eq #(.WIDTH(32)) icmp_icmp9(.in0(icmp_icmp9_in0), .in1(icmp_icmp9_in1), .out(icmp_icmp9_out));

	wire [31:0] icmp_icmp13_in0;
	wire [31:0] icmp_icmp13_in1;
	wire [0:0] icmp_icmp13_out;
	eq #(.WIDTH(32)) icmp_icmp13(.in0(icmp_icmp13_in0), .in1(icmp_icmp13_in1), .out(icmp_icmp13_out));

	wire [15:0] phi_phi14_in;
	wire [31:0] phi_phi14_last_block;
	wire [63:0] phi_phi14_s;
	wire [31:0] phi_phi14_out;
	phi #(.NB_PAIR(2), .WIDTH(8)) phi_phi14(.in(phi_phi14_in), .last_block(phi_phi14_last_block), .out(phi_phi14_out), .s(phi_phi14_s));

	add call33();

	wire [31:0] sext_sext27_in;
	wire [63:0] sext_sext27_out;
	sext sext_sext27(.in(sext_sext27_in), .out(sext_sext27_out));

	wire [31:0] icmp_icmp28_in0;
	wire [31:0] icmp_icmp28_in1;
	wire [0:0] icmp_icmp28_out;
	eq #(.WIDTH(32)) icmp_icmp28(.in0(icmp_icmp28_in0), .in1(icmp_icmp28_in1), .out(icmp_icmp28_out));

	wire [31:0] sext_sext30_in;
	wire [63:0] sext_sext30_out;
	sext sext_sext30(.in(sext_sext30_in), .out(sext_sext30_out));

	wire [7:0] icmp_icmp35_in0;
	wire [7:0] icmp_icmp35_in1;
	wire [0:0] icmp_icmp35_out;
	slt #(.WIDTH(8)) icmp_icmp35(.in0(icmp_icmp35_in0), .in1(icmp_icmp35_in1), .out(icmp_icmp35_out));

	wire [31:0] add_add31_in0;
	wire [31:0] add_add31_in1;
	wire [31:0] add_add31_out;
	add #(.WIDTH(32)) add_add31(.in0(add_add31_in0), .in1(add_add31_in1), .out(add_add31_out));

	wire [31:0] trunc_trunc32_in;
	wire [7:0] trunc_trunc32_out;
	trunc #(.IN_WIDTH(32), .OUT_WIDTH(8)) trunc_trunc32(.in(trunc_trunc32_in), .out(trunc_trunc32_out));

	reg [0:0] bb_3_active_in_state_0_in_data;
	wire [0:0] bb_3_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_0(.in_data(bb_3_active_in_state_0_in_data), .out_data(bb_3_active_in_state_0_out_data));

	reg [31:0] bb_3_predecessor_in_state_0_in_data;
	wire [31:0] bb_3_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_0(.in_data(bb_3_predecessor_in_state_0_in_data), .out_data(bb_3_predecessor_in_state_0_out_data));

	reg [0:0] br_3_happened_in_state_0_in_data;
	wire [0:0] br_3_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_0(.in_data(br_3_happened_in_state_0_in_data), .out_data(br_3_happened_in_state_0_out_data));

	reg [0:0] bb_4_active_in_state_0_in_data;
	wire [0:0] bb_4_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_0(.in_data(bb_4_active_in_state_0_in_data), .out_data(bb_4_active_in_state_0_out_data));

	reg [31:0] bb_4_predecessor_in_state_0_in_data;
	wire [31:0] bb_4_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_0(.in_data(bb_4_predecessor_in_state_0_in_data), .out_data(bb_4_predecessor_in_state_0_out_data));

	reg [0:0] br_4_happened_in_state_0_in_data;
	wire [0:0] br_4_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_0(.in_data(br_4_happened_in_state_0_in_data), .out_data(br_4_happened_in_state_0_out_data));

	reg [0:0] bb_5_active_in_state_0_in_data;
	wire [0:0] bb_5_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_5_active_in_state_0(.in_data(bb_5_active_in_state_0_in_data), .out_data(bb_5_active_in_state_0_out_data));

	reg [31:0] bb_5_predecessor_in_state_0_in_data;
	wire [31:0] bb_5_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_5_predecessor_in_state_0(.in_data(bb_5_predecessor_in_state_0_in_data), .out_data(bb_5_predecessor_in_state_0_out_data));

	reg [0:0] br_5_happened_in_state_0_in_data;
	wire [0:0] br_5_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_5_happened_in_state_0(.in_data(br_5_happened_in_state_0_in_data), .out_data(br_5_happened_in_state_0_out_data));

	reg [0:0] bb_1_active_in_state_0_in_data;
	wire [0:0] bb_1_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_0(.in_data(bb_1_active_in_state_0_in_data), .out_data(bb_1_active_in_state_0_out_data));

	reg [31:0] bb_1_predecessor_in_state_0_in_data;
	wire [31:0] bb_1_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_0(.in_data(bb_1_predecessor_in_state_0_in_data), .out_data(bb_1_predecessor_in_state_0_out_data));

	reg [0:0] br_1_happened_in_state_0_in_data;
	wire [0:0] br_1_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened_in_state_0(.in_data(br_1_happened_in_state_0_in_data), .out_data(br_1_happened_in_state_0_out_data));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] bb_6_active_in_state_1_in_data;
	wire [0:0] bb_6_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_6_active_in_state_1(.in_data(bb_6_active_in_state_1_in_data), .out_data(bb_6_active_in_state_1_out_data));

	reg [31:0] bb_6_predecessor_in_state_1_in_data;
	wire [31:0] bb_6_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_6_predecessor_in_state_1(.in_data(bb_6_predecessor_in_state_1_in_data), .out_data(bb_6_predecessor_in_state_1_out_data));

	reg [0:0] br_6_happened_in_state_1_in_data;
	wire [0:0] br_6_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_6_happened_in_state_1(.in_data(br_6_happened_in_state_1_in_data), .out_data(br_6_happened_in_state_1_out_data));

	reg [0:0] bb_6_active_in_state_2_in_data;
	wire [0:0] bb_6_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_6_active_in_state_2(.in_data(bb_6_active_in_state_2_in_data), .out_data(bb_6_active_in_state_2_out_data));

	reg [31:0] bb_6_predecessor_in_state_2_in_data;
	wire [31:0] bb_6_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_6_predecessor_in_state_2(.in_data(bb_6_predecessor_in_state_2_in_data), .out_data(bb_6_predecessor_in_state_2_out_data));

	reg [0:0] br_6_happened_in_state_2_in_data;
	wire [0:0] br_6_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_6_happened_in_state_2(.in_data(br_6_happened_in_state_2_in_data), .out_data(br_6_happened_in_state_2_out_data));

	reg [0:0] bb_7_active_in_state_2_in_data;
	wire [0:0] bb_7_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_7_active_in_state_2(.in_data(bb_7_active_in_state_2_in_data), .out_data(bb_7_active_in_state_2_out_data));

	reg [31:0] bb_7_predecessor_in_state_2_in_data;
	wire [31:0] bb_7_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_7_predecessor_in_state_2(.in_data(bb_7_predecessor_in_state_2_in_data), .out_data(bb_7_predecessor_in_state_2_out_data));

	reg [0:0] br_7_happened_in_state_2_in_data;
	wire [0:0] br_7_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_7_happened_in_state_2(.in_data(br_7_happened_in_state_2_in_data), .out_data(br_7_happened_in_state_2_out_data));

	reg [0:0] bb_8_active_in_state_2_in_data;
	wire [0:0] bb_8_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active_in_state_2(.in_data(bb_8_active_in_state_2_in_data), .out_data(bb_8_active_in_state_2_out_data));

	reg [31:0] bb_8_predecessor_in_state_2_in_data;
	wire [31:0] bb_8_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor_in_state_2(.in_data(bb_8_predecessor_in_state_2_in_data), .out_data(bb_8_predecessor_in_state_2_out_data));

	reg [0:0] br_8_happened_in_state_2_in_data;
	wire [0:0] br_8_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_8_happened_in_state_2(.in_data(br_8_happened_in_state_2_in_data), .out_data(br_8_happened_in_state_2_out_data));

	reg [0:0] bb_8_active_in_state_3_in_data;
	wire [0:0] bb_8_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active_in_state_3(.in_data(bb_8_active_in_state_3_in_data), .out_data(bb_8_active_in_state_3_out_data));

	reg [31:0] bb_8_predecessor_in_state_3_in_data;
	wire [31:0] bb_8_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor_in_state_3(.in_data(bb_8_predecessor_in_state_3_in_data), .out_data(bb_8_predecessor_in_state_3_out_data));

	reg [0:0] br_8_happened_in_state_3_in_data;
	wire [0:0] br_8_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_8_happened_in_state_3(.in_data(br_8_happened_in_state_3_in_data), .out_data(br_8_happened_in_state_3_out_data));

	reg [0:0] bb_2_active_in_state_3_in_data;
	wire [0:0] bb_2_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_3(.in_data(bb_2_active_in_state_3_in_data), .out_data(bb_2_active_in_state_3_out_data));

	reg [31:0] bb_2_predecessor_in_state_3_in_data;
	wire [31:0] bb_2_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_3(.in_data(bb_2_predecessor_in_state_3_in_data), .out_data(bb_2_predecessor_in_state_3_out_data));

	reg [0:0] bb_2_active_in_state_4_in_data;
	wire [0:0] bb_2_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_4(.in_data(bb_2_active_in_state_4_in_data), .out_data(bb_2_active_in_state_4_out_data));

	reg [31:0] bb_2_predecessor_in_state_4_in_data;
	wire [31:0] bb_2_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_4(.in_data(bb_2_predecessor_in_state_4_in_data), .out_data(bb_2_predecessor_in_state_4_out_data));

	reg [0:0] bb_2_active_in_state_5_in_data;
	wire [0:0] bb_2_active_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_5(.in_data(bb_2_active_in_state_5_in_data), .out_data(bb_2_active_in_state_5_out_data));

	reg [31:0] bb_2_predecessor_in_state_5_in_data;
	wire [31:0] bb_2_predecessor_in_state_5_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_5(.in_data(bb_2_predecessor_in_state_5_in_data), .out_data(bb_2_predecessor_in_state_5_out_data));

	reg [7:0] data_in_0_1_in_data;
	wire [7:0] data_in_0_1_out_data;
	hls_wire #(.WIDTH(8)) data_in_0_1(.in_data(data_in_0_1_in_data), .out_data(data_in_0_1_out_data));

	reg [31:0] data_in_0_3_in_data;
	wire [31:0] data_in_0_3_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_3(.in_data(data_in_0_3_in_data), .out_data(data_in_0_3_out_data));

	reg [15:0] data_in_0_5_in_data;
	wire [15:0] data_in_0_5_out_data;
	hls_wire #(.WIDTH(16)) data_in_0_5(.in_data(data_in_0_5_in_data), .out_data(data_in_0_5_out_data));

	reg [7:0] data_in_0_7_in_data;
	wire [7:0] data_in_0_7_out_data;
	hls_wire #(.WIDTH(8)) data_in_0_7(.in_data(data_in_0_7_in_data), .out_data(data_in_0_7_out_data));

	reg [7:0] data_in_0_9_in_data;
	wire [7:0] data_in_0_9_out_data;
	hls_wire #(.WIDTH(8)) data_in_0_9(.in_data(data_in_0_9_in_data), .out_data(data_in_0_9_out_data));

	reg [7:0] data_in_1_11_in_data;
	wire [7:0] data_in_1_11_out_data;
	hls_wire #(.WIDTH(8)) data_in_1_11(.in_data(data_in_1_11_in_data), .out_data(data_in_1_11_out_data));

	reg [31:0] data_in_1_13_in_data;
	wire [31:0] data_in_1_13_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_13(.in_data(data_in_1_13_in_data), .out_data(data_in_1_13_out_data));

	reg [15:0] data_in_1_15_in_data;
	wire [15:0] data_in_1_15_out_data;
	hls_wire #(.WIDTH(16)) data_in_1_15(.in_data(data_in_1_15_in_data), .out_data(data_in_1_15_out_data));

	reg [7:0] data_in_1_17_in_data;
	wire [7:0] data_in_1_17_out_data;
	hls_wire #(.WIDTH(8)) data_in_1_17(.in_data(data_in_1_17_in_data), .out_data(data_in_1_17_out_data));

	reg [7:0] data_in_1_19_in_data;
	wire [7:0] data_in_1_19_out_data;
	hls_wire #(.WIDTH(8)) data_in_1_19(.in_data(data_in_1_19_in_data), .out_data(data_in_1_19_out_data));

	reg [7:0] data_in_2_21_in_data;
	wire [7:0] data_in_2_21_out_data;
	hls_wire #(.WIDTH(8)) data_in_2_21(.in_data(data_in_2_21_in_data), .out_data(data_in_2_21_out_data));

	reg [31:0] data_in_2_23_in_data;
	wire [31:0] data_in_2_23_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_23(.in_data(data_in_2_23_in_data), .out_data(data_in_2_23_out_data));

	reg [15:0] data_in_2_25_in_data;
	wire [15:0] data_in_2_25_out_data;
	hls_wire #(.WIDTH(16)) data_in_2_25(.in_data(data_in_2_25_in_data), .out_data(data_in_2_25_out_data));

	reg [7:0] data_in_2_27_in_data;
	wire [7:0] data_in_2_27_out_data;
	hls_wire #(.WIDTH(8)) data_in_2_27(.in_data(data_in_2_27_in_data), .out_data(data_in_2_27_out_data));

	reg [7:0] data_in_2_29_in_data;
	wire [7:0] data_in_2_29_out_data;
	hls_wire #(.WIDTH(8)) data_in_2_29(.in_data(data_in_2_29_in_data), .out_data(data_in_2_29_out_data));

	reg [7:0] data_in_3_31_in_data;
	wire [7:0] data_in_3_31_out_data;
	hls_wire #(.WIDTH(8)) data_in_3_31(.in_data(data_in_3_31_in_data), .out_data(data_in_3_31_out_data));

	reg [31:0] data_in_3_33_in_data;
	wire [31:0] data_in_3_33_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_33(.in_data(data_in_3_33_in_data), .out_data(data_in_3_33_out_data));

	reg [15:0] data_in_3_35_in_data;
	wire [15:0] data_in_3_35_out_data;
	hls_wire #(.WIDTH(16)) data_in_3_35(.in_data(data_in_3_35_in_data), .out_data(data_in_3_35_out_data));

	reg [7:0] data_in_3_37_in_data;
	wire [7:0] data_in_3_37_out_data;
	hls_wire #(.WIDTH(8)) data_in_3_37(.in_data(data_in_3_37_in_data), .out_data(data_in_3_37_out_data));

	reg [7:0] data_in_3_39_in_data;
	wire [7:0] data_in_3_39_out_data;
	hls_wire #(.WIDTH(8)) data_in_3_39(.in_data(data_in_3_39_in_data), .out_data(data_in_3_39_out_data));

	wire [0:0] andOp_40_in0;
	wire [0:0] andOp_40_in1;
	wire [0:0] andOp_40_out;
	andOp #(.WIDTH(1)) andOp_40(.in0(andOp_40_in0), .in1(andOp_40_in1), .out(andOp_40_out));

	wire [0:0] notOp_41_in0;
	wire [0:0] notOp_41_out;
	notOp #(.WIDTH(1)) notOp_41(.in(notOp_41_in0), .out(notOp_41_out));

	wire [0:0] andOp_42_in0;
	wire [0:0] andOp_42_in1;
	wire [0:0] andOp_42_out;
	andOp #(.WIDTH(1)) andOp_42(.in0(andOp_42_in0), .in1(andOp_42_in1), .out(andOp_42_out));

	wire [0:0] notOp_43_in0;
	wire [0:0] notOp_43_out;
	notOp #(.WIDTH(1)) notOp_43(.in(notOp_43_in0), .out(notOp_43_out));

	wire [0:0] andOp_44_in0;
	wire [0:0] andOp_44_in1;
	wire [0:0] andOp_44_out;
	andOp #(.WIDTH(1)) andOp_44(.in0(andOp_44_in0), .in1(andOp_44_in1), .out(andOp_44_out));

	wire [0:0] andOp_45_in0;
	wire [0:0] andOp_45_in1;
	wire [0:0] andOp_45_out;
	andOp #(.WIDTH(1)) andOp_45(.in0(andOp_45_in0), .in1(andOp_45_in1), .out(andOp_45_out));

	wire [0:0] notOp_46_in0;
	wire [0:0] notOp_46_out;
	notOp #(.WIDTH(1)) notOp_46(.in(notOp_46_in0), .out(notOp_46_out));

	wire [0:0] andOp_47_in0;
	wire [0:0] andOp_47_in1;
	wire [0:0] andOp_47_out;
	andOp #(.WIDTH(1)) andOp_47(.in0(andOp_47_in0), .in1(andOp_47_in1), .out(andOp_47_out));

	wire [0:0] notOp_48_in0;
	wire [0:0] notOp_48_out;
	notOp #(.WIDTH(1)) notOp_48(.in(notOp_48_in0), .out(notOp_48_out));

	wire [0:0] andOp_49_in0;
	wire [0:0] andOp_49_in1;
	wire [0:0] andOp_49_out;
	andOp #(.WIDTH(1)) andOp_49(.in0(andOp_49_in0), .in1(andOp_49_in1), .out(andOp_49_out));

	wire [0:0] notOp_50_in0;
	wire [0:0] notOp_50_out;
	notOp #(.WIDTH(1)) notOp_50(.in(notOp_50_in0), .out(notOp_50_out));

	wire [0:0] andOp_51_in0;
	wire [0:0] andOp_51_in1;
	wire [0:0] andOp_51_out;
	andOp #(.WIDTH(1)) andOp_51(.in0(andOp_51_in0), .in1(andOp_51_in1), .out(andOp_51_out));

	wire [0:0] andOp_52_in0;
	wire [0:0] andOp_52_in1;
	wire [0:0] andOp_52_out;
	andOp #(.WIDTH(1)) andOp_52(.in0(andOp_52_in0), .in1(andOp_52_in1), .out(andOp_52_out));

	wire [0:0] notOp_53_in0;
	wire [0:0] notOp_53_out;
	notOp #(.WIDTH(1)) notOp_53(.in(notOp_53_in0), .out(notOp_53_out));

	wire [0:0] andOp_54_in0;
	wire [0:0] andOp_54_in1;
	wire [0:0] andOp_54_out;
	andOp #(.WIDTH(1)) andOp_54(.in0(andOp_54_in0), .in1(andOp_54_in1), .out(andOp_54_out));

	wire [0:0] notOp_55_in0;
	wire [0:0] notOp_55_out;
	notOp #(.WIDTH(1)) notOp_55(.in(notOp_55_in0), .out(notOp_55_out));

	wire [0:0] andOp_56_in0;
	wire [0:0] andOp_56_in1;
	wire [0:0] andOp_56_out;
	andOp #(.WIDTH(1)) andOp_56(.in0(andOp_56_in0), .in1(andOp_56_in1), .out(andOp_56_out));

	wire [0:0] notOp_57_in0;
	wire [0:0] notOp_57_out;
	notOp #(.WIDTH(1)) notOp_57(.in(notOp_57_in0), .out(notOp_57_out));

	wire [0:0] andOp_58_in0;
	wire [0:0] andOp_58_in1;
	wire [0:0] andOp_58_out;
	andOp #(.WIDTH(1)) andOp_58(.in0(andOp_58_in0), .in1(andOp_58_in1), .out(andOp_58_out));

	wire [0:0] notOp_59_in0;
	wire [0:0] notOp_59_out;
	notOp #(.WIDTH(1)) notOp_59(.in(notOp_59_in0), .out(notOp_59_out));

	wire [0:0] andOp_60_in0;
	wire [0:0] andOp_60_in1;
	wire [0:0] andOp_60_out;
	andOp #(.WIDTH(1)) andOp_60(.in0(andOp_60_in0), .in1(andOp_60_in1), .out(andOp_60_out));

	wire [0:0] notOp_61_in0;
	wire [0:0] notOp_61_out;
	notOp #(.WIDTH(1)) notOp_61(.in(notOp_61_in0), .out(notOp_61_out));

	wire [0:0] andOp_62_in0;
	wire [0:0] andOp_62_in1;
	wire [0:0] andOp_62_out;
	andOp #(.WIDTH(1)) andOp_62(.in0(andOp_62_in0), .in1(andOp_62_in1), .out(andOp_62_out));

	wire [0:0] notOp_63_in0;
	wire [0:0] notOp_63_out;
	notOp #(.WIDTH(1)) notOp_63(.in(notOp_63_in0), .out(notOp_63_out));

	wire [0:0] andOp_64_in0;
	wire [0:0] andOp_64_in1;
	wire [0:0] andOp_64_out;
	andOp #(.WIDTH(1)) andOp_64(.in0(andOp_64_in0), .in1(andOp_64_in1), .out(andOp_64_out));

	wire [0:0] andOp_65_in0;
	wire [0:0] andOp_65_in1;
	wire [0:0] andOp_65_out;
	andOp #(.WIDTH(1)) andOp_65(.in0(andOp_65_in0), .in1(andOp_65_in1), .out(andOp_65_out));

	wire [0:0] notOp_66_in0;
	wire [0:0] notOp_66_out;
	notOp #(.WIDTH(1)) notOp_66(.in(notOp_66_in0), .out(notOp_66_out));

	wire [0:0] andOp_67_in0;
	wire [0:0] andOp_67_in1;
	wire [0:0] andOp_67_out;
	andOp #(.WIDTH(1)) andOp_67(.in0(andOp_67_in0), .in1(andOp_67_in1), .out(andOp_67_out));

	wire [0:0] notOp_68_in0;
	wire [0:0] notOp_68_out;
	notOp #(.WIDTH(1)) notOp_68(.in(notOp_68_in0), .out(notOp_68_out));

	wire [0:0] andOp_69_in0;
	wire [0:0] andOp_69_in1;
	wire [0:0] andOp_69_out;
	andOp #(.WIDTH(1)) andOp_69(.in0(andOp_69_in0), .in1(andOp_69_in1), .out(andOp_69_out));

	wire [0:0] andOp_70_in0;
	wire [0:0] andOp_70_in1;
	wire [0:0] andOp_70_out;
	andOp #(.WIDTH(1)) andOp_70(.in0(andOp_70_in0), .in1(andOp_70_in1), .out(andOp_70_out));

	wire [0:0] notOp_71_in0;
	wire [0:0] notOp_71_out;
	notOp #(.WIDTH(1)) notOp_71(.in(notOp_71_in0), .out(notOp_71_out));

	wire [0:0] andOp_72_in0;
	wire [0:0] andOp_72_in1;
	wire [0:0] andOp_72_out;
	andOp #(.WIDTH(1)) andOp_72(.in0(andOp_72_in0), .in1(andOp_72_in1), .out(andOp_72_out));

	wire [0:0] notOp_73_in0;
	wire [0:0] notOp_73_out;
	notOp #(.WIDTH(1)) notOp_73(.in(notOp_73_in0), .out(notOp_73_out));

	wire [0:0] andOp_74_in0;
	wire [0:0] andOp_74_in1;
	wire [0:0] andOp_74_out;
	andOp #(.WIDTH(1)) andOp_74(.in0(andOp_74_in0), .in1(andOp_74_in1), .out(andOp_74_out));

	wire [31:0] eq_75_in0;
	wire [31:0] eq_75_in1;
	wire [0:0] eq_75_out;
	eq #(.WIDTH(32)) eq_75(.in0(eq_75_in0), .in1(eq_75_in1), .out(eq_75_out));

	wire [0:0] orOp_76_in0;
	wire [0:0] orOp_76_in1;
	wire [0:0] orOp_76_out;
	orOp #(.WIDTH(1)) orOp_76(.in0(orOp_76_in0), .in1(orOp_76_in1), .out(orOp_76_out));

	wire [31:0] eq_77_in0;
	wire [31:0] eq_77_in1;
	wire [0:0] eq_77_out;
	eq #(.WIDTH(32)) eq_77(.in0(eq_77_in0), .in1(eq_77_in1), .out(eq_77_out));

	wire [0:0] orOp_78_in0;
	wire [0:0] orOp_78_in1;
	wire [0:0] orOp_78_out;
	orOp #(.WIDTH(1)) orOp_78(.in0(orOp_78_in0), .in1(orOp_78_in1), .out(orOp_78_out));

	wire [31:0] eq_79_in0;
	wire [31:0] eq_79_in1;
	wire [0:0] eq_79_out;
	eq #(.WIDTH(32)) eq_79(.in0(eq_79_in0), .in1(eq_79_in1), .out(eq_79_out));

	wire [0:0] orOp_80_in0;
	wire [0:0] orOp_80_in1;
	wire [0:0] orOp_80_out;
	orOp #(.WIDTH(1)) orOp_80(.in0(orOp_80_in0), .in1(orOp_80_in1), .out(orOp_80_out));

	wire [31:0] eq_81_in0;
	wire [31:0] eq_81_in1;
	wire [0:0] eq_81_out;
	eq #(.WIDTH(32)) eq_81(.in0(eq_81_in0), .in1(eq_81_in1), .out(eq_81_out));

	wire [0:0] orOp_82_in0;
	wire [0:0] orOp_82_in1;
	wire [0:0] orOp_82_out;
	orOp #(.WIDTH(1)) orOp_82(.in0(orOp_82_in0), .in1(orOp_82_in1), .out(orOp_82_out));

	wire [31:0] eq_83_in0;
	wire [31:0] eq_83_in1;
	wire [0:0] eq_83_out;
	eq #(.WIDTH(32)) eq_83(.in0(eq_83_in0), .in1(eq_83_in1), .out(eq_83_out));

	wire [31:0] eq_84_in0;
	wire [31:0] eq_84_in1;
	wire [0:0] eq_84_out;
	eq #(.WIDTH(32)) eq_84(.in0(eq_84_in0), .in1(eq_84_in1), .out(eq_84_out));

	wire [31:0] eq_85_in0;
	wire [31:0] eq_85_in1;
	wire [0:0] eq_85_out;
	eq #(.WIDTH(32)) eq_85(.in0(eq_85_in0), .in1(eq_85_in1), .out(eq_85_out));

	wire [31:0] eq_86_in0;
	wire [31:0] eq_86_in1;
	wire [0:0] eq_86_out;
	eq #(.WIDTH(32)) eq_86(.in0(eq_86_in0), .in1(eq_86_in1), .out(eq_86_out));

	wire [0:0] orOp_87_in0;
	wire [0:0] orOp_87_in1;
	wire [0:0] orOp_87_out;
	orOp #(.WIDTH(1)) orOp_87(.in0(orOp_87_in0), .in1(orOp_87_in1), .out(orOp_87_out));

	wire [31:0] eq_88_in0;
	wire [31:0] eq_88_in1;
	wire [0:0] eq_88_out;
	eq #(.WIDTH(32)) eq_88(.in0(eq_88_in0), .in1(eq_88_in1), .out(eq_88_out));

	wire [0:0] orOp_89_in0;
	wire [0:0] orOp_89_in1;
	wire [0:0] orOp_89_out;
	orOp #(.WIDTH(1)) orOp_89(.in0(orOp_89_in0), .in1(orOp_89_in1), .out(orOp_89_out));

	wire [31:0] eq_90_in0;
	wire [31:0] eq_90_in1;
	wire [0:0] eq_90_out;
	eq #(.WIDTH(32)) eq_90(.in0(eq_90_in0), .in1(eq_90_in1), .out(eq_90_out));

	wire [31:0] eq_91_in0;
	wire [31:0] eq_91_in1;
	wire [0:0] eq_91_out;
	eq #(.WIDTH(32)) eq_91(.in0(eq_91_in0), .in1(eq_91_in1), .out(eq_91_out));

	wire [0:0] orOp_92_in0;
	wire [0:0] orOp_92_in1;
	wire [0:0] orOp_92_out;
	orOp #(.WIDTH(1)) orOp_92(.in0(orOp_92_in0), .in1(orOp_92_in1), .out(orOp_92_out));

	wire [31:0] eq_93_in0;
	wire [31:0] eq_93_in1;
	wire [0:0] eq_93_out;
	eq #(.WIDTH(32)) eq_93(.in0(eq_93_in0), .in1(eq_93_in1), .out(eq_93_out));

	wire [31:0] eq_94_in0;
	wire [31:0] eq_94_in1;
	wire [0:0] eq_94_out;
	eq #(.WIDTH(32)) eq_94(.in0(eq_94_in0), .in1(eq_94_in1), .out(eq_94_out));

	wire [31:0] eq_95_in0;
	wire [31:0] eq_95_in1;
	wire [0:0] eq_95_out;
	eq #(.WIDTH(32)) eq_95(.in0(eq_95_in0), .in1(eq_95_in1), .out(eq_95_out));

	wire [0:0] notOp_96_in0;
	wire [0:0] notOp_96_out;
	notOp #(.WIDTH(1)) notOp_96(.in(notOp_96_in0), .out(notOp_96_out));

	wire [0:0] andOp_97_in0;
	wire [0:0] andOp_97_in1;
	wire [0:0] andOp_97_out;
	andOp #(.WIDTH(1)) andOp_97(.in0(andOp_97_in0), .in1(andOp_97_in1), .out(andOp_97_out));

	wire [31:0] eq_98_in0;
	wire [31:0] eq_98_in1;
	wire [0:0] eq_98_out;
	eq #(.WIDTH(32)) eq_98(.in0(eq_98_in0), .in1(eq_98_in1), .out(eq_98_out));

	wire [0:0] notOp_99_in0;
	wire [0:0] notOp_99_out;
	notOp #(.WIDTH(1)) notOp_99(.in(notOp_99_in0), .out(notOp_99_out));

	wire [0:0] andOp_100_in0;
	wire [0:0] andOp_100_in1;
	wire [0:0] andOp_100_out;
	andOp #(.WIDTH(1)) andOp_100(.in0(andOp_100_in0), .in1(andOp_100_in1), .out(andOp_100_out));

	wire [31:0] eq_101_in0;
	wire [31:0] eq_101_in1;
	wire [0:0] eq_101_out;
	eq #(.WIDTH(32)) eq_101(.in0(eq_101_in0), .in1(eq_101_in1), .out(eq_101_out));

	wire [0:0] notOp_102_in0;
	wire [0:0] notOp_102_out;
	notOp #(.WIDTH(1)) notOp_102(.in(notOp_102_in0), .out(notOp_102_out));

	wire [0:0] andOp_103_in0;
	wire [0:0] andOp_103_in1;
	wire [0:0] andOp_103_out;
	andOp #(.WIDTH(1)) andOp_103(.in0(andOp_103_in0), .in1(andOp_103_in1), .out(andOp_103_out));

	wire [31:0] eq_104_in0;
	wire [31:0] eq_104_in1;
	wire [0:0] eq_104_out;
	eq #(.WIDTH(32)) eq_104(.in0(eq_104_in0), .in1(eq_104_in1), .out(eq_104_out));

	wire [0:0] notOp_105_in0;
	wire [0:0] notOp_105_out;
	notOp #(.WIDTH(1)) notOp_105(.in(notOp_105_in0), .out(notOp_105_out));

	wire [0:0] andOp_106_in0;
	wire [0:0] andOp_106_in1;
	wire [0:0] andOp_106_out;
	andOp #(.WIDTH(1)) andOp_106(.in0(andOp_106_in0), .in1(andOp_106_in1), .out(andOp_106_out));

	wire [31:0] eq_107_in0;
	wire [31:0] eq_107_in1;
	wire [0:0] eq_107_out;
	eq #(.WIDTH(32)) eq_107(.in0(eq_107_in0), .in1(eq_107_in1), .out(eq_107_out));

	wire [31:0] eq_108_in0;
	wire [31:0] eq_108_in1;
	wire [0:0] eq_108_out;
	eq #(.WIDTH(32)) eq_108(.in0(eq_108_in0), .in1(eq_108_in1), .out(eq_108_out));

	wire [31:0] eq_109_in0;
	wire [31:0] eq_109_in1;
	wire [0:0] eq_109_out;
	eq #(.WIDTH(32)) eq_109(.in0(eq_109_in0), .in1(eq_109_in1), .out(eq_109_out));

	wire [31:0] eq_110_in0;
	wire [31:0] eq_110_in1;
	wire [0:0] eq_110_out;
	eq #(.WIDTH(32)) eq_110(.in0(eq_110_in0), .in1(eq_110_in1), .out(eq_110_out));

	wire [0:0] notOp_111_in0;
	wire [0:0] notOp_111_out;
	notOp #(.WIDTH(1)) notOp_111(.in(notOp_111_in0), .out(notOp_111_out));

	wire [0:0] andOp_112_in0;
	wire [0:0] andOp_112_in1;
	wire [0:0] andOp_112_out;
	andOp #(.WIDTH(1)) andOp_112(.in0(andOp_112_in0), .in1(andOp_112_in1), .out(andOp_112_out));

	wire [31:0] eq_113_in0;
	wire [31:0] eq_113_in1;
	wire [0:0] eq_113_out;
	eq #(.WIDTH(32)) eq_113(.in0(eq_113_in0), .in1(eq_113_in1), .out(eq_113_out));

	wire [0:0] notOp_114_in0;
	wire [0:0] notOp_114_out;
	notOp #(.WIDTH(1)) notOp_114(.in(notOp_114_in0), .out(notOp_114_out));

	wire [0:0] andOp_115_in0;
	wire [0:0] andOp_115_in1;
	wire [0:0] andOp_115_out;
	andOp #(.WIDTH(1)) andOp_115(.in0(andOp_115_in0), .in1(andOp_115_in1), .out(andOp_115_out));

	wire [31:0] eq_116_in0;
	wire [31:0] eq_116_in1;
	wire [0:0] eq_116_out;
	eq #(.WIDTH(32)) eq_116(.in0(eq_116_in0), .in1(eq_116_in1), .out(eq_116_out));

	wire [31:0] eq_117_in0;
	wire [31:0] eq_117_in1;
	wire [0:0] eq_117_out;
	eq #(.WIDTH(32)) eq_117(.in0(eq_117_in0), .in1(eq_117_in1), .out(eq_117_out));

	wire [0:0] notOp_118_in0;
	wire [0:0] notOp_118_out;
	notOp #(.WIDTH(1)) notOp_118(.in(notOp_118_in0), .out(notOp_118_out));

	wire [0:0] andOp_119_in0;
	wire [0:0] andOp_119_in1;
	wire [0:0] andOp_119_out;
	andOp #(.WIDTH(1)) andOp_119(.in0(andOp_119_in0), .in1(andOp_119_in1), .out(andOp_119_out));

	wire [31:0] eq_120_in0;
	wire [31:0] eq_120_in1;
	wire [0:0] eq_120_out;
	eq #(.WIDTH(32)) eq_120(.in0(eq_120_in0), .in1(eq_120_in1), .out(eq_120_out));

	wire [31:0] eq_121_in0;
	wire [31:0] eq_121_in1;
	wire [0:0] eq_121_out;
	eq #(.WIDTH(32)) eq_121(.in0(eq_121_in0), .in1(eq_121_in1), .out(eq_121_out));

	wire [0:0] andOp_122_in0;
	wire [0:0] andOp_122_in1;
	wire [0:0] andOp_122_out;
	andOp #(.WIDTH(1)) andOp_122(.in0(andOp_122_in0), .in1(andOp_122_in1), .out(andOp_122_out));

	wire [0:0] andOp_123_in0;
	wire [0:0] andOp_123_in1;
	wire [0:0] andOp_123_out;
	andOp #(.WIDTH(1)) andOp_123(.in0(andOp_123_in0), .in1(andOp_123_in1), .out(andOp_123_out));

	reg [7:0] tmp_output_124_in_data;
	wire [7:0] tmp_output_124_out_data;
	hls_wire #(.WIDTH(8)) tmp_output_124(.in_data(tmp_output_124_in_data), .out_data(tmp_output_124_out_data));

	wire [31:0] eq_125_in0;
	wire [31:0] eq_125_in1;
	wire [0:0] eq_125_out;
	eq #(.WIDTH(32)) eq_125(.in0(eq_125_in0), .in1(eq_125_in1), .out(eq_125_out));

	wire [31:0] eq_126_in0;
	wire [31:0] eq_126_in1;
	wire [0:0] eq_126_out;
	eq #(.WIDTH(32)) eq_126(.in0(eq_126_in0), .in1(eq_126_in1), .out(eq_126_out));

	wire [31:0] eq_127_in0;
	wire [31:0] eq_127_in1;
	wire [0:0] eq_127_out;
	eq #(.WIDTH(32)) eq_127(.in0(eq_127_in0), .in1(eq_127_in1), .out(eq_127_out));

	wire [31:0] eq_128_in0;
	wire [31:0] eq_128_in1;
	wire [0:0] eq_128_out;
	eq #(.WIDTH(32)) eq_128(.in0(eq_128_in0), .in1(eq_128_in1), .out(eq_128_out));

	wire [0:0] andOp_129_in0;
	wire [0:0] andOp_129_in1;
	wire [0:0] andOp_129_out;
	andOp #(.WIDTH(1)) andOp_129(.in0(andOp_129_in0), .in1(andOp_129_in1), .out(andOp_129_out));

	wire [0:0] andOp_130_in0;
	wire [0:0] andOp_130_in1;
	wire [0:0] andOp_130_out;
	andOp #(.WIDTH(1)) andOp_130(.in0(andOp_130_in0), .in1(andOp_130_in1), .out(andOp_130_out));

	wire [0:0] andOp_131_in0;
	wire [0:0] andOp_131_in1;
	wire [0:0] andOp_131_out;
	andOp #(.WIDTH(1)) andOp_131(.in0(andOp_131_in0), .in1(andOp_131_in1), .out(andOp_131_out));

	reg [15:0] tmp_output_132_in_data;
	wire [15:0] tmp_output_132_out_data;
	hls_wire #(.WIDTH(16)) tmp_output_132(.in_data(tmp_output_132_in_data), .out_data(tmp_output_132_out_data));

	wire [31:0] eq_133_in0;
	wire [31:0] eq_133_in1;
	wire [0:0] eq_133_out;
	eq #(.WIDTH(32)) eq_133(.in0(eq_133_in0), .in1(eq_133_in1), .out(eq_133_out));

	wire [31:0] eq_134_in0;
	wire [31:0] eq_134_in1;
	wire [0:0] eq_134_out;
	eq #(.WIDTH(32)) eq_134(.in0(eq_134_in0), .in1(eq_134_in1), .out(eq_134_out));

	wire [31:0] eq_135_in0;
	wire [31:0] eq_135_in1;
	wire [0:0] eq_135_out;
	eq #(.WIDTH(32)) eq_135(.in0(eq_135_in0), .in1(eq_135_in1), .out(eq_135_out));

	wire [31:0] eq_136_in0;
	wire [31:0] eq_136_in1;
	wire [0:0] eq_136_out;
	eq #(.WIDTH(32)) eq_136(.in0(eq_136_in0), .in1(eq_136_in1), .out(eq_136_out));

	wire [0:0] andOp_137_in0;
	wire [0:0] andOp_137_in1;
	wire [0:0] andOp_137_out;
	andOp #(.WIDTH(1)) andOp_137(.in0(andOp_137_in0), .in1(andOp_137_in1), .out(andOp_137_out));

	wire [0:0] andOp_138_in0;
	wire [0:0] andOp_138_in1;
	wire [0:0] andOp_138_out;
	andOp #(.WIDTH(1)) andOp_138(.in0(andOp_138_in0), .in1(andOp_138_in1), .out(andOp_138_out));

	wire [0:0] andOp_139_in0;
	wire [0:0] andOp_139_in1;
	wire [0:0] andOp_139_out;
	andOp #(.WIDTH(1)) andOp_139(.in0(andOp_139_in0), .in1(andOp_139_in1), .out(andOp_139_out));

	wire [0:0] andOp_140_in0;
	wire [0:0] andOp_140_in1;
	wire [0:0] andOp_140_out;
	andOp #(.WIDTH(1)) andOp_140(.in0(andOp_140_in0), .in1(andOp_140_in1), .out(andOp_140_out));

	wire [0:0] andOp_141_in0;
	wire [0:0] andOp_141_in1;
	wire [0:0] andOp_141_out;
	andOp #(.WIDTH(1)) andOp_141(.in0(andOp_141_in0), .in1(andOp_141_in1), .out(andOp_141_out));

	wire [0:0] andOp_142_in0;
	wire [0:0] andOp_142_in1;
	wire [0:0] andOp_142_out;
	andOp #(.WIDTH(1)) andOp_142(.in0(andOp_142_in0), .in1(andOp_142_in1), .out(andOp_142_out));

	reg [31:0] tmp_output_143_in_data;
	wire [31:0] tmp_output_143_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_143(.in_data(tmp_output_143_in_data), .out_data(tmp_output_143_out_data));

	wire [31:0] eq_144_in0;
	wire [31:0] eq_144_in1;
	wire [0:0] eq_144_out;
	eq #(.WIDTH(32)) eq_144(.in0(eq_144_in0), .in1(eq_144_in1), .out(eq_144_out));

	wire [31:0] eq_145_in0;
	wire [31:0] eq_145_in1;
	wire [0:0] eq_145_out;
	eq #(.WIDTH(32)) eq_145(.in0(eq_145_in0), .in1(eq_145_in1), .out(eq_145_out));

	wire [0:0] andOp_146_in0;
	wire [0:0] andOp_146_in1;
	wire [0:0] andOp_146_out;
	andOp #(.WIDTH(1)) andOp_146(.in0(andOp_146_in0), .in1(andOp_146_in1), .out(andOp_146_out));

	wire [0:0] andOp_147_in0;
	wire [0:0] andOp_147_in1;
	wire [0:0] andOp_147_out;
	andOp #(.WIDTH(1)) andOp_147(.in0(andOp_147_in0), .in1(andOp_147_in1), .out(andOp_147_out));

	wire [0:0] andOp_148_in0;
	wire [0:0] andOp_148_in1;
	wire [0:0] andOp_148_out;
	andOp #(.WIDTH(1)) andOp_148(.in0(andOp_148_in0), .in1(andOp_148_in1), .out(andOp_148_out));

	wire [0:0] andOp_149_in0;
	wire [0:0] andOp_149_in1;
	wire [0:0] andOp_149_out;
	andOp #(.WIDTH(1)) andOp_149(.in0(andOp_149_in0), .in1(andOp_149_in1), .out(andOp_149_out));

	wire [0:0] andOp_150_in0;
	wire [0:0] andOp_150_in1;
	wire [0:0] andOp_150_out;
	andOp #(.WIDTH(1)) andOp_150(.in0(andOp_150_in0), .in1(andOp_150_in1), .out(andOp_150_out));

	wire [0:0] andOp_151_in0;
	wire [0:0] andOp_151_in1;
	wire [0:0] andOp_151_out;
	andOp #(.WIDTH(1)) andOp_151(.in0(andOp_151_in0), .in1(andOp_151_in1), .out(andOp_151_out));

	wire [0:0] andOp_152_in0;
	wire [0:0] andOp_152_in1;
	wire [0:0] andOp_152_out;
	andOp #(.WIDTH(1)) andOp_152(.in0(andOp_152_in0), .in1(andOp_152_in1), .out(andOp_152_out));

	wire [0:0] andOp_153_in0;
	wire [0:0] andOp_153_in1;
	wire [0:0] andOp_153_out;
	andOp #(.WIDTH(1)) andOp_153(.in0(andOp_153_in0), .in1(andOp_153_in1), .out(andOp_153_out));

	wire [0:0] andOp_154_in0;
	wire [0:0] andOp_154_in1;
	wire [0:0] andOp_154_out;
	andOp #(.WIDTH(1)) andOp_154(.in0(andOp_154_in0), .in1(andOp_154_in1), .out(andOp_154_out));

	wire [0:0] andOp_155_in0;
	wire [0:0] andOp_155_in1;
	wire [0:0] andOp_155_out;
	andOp #(.WIDTH(1)) andOp_155(.in0(andOp_155_in0), .in1(andOp_155_in1), .out(andOp_155_out));

	wire [0:0] andOp_156_in0;
	wire [0:0] andOp_156_in1;
	wire [0:0] andOp_156_out;
	andOp #(.WIDTH(1)) andOp_156(.in0(andOp_156_in0), .in1(andOp_156_in1), .out(andOp_156_out));

	wire [0:0] andOp_157_in0;
	wire [0:0] andOp_157_in1;
	wire [0:0] andOp_157_out;
	andOp #(.WIDTH(1)) andOp_157(.in0(andOp_157_in0), .in1(andOp_157_in1), .out(andOp_157_out));

	wire [7:0] concat_158_in0;
	wire [7:0] concat_158_in1;
	wire [15:0] concat_158_out;
	concat #(.IN0_WIDTH(8), .IN1_WIDTH(8)) concat_158(.in0(concat_158_in0), .in1(concat_158_in1), .out(concat_158_out));

	wire [31:0] concat_159_in0;
	wire [31:0] concat_159_in1;
	wire [63:0] concat_159_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_159(.in0(concat_159_in0), .in1(concat_159_in1), .out(concat_159_out));

	wire [0:0] andOp_160_in0;
	wire [0:0] andOp_160_in1;
	wire [0:0] andOp_160_out;
	andOp #(.WIDTH(1)) andOp_160(.in0(andOp_160_in0), .in1(andOp_160_in1), .out(andOp_160_out));

	wire [0:0] andOp_161_in0;
	wire [0:0] andOp_161_in1;
	wire [0:0] andOp_161_out;
	andOp #(.WIDTH(1)) andOp_161(.in0(andOp_161_in0), .in1(andOp_161_in1), .out(andOp_161_out));

	wire [0:0] andOp_162_in0;
	wire [0:0] andOp_162_in1;
	wire [0:0] andOp_162_out;
	andOp #(.WIDTH(1)) andOp_162(.in0(andOp_162_in0), .in1(andOp_162_in1), .out(andOp_162_out));

	wire [0:0] andOp_163_in0;
	wire [0:0] andOp_163_in1;
	wire [0:0] andOp_163_out;
	andOp #(.WIDTH(1)) andOp_163(.in0(andOp_163_in0), .in1(andOp_163_in1), .out(andOp_163_out));

	wire [0:0] andOp_164_in0;
	wire [0:0] andOp_164_in1;
	wire [0:0] andOp_164_out;
	andOp #(.WIDTH(1)) andOp_164(.in0(andOp_164_in0), .in1(andOp_164_in1), .out(andOp_164_out));

	wire [0:0] andOp_165_in0;
	wire [0:0] andOp_165_in1;
	wire [0:0] andOp_165_out;
	andOp #(.WIDTH(1)) andOp_165(.in0(andOp_165_in0), .in1(andOp_165_in1), .out(andOp_165_out));

	wire [0:0] andOp_166_in0;
	wire [0:0] andOp_166_in1;
	wire [0:0] andOp_166_out;
	andOp #(.WIDTH(1)) andOp_166(.in0(andOp_166_in0), .in1(andOp_166_in1), .out(andOp_166_out));

	wire [0:0] andOp_167_in0;
	wire [0:0] andOp_167_in1;
	wire [0:0] andOp_167_out;
	andOp #(.WIDTH(1)) andOp_167(.in0(andOp_167_in0), .in1(andOp_167_in1), .out(andOp_167_out));

	wire [0:0] andOp_168_in0;
	wire [0:0] andOp_168_in1;
	wire [0:0] andOp_168_out;
	andOp #(.WIDTH(1)) andOp_168(.in0(andOp_168_in0), .in1(andOp_168_in1), .out(andOp_168_out));

	wire [0:0] andOp_169_in0;
	wire [0:0] andOp_169_in1;
	wire [0:0] andOp_169_out;
	andOp #(.WIDTH(1)) andOp_169(.in0(andOp_169_in0), .in1(andOp_169_in1), .out(andOp_169_out));

	wire [0:0] andOp_170_in0;
	wire [0:0] andOp_170_in1;
	wire [0:0] andOp_170_out;
	andOp #(.WIDTH(1)) andOp_170(.in0(andOp_170_in0), .in1(andOp_170_in1), .out(andOp_170_out));

	wire [0:0] andOp_171_in0;
	wire [0:0] andOp_171_in1;
	wire [0:0] andOp_171_out;
	andOp #(.WIDTH(1)) andOp_171(.in0(andOp_171_in0), .in1(andOp_171_in1), .out(andOp_171_out));

	wire [0:0] andOp_172_in0;
	wire [0:0] andOp_172_in1;
	wire [0:0] andOp_172_out;
	andOp #(.WIDTH(1)) andOp_172(.in0(andOp_172_in0), .in1(andOp_172_in1), .out(andOp_172_out));

	wire [0:0] andOp_173_in0;
	wire [0:0] andOp_173_in1;
	wire [0:0] andOp_173_out;
	andOp #(.WIDTH(1)) andOp_173(.in0(andOp_173_in0), .in1(andOp_173_in1), .out(andOp_173_out));

	wire [0:0] andOp_174_in0;
	wire [0:0] andOp_174_in1;
	wire [0:0] andOp_174_out;
	andOp #(.WIDTH(1)) andOp_174(.in0(andOp_174_in0), .in1(andOp_174_in1), .out(andOp_174_out));

	wire [0:0] notOp_175_in0;
	wire [0:0] notOp_175_out;
	notOp #(.WIDTH(1)) notOp_175(.in(notOp_175_in0), .out(notOp_175_out));

	wire [0:0] andOp_176_in0;
	wire [0:0] andOp_176_in1;
	wire [0:0] andOp_176_out;
	andOp #(.WIDTH(1)) andOp_176(.in0(andOp_176_in0), .in1(andOp_176_in1), .out(andOp_176_out));

	wire [0:0] notOp_177_in0;
	wire [0:0] notOp_177_out;
	notOp #(.WIDTH(1)) notOp_177(.in(notOp_177_in0), .out(notOp_177_out));

	wire [0:0] andOp_178_in0;
	wire [0:0] andOp_178_in1;
	wire [0:0] andOp_178_out;
	andOp #(.WIDTH(1)) andOp_178(.in0(andOp_178_in0), .in1(andOp_178_in1), .out(andOp_178_out));

	wire [0:0] notOp_179_in0;
	wire [0:0] notOp_179_out;
	notOp #(.WIDTH(1)) notOp_179(.in(notOp_179_in0), .out(notOp_179_out));

	wire [0:0] andOp_180_in0;
	wire [0:0] andOp_180_in1;
	wire [0:0] andOp_180_out;
	andOp #(.WIDTH(1)) andOp_180(.in0(andOp_180_in0), .in1(andOp_180_in1), .out(andOp_180_out));

	wire [0:0] notOp_181_in0;
	wire [0:0] notOp_181_out;
	notOp #(.WIDTH(1)) notOp_181(.in(notOp_181_in0), .out(notOp_181_out));

	wire [0:0] andOp_182_in0;
	wire [0:0] andOp_182_in1;
	wire [0:0] andOp_182_out;
	andOp #(.WIDTH(1)) andOp_182(.in0(andOp_182_in0), .in1(andOp_182_in1), .out(andOp_182_out));

	wire [0:0] notOp_183_in0;
	wire [0:0] notOp_183_out;
	notOp #(.WIDTH(1)) notOp_183(.in(notOp_183_in0), .out(notOp_183_out));

	wire [0:0] andOp_184_in0;
	wire [0:0] andOp_184_in1;
	wire [0:0] andOp_184_out;
	andOp #(.WIDTH(1)) andOp_184(.in0(andOp_184_in0), .in1(andOp_184_in1), .out(andOp_184_out));

	wire [0:0] notOp_185_in0;
	wire [0:0] notOp_185_out;
	notOp #(.WIDTH(1)) notOp_185(.in(notOp_185_in0), .out(notOp_185_out));

	wire [0:0] andOp_186_in0;
	wire [0:0] andOp_186_in1;
	wire [0:0] andOp_186_out;
	andOp #(.WIDTH(1)) andOp_186(.in0(andOp_186_in0), .in1(andOp_186_in1), .out(andOp_186_out));

	wire [0:0] notOp_187_in0;
	wire [0:0] notOp_187_out;
	notOp #(.WIDTH(1)) notOp_187(.in(notOp_187_in0), .out(notOp_187_out));

	wire [0:0] andOp_188_in0;
	wire [0:0] andOp_188_in1;
	wire [0:0] andOp_188_out;
	andOp #(.WIDTH(1)) andOp_188(.in0(andOp_188_in0), .in1(andOp_188_in1), .out(andOp_188_out));

	wire [0:0] notOp_189_in0;
	wire [0:0] notOp_189_out;
	notOp #(.WIDTH(1)) notOp_189(.in(notOp_189_in0), .out(notOp_189_out));

	wire [0:0] andOp_190_in0;
	wire [0:0] andOp_190_in1;
	wire [0:0] andOp_190_out;
	andOp #(.WIDTH(1)) andOp_190(.in0(andOp_190_in0), .in1(andOp_190_in1), .out(andOp_190_out));

	wire [0:0] notOp_191_in0;
	wire [0:0] notOp_191_out;
	notOp #(.WIDTH(1)) notOp_191(.in(notOp_191_in0), .out(notOp_191_out));

	wire [0:0] andOp_192_in0;
	wire [0:0] andOp_192_in1;
	wire [0:0] andOp_192_out;
	andOp #(.WIDTH(1)) andOp_192(.in0(andOp_192_in0), .in1(andOp_192_in1), .out(andOp_192_out));

	wire [0:0] notOp_193_in0;
	wire [0:0] notOp_193_out;
	notOp #(.WIDTH(1)) notOp_193(.in(notOp_193_in0), .out(notOp_193_out));

	wire [0:0] andOp_194_in0;
	wire [0:0] andOp_194_in1;
	wire [0:0] andOp_194_out;
	andOp #(.WIDTH(1)) andOp_194(.in0(andOp_194_in0), .in1(andOp_194_in1), .out(andOp_194_out));

	wire [31:0] eq_195_in0;
	wire [31:0] eq_195_in1;
	wire [0:0] eq_195_out;
	eq #(.WIDTH(32)) eq_195(.in0(eq_195_in0), .in1(eq_195_in1), .out(eq_195_out));

	wire [31:0] eq_196_in0;
	wire [31:0] eq_196_in1;
	wire [0:0] eq_196_out;
	eq #(.WIDTH(32)) eq_196(.in0(eq_196_in0), .in1(eq_196_in1), .out(eq_196_out));

	wire [0:0] andOp_197_in0;
	wire [0:0] andOp_197_in1;
	wire [0:0] andOp_197_out;
	andOp #(.WIDTH(1)) andOp_197(.in0(andOp_197_in0), .in1(andOp_197_in1), .out(andOp_197_out));

	wire [0:0] andOp_198_in0;
	wire [0:0] andOp_198_in1;
	wire [0:0] andOp_198_out;
	andOp #(.WIDTH(1)) andOp_198(.in0(andOp_198_in0), .in1(andOp_198_in1), .out(andOp_198_out));

	wire [0:0] andOp_199_in0;
	wire [0:0] andOp_199_in1;
	wire [0:0] andOp_199_out;
	andOp #(.WIDTH(1)) andOp_199(.in0(andOp_199_in0), .in1(andOp_199_in1), .out(andOp_199_out));

	wire [31:0] eq_200_in0;
	wire [31:0] eq_200_in1;
	wire [0:0] eq_200_out;
	eq #(.WIDTH(32)) eq_200(.in0(eq_200_in0), .in1(eq_200_in1), .out(eq_200_out));

	wire [31:0] eq_201_in0;
	wire [31:0] eq_201_in1;
	wire [0:0] eq_201_out;
	eq #(.WIDTH(32)) eq_201(.in0(eq_201_in0), .in1(eq_201_in1), .out(eq_201_out));

	wire [31:0] eq_202_in0;
	wire [31:0] eq_202_in1;
	wire [0:0] eq_202_out;
	eq #(.WIDTH(32)) eq_202(.in0(eq_202_in0), .in1(eq_202_in1), .out(eq_202_out));

	wire [31:0] eq_203_in0;
	wire [31:0] eq_203_in1;
	wire [0:0] eq_203_out;
	eq #(.WIDTH(32)) eq_203(.in0(eq_203_in0), .in1(eq_203_in1), .out(eq_203_out));

	wire [0:0] andOp_204_in0;
	wire [0:0] andOp_204_in1;
	wire [0:0] andOp_204_out;
	andOp #(.WIDTH(1)) andOp_204(.in0(andOp_204_in0), .in1(andOp_204_in1), .out(andOp_204_out));

	wire [0:0] andOp_205_in0;
	wire [0:0] andOp_205_in1;
	wire [0:0] andOp_205_out;
	andOp #(.WIDTH(1)) andOp_205(.in0(andOp_205_in0), .in1(andOp_205_in1), .out(andOp_205_out));

	wire [31:0] eq_206_in0;
	wire [31:0] eq_206_in1;
	wire [0:0] eq_206_out;
	eq #(.WIDTH(32)) eq_206(.in0(eq_206_in0), .in1(eq_206_in1), .out(eq_206_out));

	wire [31:0] eq_207_in0;
	wire [31:0] eq_207_in1;
	wire [0:0] eq_207_out;
	eq #(.WIDTH(32)) eq_207(.in0(eq_207_in0), .in1(eq_207_in1), .out(eq_207_out));

	wire [31:0] eq_208_in0;
	wire [31:0] eq_208_in1;
	wire [0:0] eq_208_out;
	eq #(.WIDTH(32)) eq_208(.in0(eq_208_in0), .in1(eq_208_in1), .out(eq_208_out));

	wire [31:0] eq_209_in0;
	wire [31:0] eq_209_in1;
	wire [0:0] eq_209_out;
	eq #(.WIDTH(32)) eq_209(.in0(eq_209_in0), .in1(eq_209_in1), .out(eq_209_out));

	wire [31:0] eq_210_in0;
	wire [31:0] eq_210_in1;
	wire [0:0] eq_210_out;
	eq #(.WIDTH(32)) eq_210(.in0(eq_210_in0), .in1(eq_210_in1), .out(eq_210_out));

	wire [31:0] eq_211_in0;
	wire [31:0] eq_211_in1;
	wire [0:0] eq_211_out;
	eq #(.WIDTH(32)) eq_211(.in0(eq_211_in0), .in1(eq_211_in1), .out(eq_211_out));

	// End Functional Units

	reg [7:0] data_store_0_0;
	reg [31:0] data_store_0_2;
	reg [15:0] data_store_0_4;
	reg [7:0] data_store_0_6;
	reg [7:0] data_store_0_8;
	reg [7:0] data_store_1_10;
	reg [31:0] data_store_1_12;
	reg [15:0] data_store_1_14;
	reg [7:0] data_store_1_16;
	reg [7:0] data_store_1_18;
	reg [7:0] data_store_2_20;
	reg [31:0] data_store_2_22;
	reg [15:0] data_store_2_24;
	reg [7:0] data_store_2_26;
	reg [7:0] data_store_2_28;
	reg [7:0] data_store_3_30;
	reg [31:0] data_store_3_32;
	reg [15:0] data_store_3_34;
	reg [7:0] data_store_3_36;
	reg [7:0] data_store_3_38;
	reg [31:0] global_state;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_3_last_state;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;
	reg [31:0] state_4_last_state;
	reg [31:0] state_5_entry_BB_reg;
	reg [0:0] state_5_is_active;
	reg [31:0] state_5_last_BB_reg;
	reg [31:0] state_5_last_state;

	// controller for add_add31.add_add31_in0
	// controller for add_add31.add_add31_in1
	// Insensitive connections
	assign add_add31_in0 = sext_sext30_out;
	assign add_add31_in1 = 32'd1;
	// controller for andOp_100.andOp_100_in0
	// controller for andOp_100.andOp_100_in1
	// Insensitive connections
	assign andOp_100_in0 = notOp_99_out;
	assign andOp_100_in1 = andOp_44_out;
	// controller for andOp_103.andOp_103_in0
	// controller for andOp_103.andOp_103_in1
	// Insensitive connections
	assign andOp_103_in0 = notOp_102_out;
	assign andOp_103_in1 = andOp_52_out;
	// controller for andOp_106.andOp_106_in0
	// controller for andOp_106.andOp_106_in1
	// Insensitive connections
	assign andOp_106_in0 = notOp_105_out;
	assign andOp_106_in1 = andOp_45_out;
	// controller for andOp_112.andOp_112_in0
	// controller for andOp_112.andOp_112_in1
	// Insensitive connections
	assign andOp_112_in0 = notOp_111_out;
	assign andOp_112_in1 = andOp_56_out;
	// controller for andOp_115.andOp_115_in0
	// controller for andOp_115.andOp_115_in1
	// Insensitive connections
	assign andOp_115_in0 = notOp_114_out;
	assign andOp_115_in1 = andOp_64_out;
	// controller for andOp_119.andOp_119_in0
	// controller for andOp_119.andOp_119_in1
	// Insensitive connections
	assign andOp_119_in0 = notOp_118_out;
	assign andOp_119_in1 = andOp_69_out;
	// controller for andOp_122.andOp_122_in0
	// controller for andOp_122.andOp_122_in1
	// Insensitive connections
	assign andOp_122_in0 = bb_5_active_in_state_0_out_data;
	assign andOp_122_in1 = state_0_is_active;
	// controller for andOp_123.andOp_123_in0
	// controller for andOp_123.andOp_123_in1
	// Insensitive connections
	assign andOp_123_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_123_in1 = state_0_is_active;
	// controller for andOp_129.andOp_129_in0
	// controller for andOp_129.andOp_129_in1
	// Insensitive connections
	assign andOp_129_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_129_in1 = state_0_is_active;
	// controller for andOp_130.andOp_130_in0
	// controller for andOp_130.andOp_130_in1
	// Insensitive connections
	assign andOp_130_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_130_in1 = state_0_is_active;
	// controller for andOp_131.andOp_131_in0
	// controller for andOp_131.andOp_131_in1
	// Insensitive connections
	assign andOp_131_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_131_in1 = state_0_is_active;
	// controller for andOp_137.andOp_137_in0
	// controller for andOp_137.andOp_137_in1
	// Insensitive connections
	assign andOp_137_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_137_in1 = state_0_is_active;
	// controller for andOp_138.andOp_138_in0
	// controller for andOp_138.andOp_138_in1
	// Insensitive connections
	assign andOp_138_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_138_in1 = state_0_is_active;
	// controller for andOp_139.andOp_139_in0
	// controller for andOp_139.andOp_139_in1
	// Insensitive connections
	assign andOp_139_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_139_in1 = state_0_is_active;
	// controller for andOp_140.andOp_140_in0
	// controller for andOp_140.andOp_140_in1
	// Insensitive connections
	assign andOp_140_in0 = bb_7_active_in_state_2_out_data;
	assign andOp_140_in1 = state_2_is_active;
	// controller for andOp_141.andOp_141_in0
	// controller for andOp_141.andOp_141_in1
	// Insensitive connections
	assign andOp_141_in0 = bb_7_active_in_state_2_out_data;
	assign andOp_141_in1 = state_2_is_active;
	// controller for andOp_142.andOp_142_in0
	// controller for andOp_142.andOp_142_in1
	// Insensitive connections
	assign andOp_142_in0 = bb_7_active_in_state_2_out_data;
	assign andOp_142_in1 = state_2_is_active;
	// controller for andOp_146.andOp_146_in0
	// controller for andOp_146.andOp_146_in1
	// Insensitive connections
	assign andOp_146_in0 = bb_7_active_in_state_2_out_data;
	assign andOp_146_in1 = state_2_is_active;
	// controller for andOp_147.andOp_147_in0
	// controller for andOp_147.andOp_147_in1
	// Insensitive connections
	assign andOp_147_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_147_in1 = state_3_is_active;
	// controller for andOp_148.andOp_148_in0
	// controller for andOp_148.andOp_148_in1
	// Insensitive connections
	assign andOp_148_in0 = bb_2_active_in_state_4_out_data;
	assign andOp_148_in1 = state_4_is_active;
	// controller for andOp_149.andOp_149_in0
	// controller for andOp_149.andOp_149_in1
	// Insensitive connections
	assign andOp_149_in0 = bb_2_active_in_state_4_out_data;
	assign andOp_149_in1 = state_4_is_active;
	// controller for andOp_150.andOp_150_in0
	// controller for andOp_150.andOp_150_in1
	// Insensitive connections
	assign andOp_150_in0 = bb_2_active_in_state_4_out_data;
	assign andOp_150_in1 = state_4_is_active;
	// controller for andOp_151.andOp_151_in0
	// controller for andOp_151.andOp_151_in1
	// Insensitive connections
	assign andOp_151_in0 = bb_5_active_in_state_0_out_data;
	assign andOp_151_in1 = state_0_is_active;
	// controller for andOp_152.andOp_152_in0
	// controller for andOp_152.andOp_152_in1
	// Insensitive connections
	assign andOp_152_in0 = bb_6_active_in_state_1_out_data;
	assign andOp_152_in1 = state_1_is_active;
	// controller for andOp_153.andOp_153_in0
	// controller for andOp_153.andOp_153_in1
	// Insensitive connections
	assign andOp_153_in0 = bb_6_active_in_state_2_out_data;
	assign andOp_153_in1 = state_2_is_active;
	// controller for andOp_154.andOp_154_in0
	// controller for andOp_154.andOp_154_in1
	// Insensitive connections
	assign andOp_154_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_154_in1 = state_0_is_active;
	// controller for andOp_155.andOp_155_in0
	// controller for andOp_155.andOp_155_in1
	// Insensitive connections
	assign andOp_155_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_155_in1 = state_0_is_active;
	// controller for andOp_156.andOp_156_in0
	// controller for andOp_156.andOp_156_in1
	// Insensitive connections
	assign andOp_156_in0 = bb_5_active_in_state_0_out_data;
	assign andOp_156_in1 = state_0_is_active;
	// controller for andOp_157.andOp_157_in0
	// controller for andOp_157.andOp_157_in1
	// Insensitive connections
	assign andOp_157_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_157_in1 = state_0_is_active;
	// controller for andOp_160.andOp_160_in0
	// controller for andOp_160.andOp_160_in1
	// Insensitive connections
	assign andOp_160_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_160_in1 = state_0_is_active;
	// controller for andOp_161.andOp_161_in0
	// controller for andOp_161.andOp_161_in1
	// Insensitive connections
	assign andOp_161_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_161_in1 = state_0_is_active;
	// controller for andOp_162.andOp_162_in0
	// controller for andOp_162.andOp_162_in1
	// Insensitive connections
	assign andOp_162_in0 = bb_7_active_in_state_2_out_data;
	assign andOp_162_in1 = state_2_is_active;
	// controller for andOp_163.andOp_163_in0
	// controller for andOp_163.andOp_163_in1
	// Insensitive connections
	assign andOp_163_in0 = bb_7_active_in_state_2_out_data;
	assign andOp_163_in1 = state_2_is_active;
	// controller for andOp_164.andOp_164_in0
	// controller for andOp_164.andOp_164_in1
	// Insensitive connections
	assign andOp_164_in0 = bb_8_active_in_state_2_out_data;
	assign andOp_164_in1 = state_2_is_active;
	// controller for andOp_165.andOp_165_in0
	// controller for andOp_165.andOp_165_in1
	// Insensitive connections
	assign andOp_165_in0 = bb_8_active_in_state_2_out_data;
	assign andOp_165_in1 = state_2_is_active;
	// controller for andOp_166.andOp_166_in0
	// controller for andOp_166.andOp_166_in1
	// Insensitive connections
	assign andOp_166_in0 = bb_8_active_in_state_2_out_data;
	assign andOp_166_in1 = state_2_is_active;
	// controller for andOp_167.andOp_167_in0
	// controller for andOp_167.andOp_167_in1
	// Insensitive connections
	assign andOp_167_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_167_in1 = state_3_is_active;
	// controller for andOp_168.andOp_168_in0
	// controller for andOp_168.andOp_168_in1
	// Insensitive connections
	assign andOp_168_in0 = bb_8_active_in_state_3_out_data;
	assign andOp_168_in1 = state_3_is_active;
	// controller for andOp_169.andOp_169_in0
	// controller for andOp_169.andOp_169_in1
	// Insensitive connections
	assign andOp_169_in0 = bb_2_active_in_state_5_out_data;
	assign andOp_169_in1 = state_5_is_active;
	// controller for andOp_170.andOp_170_in0
	// controller for andOp_170.andOp_170_in1
	// Insensitive connections
	assign andOp_170_in0 = bb_6_active_in_state_1_out_data;
	assign andOp_170_in1 = state_1_is_active;
	// controller for andOp_171.andOp_171_in0
	// controller for andOp_171.andOp_171_in1
	// Insensitive connections
	assign andOp_171_in0 = bb_8_active_in_state_2_out_data;
	assign andOp_171_in1 = state_2_is_active;
	// controller for andOp_172.andOp_172_in0
	// controller for andOp_172.andOp_172_in1
	// Insensitive connections
	assign andOp_172_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_172_in1 = state_3_is_active;
	// controller for andOp_173.andOp_173_in0
	// controller for andOp_173.andOp_173_in1
	// Insensitive connections
	assign andOp_173_in0 = bb_2_active_in_state_4_out_data;
	assign andOp_173_in1 = state_4_is_active;
	// controller for andOp_174.andOp_174_in0
	// controller for andOp_174.andOp_174_in1
	// Insensitive connections
	assign andOp_174_in0 = bb_2_active_in_state_5_out_data;
	assign andOp_174_in1 = state_5_is_active;
	// controller for andOp_176.andOp_176_in0
	// controller for andOp_176.andOp_176_in1
	// Insensitive connections
	assign andOp_176_in0 = notOp_175_out;
	assign andOp_176_in1 = 1'd1;
	// controller for andOp_178.andOp_178_in0
	// controller for andOp_178.andOp_178_in1
	// Insensitive connections
	assign andOp_178_in0 = notOp_177_out;
	assign andOp_178_in1 = andOp_176_out;
	// controller for andOp_180.andOp_180_in0
	// controller for andOp_180.andOp_180_in1
	// Insensitive connections
	assign andOp_180_in0 = notOp_179_out;
	assign andOp_180_in1 = andOp_178_out;
	// controller for andOp_182.andOp_182_in0
	// controller for andOp_182.andOp_182_in1
	// Insensitive connections
	assign andOp_182_in0 = notOp_181_out;
	assign andOp_182_in1 = 1'd1;
	// controller for andOp_184.andOp_184_in0
	// controller for andOp_184.andOp_184_in1
	// Insensitive connections
	assign andOp_184_in0 = notOp_183_out;
	assign andOp_184_in1 = 1'd1;
	// controller for andOp_186.andOp_186_in0
	// controller for andOp_186.andOp_186_in1
	// Insensitive connections
	assign andOp_186_in0 = notOp_185_out;
	assign andOp_186_in1 = andOp_184_out;
	// controller for andOp_188.andOp_188_in0
	// controller for andOp_188.andOp_188_in1
	// Insensitive connections
	assign andOp_188_in0 = notOp_187_out;
	assign andOp_188_in1 = 1'd1;
	// controller for andOp_190.andOp_190_in0
	// controller for andOp_190.andOp_190_in1
	// Insensitive connections
	assign andOp_190_in0 = notOp_189_out;
	assign andOp_190_in1 = 1'd1;
	// controller for andOp_192.andOp_192_in0
	// controller for andOp_192.andOp_192_in1
	// Insensitive connections
	assign andOp_192_in0 = notOp_191_out;
	assign andOp_192_in1 = 1'd1;
	// controller for andOp_194.andOp_194_in0
	// controller for andOp_194.andOp_194_in1
	// Insensitive connections
	assign andOp_194_in0 = notOp_193_out;
	assign andOp_194_in1 = andOp_192_out;
	// controller for andOp_197.andOp_197_in0
	// controller for andOp_197.andOp_197_in1
	// Insensitive connections
	assign andOp_197_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_197_in1 = state_0_is_active;
	// controller for andOp_198.andOp_198_in0
	// controller for andOp_198.andOp_198_in1
	// Insensitive connections
	assign andOp_198_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_198_in1 = state_0_is_active;
	// controller for andOp_199.andOp_199_in0
	// controller for andOp_199.andOp_199_in1
	// Insensitive connections
	assign andOp_199_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_199_in1 = state_0_is_active;
	// controller for andOp_204.andOp_204_in0
	// controller for andOp_204.andOp_204_in1
	// Insensitive connections
	assign andOp_204_in0 = bb_6_active_in_state_2_out_data;
	assign andOp_204_in1 = state_2_is_active;
	// controller for andOp_205.andOp_205_in0
	// controller for andOp_205.andOp_205_in1
	// Insensitive connections
	assign andOp_205_in0 = bb_8_active_in_state_2_out_data;
	assign andOp_205_in1 = state_2_is_active;
	// controller for andOp_40.andOp_40_in0
	// controller for andOp_40.andOp_40_in1
	// Insensitive connections
	assign andOp_40_in0 = bb_3_active_in_state_0_out_data;
	assign andOp_40_in1 = state_0_is_active;
	// controller for andOp_42.andOp_42_in0
	// controller for andOp_42.andOp_42_in1
	// Insensitive connections
	assign andOp_42_in0 = andOp_40_out;
	assign andOp_42_in1 = icmp_icmp9_out;
	// controller for andOp_44.andOp_44_in0
	// controller for andOp_44.andOp_44_in1
	// Insensitive connections
	assign andOp_44_in0 = andOp_40_out;
	assign andOp_44_in1 = notOp_43_out;
	// controller for andOp_45.andOp_45_in0
	// controller for andOp_45.andOp_45_in1
	// Insensitive connections
	assign andOp_45_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_45_in1 = state_0_is_active;
	// controller for andOp_47.andOp_47_in0
	// controller for andOp_47.andOp_47_in1
	// Insensitive connections
	assign andOp_47_in0 = bb_5_active_in_state_0_out_data;
	assign andOp_47_in1 = state_0_is_active;
	// controller for andOp_49.andOp_49_in0
	// controller for andOp_49.andOp_49_in1
	// Insensitive connections
	assign andOp_49_in0 = andOp_47_out;
	assign andOp_49_in1 = icmp_icmp13_out;
	// controller for andOp_51.andOp_51_in0
	// controller for andOp_51.andOp_51_in1
	// Insensitive connections
	assign andOp_51_in0 = andOp_47_out;
	assign andOp_51_in1 = notOp_50_out;
	// controller for andOp_52.andOp_52_in0
	// controller for andOp_52.andOp_52_in1
	// Insensitive connections
	assign andOp_52_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_52_in1 = state_0_is_active;
	// controller for andOp_54.andOp_54_in0
	// controller for andOp_54.andOp_54_in1
	// Insensitive connections
	assign andOp_54_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_54_in1 = state_0_is_active;
	// controller for andOp_56.andOp_56_in0
	// controller for andOp_56.andOp_56_in1
	// Insensitive connections
	assign andOp_56_in0 = bb_6_active_in_state_2_out_data;
	assign andOp_56_in1 = state_2_is_active;
	// controller for andOp_58.andOp_58_in0
	// controller for andOp_58.andOp_58_in1
	// Insensitive connections
	assign andOp_58_in0 = bb_6_active_in_state_2_out_data;
	assign andOp_58_in1 = state_2_is_active;
	// controller for andOp_60.andOp_60_in0
	// controller for andOp_60.andOp_60_in1
	// Insensitive connections
	assign andOp_60_in0 = bb_7_active_in_state_2_out_data;
	assign andOp_60_in1 = state_2_is_active;
	// controller for andOp_62.andOp_62_in0
	// controller for andOp_62.andOp_62_in1
	// Insensitive connections
	assign andOp_62_in0 = andOp_60_out;
	assign andOp_62_in1 = icmp_icmp28_out;
	// controller for andOp_64.andOp_64_in0
	// controller for andOp_64.andOp_64_in1
	// Insensitive connections
	assign andOp_64_in0 = andOp_60_out;
	assign andOp_64_in1 = notOp_63_out;
	// controller for andOp_65.andOp_65_in0
	// controller for andOp_65.andOp_65_in1
	// Insensitive connections
	assign andOp_65_in0 = bb_8_active_in_state_3_out_data;
	assign andOp_65_in1 = state_3_is_active;
	// controller for andOp_67.andOp_67_in0
	// controller for andOp_67.andOp_67_in1
	// Insensitive connections
	assign andOp_67_in0 = andOp_65_out;
	assign andOp_67_in1 = icmp_icmp35_out;
	// controller for andOp_69.andOp_69_in0
	// controller for andOp_69.andOp_69_in1
	// Insensitive connections
	assign andOp_69_in0 = andOp_65_out;
	assign andOp_69_in1 = notOp_68_out;
	// controller for andOp_70.andOp_70_in0
	// controller for andOp_70.andOp_70_in1
	// Insensitive connections
	assign andOp_70_in0 = bb_8_active_in_state_3_out_data;
	assign andOp_70_in1 = state_3_is_active;
	// controller for andOp_72.andOp_72_in0
	// controller for andOp_72.andOp_72_in1
	// Insensitive connections
	assign andOp_72_in0 = andOp_70_out;
	assign andOp_72_in1 = icmp_icmp35_out;
	// controller for andOp_74.andOp_74_in0
	// controller for andOp_74.andOp_74_in1
	// Insensitive connections
	assign andOp_74_in0 = andOp_70_out;
	assign andOp_74_in1 = notOp_73_out;
	// controller for andOp_97.andOp_97_in0
	// controller for andOp_97.andOp_97_in1
	// Insensitive connections
	assign andOp_97_in0 = notOp_96_out;
	assign andOp_97_in1 = andOp_54_out;
	// controller for arg_0.arg_0_read_valid_reg
	always @(*) begin
		if (andOp_152_out) begin 
			arg_0_read_valid_reg = 32'd1;
		end else begin
			arg_0_read_valid_reg = 0;
		end
	end
	// controller for arg_1.arg_1_raddr_reg
	always @(*) begin
		if (andOp_161_out) begin 
			arg_1_raddr_reg = arg_1_rdata;
		end else begin
			arg_1_raddr_reg = 0;
		end
	end
	// controller for arg_2.arg_2_raddr_reg
	always @(*) begin
		if (andOp_160_out) begin 
			arg_2_raddr_reg = arg_2_rdata;
		end else begin
			arg_2_raddr_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_awaddr_reg
	always @(*) begin
		if (andOp_131_out) begin 
			arg_3_s_axi_awaddr_reg = tmp_output_132_out_data;
		end else begin
			arg_3_s_axi_awaddr_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_awburst_reg
	always @(*) begin
		if (andOp_130_out) begin 
			arg_3_s_axi_awburst_reg = 2'd1;
		end else begin
			arg_3_s_axi_awburst_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_awlen_reg
	always @(*) begin
		if (andOp_123_out) begin 
			arg_3_s_axi_awlen_reg = tmp_output_124_out_data;
		end else begin
			arg_3_s_axi_awlen_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_awsize_reg
	always @(*) begin
		if (andOp_129_out) begin 
			arg_3_s_axi_awsize_reg = -(3'd3);
		end else begin
			arg_3_s_axi_awsize_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_awvalid_reg
	always @(*) begin
		if (andOp_138_out) begin 
			arg_3_s_axi_awvalid_reg = 32'd1;
		end else begin
			arg_3_s_axi_awvalid_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_wdata_reg
	always @(*) begin
		if (andOp_142_out) begin 
			arg_3_s_axi_wdata_reg = tmp_output_143_out_data;
		end else if (andOp_149_out) begin 
			arg_3_s_axi_wdata_reg = 32'd0;
		end else begin
			arg_3_s_axi_wdata_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_wstrb_reg
	always @(*) begin
		if (andOp_146_out) begin 
			arg_3_s_axi_wstrb_reg = -(4'd1);
		end else if (andOp_150_out) begin 
			arg_3_s_axi_wstrb_reg = 32'd0;
		end else begin
			arg_3_s_axi_wstrb_reg = 0;
		end
	end
	// controller for arg_3.arg_3_s_axi_wvalid_reg
	always @(*) begin
		if (andOp_137_out) begin 
			arg_3_s_axi_wvalid_reg = 32'd1;
		end else if (andOp_141_out) begin 
			arg_3_s_axi_wvalid_reg = 32'd1;
		end else if (andOp_148_out) begin 
			arg_3_s_axi_wvalid_reg = 32'd1;
		end else begin
			arg_3_s_axi_wvalid_reg = 0;
		end
	end
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_83_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_107_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_0.bb_1_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_0_in_data = orOp_82_out;
		end else begin
			bb_1_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_0.bb_1_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_106_out) begin 
			bb_1_predecessor_in_state_0_in_data = 32'd4;
		end else if (eq_104_out) begin 
			bb_1_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_3.bb_2_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_3_in_data = orOp_92_out;
		end else begin
			bb_2_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_4.bb_2_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_4_in_data = eq_93_out;
		end else begin
			bb_2_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_5.bb_2_active_in_state_5_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_5_in_data = eq_94_out;
		end else begin
			bb_2_active_in_state_5_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_3.bb_2_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_119_out) begin 
			bb_2_predecessor_in_state_3_in_data = 32'd8;
		end else if (eq_117_out) begin 
			bb_2_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_4.bb_2_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_120_out) begin 
			bb_2_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_5.bb_2_predecessor_in_state_5_in_data
	always @(*) begin
		if (eq_121_out) begin 
			bb_2_predecessor_in_state_5_in_data = state_5_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_5_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_0.bb_3_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_0_in_data = orOp_76_out;
		end else begin
			bb_3_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_0.bb_3_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_97_out) begin 
			bb_3_predecessor_in_state_0_in_data = 32'd0;
		end else if (eq_95_out) begin 
			bb_3_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_0.bb_4_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_0_in_data = orOp_78_out;
		end else begin
			bb_4_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_0.bb_4_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_100_out) begin 
			bb_4_predecessor_in_state_0_in_data = 32'd3;
		end else if (eq_98_out) begin 
			bb_4_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_5_active_in_state_0.bb_5_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_5_active_in_state_0_in_data = orOp_80_out;
		end else begin
			bb_5_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_5_predecessor_in_state_0.bb_5_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_103_out) begin 
			bb_5_predecessor_in_state_0_in_data = 32'd1;
		end else if (eq_101_out) begin 
			bb_5_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_5_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_6_active_in_state_1.bb_6_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_6_active_in_state_1_in_data = eq_84_out;
		end else begin
			bb_6_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_6_active_in_state_2.bb_6_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_6_active_in_state_2_in_data = eq_85_out;
		end else begin
			bb_6_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_6_predecessor_in_state_1.bb_6_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_108_out) begin 
			bb_6_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_6_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_6_predecessor_in_state_2.bb_6_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_109_out) begin 
			bb_6_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_6_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_7_active_in_state_2.bb_7_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_7_active_in_state_2_in_data = orOp_87_out;
		end else begin
			bb_7_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_7_predecessor_in_state_2.bb_7_predecessor_in_state_2_in_data
	always @(*) begin
		if (andOp_112_out) begin 
			bb_7_predecessor_in_state_2_in_data = 32'd6;
		end else if (eq_110_out) begin 
			bb_7_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_7_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_8_active_in_state_2.bb_8_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_state_2_in_data = orOp_89_out;
		end else begin
			bb_8_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_8_active_in_state_3.bb_8_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_state_3_in_data = eq_90_out;
		end else begin
			bb_8_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_8_predecessor_in_state_2.bb_8_predecessor_in_state_2_in_data
	always @(*) begin
		if (andOp_115_out) begin 
			bb_8_predecessor_in_state_2_in_data = 32'd7;
		end else if (eq_113_out) begin 
			bb_8_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_8_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_8_predecessor_in_state_3.bb_8_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_116_out) begin 
			bb_8_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_8_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_54_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_55_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_1_happened_in_state_0.br_1_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_52_out) begin 
			br_1_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_53_out) begin 
			br_1_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_1_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_0.br_3_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_40_out) begin 
			br_3_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_41_out) begin 
			br_3_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_0.br_4_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_45_out) begin 
			br_4_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_46_out) begin 
			br_4_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_5_happened_in_state_0.br_5_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_47_out) begin 
			br_5_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_48_out) begin 
			br_5_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_5_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_6_happened_in_state_1.br_6_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_56_out) begin 
			br_6_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_57_out) begin 
			br_6_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_6_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_6_happened_in_state_2.br_6_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_58_out) begin 
			br_6_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_59_out) begin 
			br_6_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_6_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_7_happened_in_state_2.br_7_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_60_out) begin 
			br_7_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_61_out) begin 
			br_7_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_7_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_8_happened_in_state_2.br_8_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_65_out) begin 
			br_8_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_66_out) begin 
			br_8_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_8_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_8_happened_in_state_3.br_8_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_70_out) begin 
			br_8_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_71_out) begin 
			br_8_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_8_happened_in_state_3_in_data = 0;
		end
	end
	// controller for concat_158.concat_158_in0
	// controller for concat_158.concat_158_in1
	// Insensitive connections
	assign concat_158_in0 = 8'd0;
	assign concat_158_in1 = data_in_0_9_out_data;
	// controller for concat_159.concat_159_in0
	// controller for concat_159.concat_159_in1
	// Insensitive connections
	assign concat_159_in0 = 32'd4;
	assign concat_159_in1 = 32'd8;
	// controller for data_in_0_1.data_in_0_1_in_data
	always @(*) begin
		if (eq_195_out) begin 
			data_in_0_1_in_data = data_store_0_0;
		end else if (eq_196_out) begin 
			data_in_0_1_in_data = data_store_3_30;
		end else begin
			data_in_0_1_in_data = 0;
		end
	end
	// controller for data_in_0_3.data_in_0_3_in_data
	always @(*) begin
		if (eq_195_out) begin 
			data_in_0_3_in_data = data_store_0_2;
		end else if (eq_196_out) begin 
			data_in_0_3_in_data = data_store_3_32;
		end else begin
			data_in_0_3_in_data = 0;
		end
	end
	// controller for data_in_0_5.data_in_0_5_in_data
	always @(*) begin
		if (eq_195_out) begin 
			data_in_0_5_in_data = data_store_0_4;
		end else if (eq_196_out) begin 
			data_in_0_5_in_data = data_store_3_34;
		end else begin
			data_in_0_5_in_data = 0;
		end
	end
	// controller for data_in_0_7.data_in_0_7_in_data
	always @(*) begin
		if (eq_195_out) begin 
			data_in_0_7_in_data = data_store_0_6;
		end else if (eq_196_out) begin 
			data_in_0_7_in_data = data_store_3_36;
		end else begin
			data_in_0_7_in_data = 0;
		end
	end
	// controller for data_in_0_9.data_in_0_9_in_data
	always @(*) begin
		if (eq_195_out) begin 
			data_in_0_9_in_data = data_store_0_8;
		end else if (eq_196_out) begin 
			data_in_0_9_in_data = data_store_3_38;
		end else begin
			data_in_0_9_in_data = 0;
		end
	end
	// controller for data_in_1_11.data_in_1_11_in_data
	always @(*) begin
		if (eq_200_out) begin 
			data_in_1_11_in_data = data_store_0_0;
		end else if (eq_201_out) begin 
			data_in_1_11_in_data = data_store_1_10;
		end else begin
			data_in_1_11_in_data = 0;
		end
	end
	// controller for data_in_1_13.data_in_1_13_in_data
	always @(*) begin
		if (eq_200_out) begin 
			data_in_1_13_in_data = data_store_0_2;
		end else if (eq_201_out) begin 
			data_in_1_13_in_data = data_store_1_12;
		end else begin
			data_in_1_13_in_data = 0;
		end
	end
	// controller for data_in_1_15.data_in_1_15_in_data
	always @(*) begin
		if (eq_200_out) begin 
			data_in_1_15_in_data = data_store_0_4;
		end else if (eq_201_out) begin 
			data_in_1_15_in_data = data_store_1_14;
		end else begin
			data_in_1_15_in_data = 0;
		end
	end
	// controller for data_in_1_17.data_in_1_17_in_data
	always @(*) begin
		if (eq_200_out) begin 
			data_in_1_17_in_data = data_store_0_6;
		end else if (eq_201_out) begin 
			data_in_1_17_in_data = data_store_1_16;
		end else begin
			data_in_1_17_in_data = 0;
		end
	end
	// controller for data_in_1_19.data_in_1_19_in_data
	always @(*) begin
		if (eq_200_out) begin 
			data_in_1_19_in_data = data_store_0_8;
		end else if (eq_201_out) begin 
			data_in_1_19_in_data = data_store_1_18;
		end else begin
			data_in_1_19_in_data = 0;
		end
	end
	// controller for data_in_2_21.data_in_2_21_in_data
	always @(*) begin
		if (eq_202_out) begin 
			data_in_2_21_in_data = data_store_1_10;
		end else if (eq_203_out) begin 
			data_in_2_21_in_data = data_store_2_20;
		end else begin
			data_in_2_21_in_data = 0;
		end
	end
	// controller for data_in_2_23.data_in_2_23_in_data
	always @(*) begin
		if (eq_202_out) begin 
			data_in_2_23_in_data = data_store_1_12;
		end else if (eq_203_out) begin 
			data_in_2_23_in_data = data_store_2_22;
		end else begin
			data_in_2_23_in_data = 0;
		end
	end
	// controller for data_in_2_25.data_in_2_25_in_data
	always @(*) begin
		if (eq_202_out) begin 
			data_in_2_25_in_data = data_store_1_14;
		end else if (eq_203_out) begin 
			data_in_2_25_in_data = data_store_2_24;
		end else begin
			data_in_2_25_in_data = 0;
		end
	end
	// controller for data_in_2_27.data_in_2_27_in_data
	always @(*) begin
		if (eq_202_out) begin 
			data_in_2_27_in_data = data_store_1_16;
		end else if (eq_203_out) begin 
			data_in_2_27_in_data = data_store_2_26;
		end else begin
			data_in_2_27_in_data = 0;
		end
	end
	// controller for data_in_2_29.data_in_2_29_in_data
	always @(*) begin
		if (eq_202_out) begin 
			data_in_2_29_in_data = data_store_1_18;
		end else if (eq_203_out) begin 
			data_in_2_29_in_data = data_store_2_28;
		end else begin
			data_in_2_29_in_data = 0;
		end
	end
	// controller for data_in_3_31.data_in_3_31_in_data
	always @(*) begin
		if (eq_206_out) begin 
			data_in_3_31_in_data = data_store_2_20;
		end else if (eq_207_out) begin 
			data_in_3_31_in_data = data_store_3_30;
		end else begin
			data_in_3_31_in_data = 0;
		end
	end
	// controller for data_in_3_33.data_in_3_33_in_data
	always @(*) begin
		if (eq_206_out) begin 
			data_in_3_33_in_data = data_store_2_22;
		end else if (eq_207_out) begin 
			data_in_3_33_in_data = data_store_3_32;
		end else begin
			data_in_3_33_in_data = 0;
		end
	end
	// controller for data_in_3_35.data_in_3_35_in_data
	always @(*) begin
		if (eq_206_out) begin 
			data_in_3_35_in_data = data_store_2_24;
		end else if (eq_207_out) begin 
			data_in_3_35_in_data = data_store_3_34;
		end else begin
			data_in_3_35_in_data = 0;
		end
	end
	// controller for data_in_3_37.data_in_3_37_in_data
	always @(*) begin
		if (eq_206_out) begin 
			data_in_3_37_in_data = data_store_2_26;
		end else if (eq_207_out) begin 
			data_in_3_37_in_data = data_store_3_36;
		end else begin
			data_in_3_37_in_data = 0;
		end
	end
	// controller for data_in_3_39.data_in_3_39_in_data
	always @(*) begin
		if (eq_206_out) begin 
			data_in_3_39_in_data = data_store_2_28;
		end else if (eq_207_out) begin 
			data_in_3_39_in_data = data_store_3_38;
		end else begin
			data_in_3_39_in_data = 0;
		end
	end
	// controller for eq_101.eq_101_in0
	// controller for eq_101.eq_101_in1
	// Insensitive connections
	assign eq_101_in0 = 32'd5;
	assign eq_101_in1 = state_0_entry_BB_reg;
	// controller for eq_104.eq_104_in0
	// controller for eq_104.eq_104_in1
	// Insensitive connections
	assign eq_104_in0 = 32'd1;
	assign eq_104_in1 = state_0_entry_BB_reg;
	// controller for eq_107.eq_107_in0
	// controller for eq_107.eq_107_in1
	// Insensitive connections
	assign eq_107_in0 = 32'd0;
	assign eq_107_in1 = state_0_entry_BB_reg;
	// controller for eq_108.eq_108_in0
	// controller for eq_108.eq_108_in1
	// Insensitive connections
	assign eq_108_in0 = 32'd6;
	assign eq_108_in1 = state_1_entry_BB_reg;
	// controller for eq_109.eq_109_in0
	// controller for eq_109.eq_109_in1
	// Insensitive connections
	assign eq_109_in0 = 32'd6;
	assign eq_109_in1 = state_2_entry_BB_reg;
	// controller for eq_110.eq_110_in0
	// controller for eq_110.eq_110_in1
	// Insensitive connections
	assign eq_110_in0 = 32'd7;
	assign eq_110_in1 = state_2_entry_BB_reg;
	// controller for eq_113.eq_113_in0
	// controller for eq_113.eq_113_in1
	// Insensitive connections
	assign eq_113_in0 = 32'd8;
	assign eq_113_in1 = state_2_entry_BB_reg;
	// controller for eq_116.eq_116_in0
	// controller for eq_116.eq_116_in1
	// Insensitive connections
	assign eq_116_in0 = 32'd8;
	assign eq_116_in1 = state_3_entry_BB_reg;
	// controller for eq_117.eq_117_in0
	// controller for eq_117.eq_117_in1
	// Insensitive connections
	assign eq_117_in0 = 32'd2;
	assign eq_117_in1 = state_3_entry_BB_reg;
	// controller for eq_120.eq_120_in0
	// controller for eq_120.eq_120_in1
	// Insensitive connections
	assign eq_120_in0 = 32'd2;
	assign eq_120_in1 = state_4_entry_BB_reg;
	// controller for eq_121.eq_121_in0
	// controller for eq_121.eq_121_in1
	// Insensitive connections
	assign eq_121_in0 = 32'd2;
	assign eq_121_in1 = state_5_entry_BB_reg;
	// controller for eq_125.eq_125_in0
	// controller for eq_125.eq_125_in1
	// Insensitive connections
	assign eq_125_in0 = 32'd3;
	assign eq_125_in1 = state_0_entry_BB_reg;
	// controller for eq_126.eq_126_in0
	// controller for eq_126.eq_126_in1
	// Insensitive connections
	assign eq_126_in0 = 32'd5;
	assign eq_126_in1 = state_0_entry_BB_reg;
	// controller for eq_127.eq_127_in0
	// controller for eq_127.eq_127_in1
	// Insensitive connections
	assign eq_127_in0 = 32'd1;
	assign eq_127_in1 = state_0_entry_BB_reg;
	// controller for eq_128.eq_128_in0
	// controller for eq_128.eq_128_in1
	// Insensitive connections
	assign eq_128_in0 = 32'd0;
	assign eq_128_in1 = state_0_entry_BB_reg;
	// controller for eq_133.eq_133_in0
	// controller for eq_133.eq_133_in1
	// Insensitive connections
	assign eq_133_in0 = 32'd3;
	assign eq_133_in1 = state_0_entry_BB_reg;
	// controller for eq_134.eq_134_in0
	// controller for eq_134.eq_134_in1
	// Insensitive connections
	assign eq_134_in0 = 32'd5;
	assign eq_134_in1 = state_0_entry_BB_reg;
	// controller for eq_135.eq_135_in0
	// controller for eq_135.eq_135_in1
	// Insensitive connections
	assign eq_135_in0 = 32'd1;
	assign eq_135_in1 = state_0_entry_BB_reg;
	// controller for eq_136.eq_136_in0
	// controller for eq_136.eq_136_in1
	// Insensitive connections
	assign eq_136_in0 = 32'd0;
	assign eq_136_in1 = state_0_entry_BB_reg;
	// controller for eq_144.eq_144_in0
	// controller for eq_144.eq_144_in1
	// Insensitive connections
	assign eq_144_in0 = 32'd6;
	assign eq_144_in1 = state_2_entry_BB_reg;
	// controller for eq_145.eq_145_in0
	// controller for eq_145.eq_145_in1
	// Insensitive connections
	assign eq_145_in0 = 32'd7;
	assign eq_145_in1 = state_2_entry_BB_reg;
	// controller for eq_195.eq_195_in0
	// controller for eq_195.eq_195_in1
	// Insensitive connections
	assign eq_195_in0 = 32'd0;
	assign eq_195_in1 = state_0_last_state;
	// controller for eq_196.eq_196_in0
	// controller for eq_196.eq_196_in1
	// Insensitive connections
	assign eq_196_in0 = 32'd3;
	assign eq_196_in1 = state_0_last_state;
	// controller for eq_200.eq_200_in0
	// controller for eq_200.eq_200_in1
	// Insensitive connections
	assign eq_200_in0 = 32'd0;
	assign eq_200_in1 = state_1_last_state;
	// controller for eq_201.eq_201_in0
	// controller for eq_201.eq_201_in1
	// Insensitive connections
	assign eq_201_in0 = 32'd1;
	assign eq_201_in1 = state_1_last_state;
	// controller for eq_202.eq_202_in0
	// controller for eq_202.eq_202_in1
	// Insensitive connections
	assign eq_202_in0 = 32'd1;
	assign eq_202_in1 = state_2_last_state;
	// controller for eq_203.eq_203_in0
	// controller for eq_203.eq_203_in1
	// Insensitive connections
	assign eq_203_in0 = 32'd2;
	assign eq_203_in1 = state_2_last_state;
	// controller for eq_206.eq_206_in0
	// controller for eq_206.eq_206_in1
	// Insensitive connections
	assign eq_206_in0 = 32'd2;
	assign eq_206_in1 = state_3_last_state;
	// controller for eq_207.eq_207_in0
	// controller for eq_207.eq_207_in1
	// Insensitive connections
	assign eq_207_in0 = 32'd3;
	assign eq_207_in1 = state_3_last_state;
	// controller for eq_208.eq_208_in0
	// controller for eq_208.eq_208_in1
	// Insensitive connections
	assign eq_208_in0 = 32'd3;
	assign eq_208_in1 = state_4_last_state;
	// controller for eq_209.eq_209_in0
	// controller for eq_209.eq_209_in1
	// Insensitive connections
	assign eq_209_in0 = 32'd4;
	assign eq_209_in1 = state_4_last_state;
	// controller for eq_210.eq_210_in0
	// controller for eq_210.eq_210_in1
	// Insensitive connections
	assign eq_210_in0 = 32'd4;
	assign eq_210_in1 = state_5_last_state;
	// controller for eq_211.eq_211_in0
	// controller for eq_211.eq_211_in1
	// Insensitive connections
	assign eq_211_in0 = 32'd5;
	assign eq_211_in1 = state_5_last_state;
	// controller for eq_75.eq_75_in0
	// controller for eq_75.eq_75_in1
	// Insensitive connections
	assign eq_75_in0 = 32'd3;
	assign eq_75_in1 = state_0_entry_BB_reg;
	// controller for eq_77.eq_77_in0
	// controller for eq_77.eq_77_in1
	// Insensitive connections
	assign eq_77_in0 = 32'd4;
	assign eq_77_in1 = state_0_entry_BB_reg;
	// controller for eq_79.eq_79_in0
	// controller for eq_79.eq_79_in1
	// Insensitive connections
	assign eq_79_in0 = 32'd5;
	assign eq_79_in1 = state_0_entry_BB_reg;
	// controller for eq_81.eq_81_in0
	// controller for eq_81.eq_81_in1
	// Insensitive connections
	assign eq_81_in0 = 32'd1;
	assign eq_81_in1 = state_0_entry_BB_reg;
	// controller for eq_83.eq_83_in0
	// controller for eq_83.eq_83_in1
	// Insensitive connections
	assign eq_83_in0 = 32'd0;
	assign eq_83_in1 = state_0_entry_BB_reg;
	// controller for eq_84.eq_84_in0
	// controller for eq_84.eq_84_in1
	// Insensitive connections
	assign eq_84_in0 = 32'd6;
	assign eq_84_in1 = state_1_entry_BB_reg;
	// controller for eq_85.eq_85_in0
	// controller for eq_85.eq_85_in1
	// Insensitive connections
	assign eq_85_in0 = 32'd6;
	assign eq_85_in1 = state_2_entry_BB_reg;
	// controller for eq_86.eq_86_in0
	// controller for eq_86.eq_86_in1
	// Insensitive connections
	assign eq_86_in0 = 32'd7;
	assign eq_86_in1 = state_2_entry_BB_reg;
	// controller for eq_88.eq_88_in0
	// controller for eq_88.eq_88_in1
	// Insensitive connections
	assign eq_88_in0 = 32'd8;
	assign eq_88_in1 = state_2_entry_BB_reg;
	// controller for eq_90.eq_90_in0
	// controller for eq_90.eq_90_in1
	// Insensitive connections
	assign eq_90_in0 = 32'd8;
	assign eq_90_in1 = state_3_entry_BB_reg;
	// controller for eq_91.eq_91_in0
	// controller for eq_91.eq_91_in1
	// Insensitive connections
	assign eq_91_in0 = 32'd2;
	assign eq_91_in1 = state_3_entry_BB_reg;
	// controller for eq_93.eq_93_in0
	// controller for eq_93.eq_93_in1
	// Insensitive connections
	assign eq_93_in0 = 32'd2;
	assign eq_93_in1 = state_4_entry_BB_reg;
	// controller for eq_94.eq_94_in0
	// controller for eq_94.eq_94_in1
	// Insensitive connections
	assign eq_94_in0 = 32'd2;
	assign eq_94_in1 = state_5_entry_BB_reg;
	// controller for eq_95.eq_95_in0
	// controller for eq_95.eq_95_in1
	// Insensitive connections
	assign eq_95_in0 = 32'd3;
	assign eq_95_in1 = state_0_entry_BB_reg;
	// controller for eq_98.eq_98_in0
	// controller for eq_98.eq_98_in1
	// Insensitive connections
	assign eq_98_in0 = 32'd4;
	assign eq_98_in1 = state_0_entry_BB_reg;
	// controller for icmp_icmp13.icmp_icmp13_in0
	// controller for icmp_icmp13.icmp_icmp13_in1
	// Insensitive connections
	assign icmp_icmp13_in0 = sext_sext0_out;
	assign icmp_icmp13_in1 = 32'd0;
	// controller for icmp_icmp28.icmp_icmp28_in0
	// controller for icmp_icmp28.icmp_icmp28_in1
	// Insensitive connections
	assign icmp_icmp28_in0 = sext_sext27_out;
	assign icmp_icmp28_in1 = 32'd0;
	// controller for icmp_icmp35.icmp_icmp35_in0
	// controller for icmp_icmp35.icmp_icmp35_in1
	// Insensitive connections
	assign icmp_icmp35_in0 = data_in_3_39_out_data;
	assign icmp_icmp35_in1 = data_in_3_37_out_data;
	// controller for icmp_icmp9.icmp_icmp9_in0
	// controller for icmp_icmp9.icmp_icmp9_in1
	// Insensitive connections
	assign icmp_icmp9_in0 = sext_sext8_out;
	assign icmp_icmp9_in1 = 32'd0;
	// controller for notOp_102.notOp_102_in0
	// Insensitive connections
	assign notOp_102_in0 = eq_101_out;
	// controller for notOp_105.notOp_105_in0
	// Insensitive connections
	assign notOp_105_in0 = eq_104_out;
	// controller for notOp_111.notOp_111_in0
	// Insensitive connections
	assign notOp_111_in0 = eq_110_out;
	// controller for notOp_114.notOp_114_in0
	// Insensitive connections
	assign notOp_114_in0 = eq_113_out;
	// controller for notOp_118.notOp_118_in0
	// Insensitive connections
	assign notOp_118_in0 = eq_117_out;
	// controller for notOp_175.notOp_175_in0
	// Insensitive connections
	assign notOp_175_in0 = andOp_42_out;
	// controller for notOp_177.notOp_177_in0
	// Insensitive connections
	assign notOp_177_in0 = andOp_49_out;
	// controller for notOp_179.notOp_179_in0
	// Insensitive connections
	assign notOp_179_in0 = andOp_67_out;
	// controller for notOp_181.notOp_181_in0
	// Insensitive connections
	assign notOp_181_in0 = andOp_51_out;
	// controller for notOp_183.notOp_183_in0
	// Insensitive connections
	assign notOp_183_in0 = andOp_170_out;
	// controller for notOp_185.notOp_185_in0
	// Insensitive connections
	assign notOp_185_in0 = andOp_62_out;
	// controller for notOp_187.notOp_187_in0
	// Insensitive connections
	assign notOp_187_in0 = andOp_171_out;
	// controller for notOp_189.notOp_189_in0
	// Insensitive connections
	assign notOp_189_in0 = andOp_172_out;
	// controller for notOp_191.notOp_191_in0
	// Insensitive connections
	assign notOp_191_in0 = andOp_173_out;
	// controller for notOp_193.notOp_193_in0
	// Insensitive connections
	assign notOp_193_in0 = andOp_174_out;
	// controller for notOp_41.notOp_41_in0
	// Insensitive connections
	assign notOp_41_in0 = andOp_40_out;
	// controller for notOp_43.notOp_43_in0
	// Insensitive connections
	assign notOp_43_in0 = icmp_icmp9_out;
	// controller for notOp_46.notOp_46_in0
	// Insensitive connections
	assign notOp_46_in0 = andOp_45_out;
	// controller for notOp_48.notOp_48_in0
	// Insensitive connections
	assign notOp_48_in0 = andOp_47_out;
	// controller for notOp_50.notOp_50_in0
	// Insensitive connections
	assign notOp_50_in0 = icmp_icmp13_out;
	// controller for notOp_53.notOp_53_in0
	// Insensitive connections
	assign notOp_53_in0 = andOp_52_out;
	// controller for notOp_55.notOp_55_in0
	// Insensitive connections
	assign notOp_55_in0 = andOp_54_out;
	// controller for notOp_57.notOp_57_in0
	// Insensitive connections
	assign notOp_57_in0 = andOp_56_out;
	// controller for notOp_59.notOp_59_in0
	// Insensitive connections
	assign notOp_59_in0 = andOp_58_out;
	// controller for notOp_61.notOp_61_in0
	// Insensitive connections
	assign notOp_61_in0 = andOp_60_out;
	// controller for notOp_63.notOp_63_in0
	// Insensitive connections
	assign notOp_63_in0 = icmp_icmp28_out;
	// controller for notOp_66.notOp_66_in0
	// Insensitive connections
	assign notOp_66_in0 = andOp_65_out;
	// controller for notOp_68.notOp_68_in0
	// Insensitive connections
	assign notOp_68_in0 = icmp_icmp35_out;
	// controller for notOp_71.notOp_71_in0
	// Insensitive connections
	assign notOp_71_in0 = andOp_70_out;
	// controller for notOp_73.notOp_73_in0
	// Insensitive connections
	assign notOp_73_in0 = icmp_icmp35_out;
	// controller for notOp_96.notOp_96_in0
	// Insensitive connections
	assign notOp_96_in0 = eq_95_out;
	// controller for notOp_99.notOp_99_in0
	// Insensitive connections
	assign notOp_99_in0 = eq_98_out;
	// controller for orOp_76.orOp_76_in0
	// controller for orOp_76.orOp_76_in1
	// Insensitive connections
	assign orOp_76_in0 = eq_75_out;
	assign orOp_76_in1 = andOp_54_out;
	// controller for orOp_78.orOp_78_in0
	// controller for orOp_78.orOp_78_in1
	// Insensitive connections
	assign orOp_78_in0 = eq_77_out;
	assign orOp_78_in1 = andOp_44_out;
	// controller for orOp_80.orOp_80_in0
	// controller for orOp_80.orOp_80_in1
	// Insensitive connections
	assign orOp_80_in0 = eq_79_out;
	assign orOp_80_in1 = andOp_52_out;
	// controller for orOp_82.orOp_82_in0
	// controller for orOp_82.orOp_82_in1
	// Insensitive connections
	assign orOp_82_in0 = eq_81_out;
	assign orOp_82_in1 = andOp_45_out;
	// controller for orOp_87.orOp_87_in0
	// controller for orOp_87.orOp_87_in1
	// Insensitive connections
	assign orOp_87_in0 = eq_86_out;
	assign orOp_87_in1 = andOp_56_out;
	// controller for orOp_89.orOp_89_in0
	// controller for orOp_89.orOp_89_in1
	// Insensitive connections
	assign orOp_89_in0 = eq_88_out;
	assign orOp_89_in1 = andOp_64_out;
	// controller for orOp_92.orOp_92_in0
	// controller for orOp_92.orOp_92_in1
	// Insensitive connections
	assign orOp_92_in0 = eq_91_out;
	assign orOp_92_in1 = andOp_69_out;
	// controller for phi_phi14.phi_phi14_in
	// controller for phi_phi14.phi_phi14_last_block
	// controller for phi_phi14.phi_phi14_s
	// Insensitive connections
	assign phi_phi14_in = concat_158_out;
	assign phi_phi14_last_block = bb_1_predecessor_in_state_0_out_data;
	assign phi_phi14_s = concat_159_out;
	// controller for ret40.valid_reg
	always @(*) begin
		if (andOp_169_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// controller for sext_sext0.sext_sext0_in
	// Insensitive connections
	assign sext_sext0_in = arg_0_read_ready;
	// controller for sext_sext27.sext_sext27_in
	// Insensitive connections
	assign sext_sext27_in = arg_3_s_axi_wready;
	// controller for sext_sext30.sext_sext30_in
	// Insensitive connections
	assign sext_sext30_in = data_in_2_21_out_data;
	// controller for sext_sext8.sext_sext8_in
	// Insensitive connections
	assign sext_sext8_in = arg_3_s_axi_awready;
	// controller for tmp_output_124.tmp_output_124_in_data
	always @(*) begin
		if (eq_125_out) begin 
			tmp_output_124_in_data = data_in_0_7_out_data;
		end else if (eq_128_out) begin 
			tmp_output_124_in_data = arg_1_rdata;
		end else begin
			tmp_output_124_in_data = 0;
		end
	end
	// controller for tmp_output_132.tmp_output_132_in_data
	always @(*) begin
		if (eq_133_out) begin 
			tmp_output_132_in_data = data_in_0_5_out_data;
		end else if (eq_136_out) begin 
			tmp_output_132_in_data = arg_2_rdata;
		end else begin
			tmp_output_132_in_data = 0;
		end
	end
	// controller for tmp_output_143.tmp_output_143_in_data
	always @(*) begin
		if (eq_144_out) begin 
			tmp_output_143_in_data = arg_0_out_data;
		end else if (eq_145_out) begin 
			tmp_output_143_in_data = data_in_2_23_out_data;
		end else begin
			tmp_output_143_in_data = 0;
		end
	end
	// controller for trunc_trunc32.trunc_trunc32_in
	// Insensitive connections
	assign trunc_trunc32_in = add_add31_out;
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			data_store_0_0 <= 0;
		end else begin
			if (andOp_197_out) begin
				data_store_0_0 <= phi_phi14_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_2 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_2 <= data_in_0_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_4 <= 0;
		end else begin
			if (andOp_198_out) begin
				data_store_0_4 <= arg_2_rdata;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_6 <= 0;
		end else begin
			if (andOp_199_out) begin
				data_store_0_6 <= arg_1_rdata;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_8 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_8 <= data_in_0_9_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_10 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_10 <= data_in_1_11_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_12 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_12 <= data_in_1_13_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_14 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_14 <= data_in_1_15_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_16 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_16 <= data_in_1_17_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_18 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_18 <= data_in_1_19_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_20 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_20 <= data_in_2_21_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_22 <= 0;
		end else begin
			if (andOp_204_out) begin
				data_store_2_22 <= arg_0_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_24 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_24 <= data_in_2_25_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_26 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_26 <= data_in_2_27_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_28 <= 0;
		end else begin
			if (andOp_205_out) begin
				data_store_2_28 <= trunc_trunc32_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_30 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_30 <= data_in_3_31_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_32 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_32 <= data_in_3_33_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_34 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_34 <= data_in_3_35_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_36 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_36 <= data_in_3_37_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_38 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_38 <= data_in_3_39_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_170_out) begin
				global_state <= 32'd2;
			end
			if (andOp_171_out) begin
				global_state <= 32'd3;
			end
			if (andOp_172_out) begin
				global_state <= 32'd4;
			end
			if (andOp_173_out) begin
				global_state <= 32'd5;
			end
			if (andOp_174_out) begin
				global_state <= 32'd5;
			end
			if (andOp_42_out) begin
				global_state <= 32'd0;
			end
			if (andOp_49_out) begin
				global_state <= 32'd0;
			end
			if (andOp_51_out) begin
				global_state <= 32'd1;
			end
			if (andOp_62_out) begin
				global_state <= 32'd2;
			end
			if (andOp_67_out) begin
				global_state <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
			if (andOp_42_out) begin
				state_0_entry_BB_reg <= 32'd3;
			end
			if (andOp_49_out) begin
				state_0_entry_BB_reg <= 32'd5;
			end
			if (andOp_67_out) begin
				state_0_entry_BB_reg <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (andOp_180_out) begin
				state_0_is_active <= 1'd0;
			end
			if (andOp_42_out) begin
				state_0_is_active <= 1'd1;
			end
			if (andOp_49_out) begin
				state_0_is_active <= 1'd1;
			end
			if (andOp_67_out) begin
				state_0_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
			if (andOp_42_out) begin
				state_0_last_BB_reg <= 32'd3;
			end
			if (andOp_49_out) begin
				state_0_last_BB_reg <= 32'd5;
			end
			if (andOp_67_out) begin
				state_0_last_BB_reg <= 32'd8;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
			if (andOp_42_out) begin
				state_0_last_state <= 32'd0;
			end
			if (andOp_49_out) begin
				state_0_last_state <= 32'd0;
			end
			if (andOp_67_out) begin
				state_0_last_state <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_51_out) begin
				state_1_entry_BB_reg <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_182_out) begin
				state_1_is_active <= 1'd0;
			end
			if (andOp_51_out) begin
				state_1_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_51_out) begin
				state_1_last_BB_reg <= 32'd5;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_51_out) begin
				state_1_last_state <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_170_out) begin
				state_2_entry_BB_reg <= 32'd6;
			end
			if (andOp_62_out) begin
				state_2_entry_BB_reg <= 32'd7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_170_out) begin
				state_2_is_active <= 1'd1;
			end
			if (andOp_186_out) begin
				state_2_is_active <= 1'd0;
			end
			if (andOp_62_out) begin
				state_2_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_170_out) begin
				state_2_last_BB_reg <= bb_6_predecessor_in_state_1_out_data;
			end
			if (andOp_62_out) begin
				state_2_last_BB_reg <= 32'd7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_170_out) begin
				state_2_last_state <= 32'd1;
			end
			if (andOp_62_out) begin
				state_2_last_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_171_out) begin
				state_3_entry_BB_reg <= 32'd8;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_171_out) begin
				state_3_is_active <= 1'd1;
			end
			if (andOp_188_out) begin
				state_3_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_171_out) begin
				state_3_last_BB_reg <= bb_8_predecessor_in_state_2_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_state <= 0;
		end else begin
			if (andOp_171_out) begin
				state_3_last_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_172_out) begin
				state_4_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_172_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_190_out) begin
				state_4_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_172_out) begin
				state_4_last_BB_reg <= bb_2_predecessor_in_state_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_state <= 0;
		end else begin
			if (andOp_172_out) begin
				state_4_last_state <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_entry_BB_reg <= 0;
		end else begin
			if (andOp_173_out) begin
				state_5_entry_BB_reg <= 32'd2;
			end
			if (andOp_174_out) begin
				state_5_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_is_active <= 0;
		end else begin
			if (andOp_173_out) begin
				state_5_is_active <= 1'd1;
			end
			if (andOp_174_out) begin
				state_5_is_active <= 1'd1;
			end
			if (andOp_194_out) begin
				state_5_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_last_BB_reg <= 0;
		end else begin
			if (andOp_173_out) begin
				state_5_last_BB_reg <= bb_2_predecessor_in_state_4_out_data;
			end
			if (andOp_174_out) begin
				state_5_last_BB_reg <= bb_2_predecessor_in_state_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_last_state <= 0;
		end else begin
			if (andOp_173_out) begin
				state_5_last_state <= 32'd4;
			end
			if (andOp_174_out) begin
				state_5_last_state <= 32'd5;
			end
		end
	end

endmodule

