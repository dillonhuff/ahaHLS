module mvmul(input [0:0] clk, input [0:0] rst, output [0:0] valid, output [4:0] ram_debug_addr, input [31:0] ram_debug_data, output [4:0] ram_debug_write_addr, output [31:0] ram_debug_write_data, output [0:0] ram_debug_write_en, output [4:0] ram_raddr_0, output [4:0] ram_raddr_1, output [4:0] ram_raddr_2, input [31:0] ram_rdata_0, input [31:0] ram_rdata_1, input [31:0] ram_rdata_2, output [0:0] ram_rst, output [4:0] ram_waddr_0, output [31:0] ram_wdata_0, output [0:0] ram_wen_0);

	reg [0:0] valid_reg;
	reg [4:0] ram_debug_addr_reg;
	reg [4:0] ram_debug_write_addr_reg;
	reg [31:0] ram_debug_write_data_reg;
	reg [0:0] ram_debug_write_en_reg;
	reg [4:0] ram_raddr_0_reg;
	reg [4:0] ram_raddr_1_reg;
	reg [4:0] ram_raddr_2_reg;
	reg [0:0] ram_rst_reg;
	reg [4:0] ram_waddr_0_reg;
	reg [31:0] ram_wdata_0_reg;
	reg [0:0] ram_wen_0_reg;

	assign valid = valid_reg;
	assign ram_debug_addr = ram_debug_addr_reg;
	assign ram_debug_write_addr = ram_debug_write_addr_reg;
	assign ram_debug_write_data = ram_debug_write_data_reg;
	assign ram_debug_write_en = ram_debug_write_en_reg;
	assign ram_raddr_0 = ram_raddr_0_reg;
	assign ram_raddr_1 = ram_raddr_1_reg;
	assign ram_raddr_2 = ram_raddr_2_reg;
	assign ram_rst = ram_rst_reg;
	assign ram_waddr_0 = ram_waddr_0_reg;
	assign ram_wdata_0 = ram_wdata_0_reg;
	assign ram_wen_0 = ram_wen_0_reg;

	// Start debug wires and ports

	initial begin
	end



	always @(posedge clk) begin
		if (!((!(andOp_192_out === 1) || andOp_99_out !== 1))) begin $display("assertion((!(andOp_192_out === 1) || andOp_99_out !== 1))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_99_out === 1) || andOp_192_out !== 1))) begin $display("assertion((!(andOp_99_out === 1) || andOp_192_out !== 1))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_196_out === 1) || andOp_197_out !== 1))) begin $display("assertion((!(andOp_196_out === 1) || andOp_197_out !== 1))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_197_out === 1) || andOp_196_out !== 1))) begin $display("assertion((!(andOp_197_out === 1) || andOp_196_out !== 1))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_192_out === 1) || andOp_99_out !== 1))) begin $display("assertion((!(andOp_192_out === 1) || andOp_99_out !== 1))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_99_out === 1) || andOp_192_out !== 1))) begin $display("assertion((!(andOp_99_out === 1) || andOp_192_out !== 1))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_196_out === 1) || andOp_197_out !== 1))) begin $display("assertion((!(andOp_196_out === 1) || andOp_197_out !== 1))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_197_out === 1) || andOp_196_out !== 1))) begin $display("assertion((!(andOp_197_out === 1) || andOp_196_out !== 1))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_119_out === 1) || andOp_199_out !== 1))) begin $display("assertion((!(andOp_119_out === 1) || andOp_199_out !== 1)) failed: Overlapping state active transition for state 0"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_199_out === 1) || andOp_119_out !== 1))) begin $display("assertion((!(andOp_199_out === 1) || andOp_119_out !== 1)) failed: Overlapping state active transition for state 0"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_190_out === 1) || andOp_201_out !== 1))) begin $display("assertion((!(andOp_190_out === 1) || andOp_201_out !== 1)) failed: Overlapping state active transition for state 1"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_201_out === 1) || andOp_190_out !== 1))) begin $display("assertion((!(andOp_201_out === 1) || andOp_190_out !== 1)) failed: Overlapping state active transition for state 1"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_191_out === 1) || andOp_203_out !== 1))) begin $display("assertion((!(andOp_191_out === 1) || andOp_203_out !== 1)) failed: Overlapping state active transition for state 2"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_203_out === 1) || andOp_191_out !== 1))) begin $display("assertion((!(andOp_203_out === 1) || andOp_191_out !== 1)) failed: Overlapping state active transition for state 2"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_192_out === 1) || andOp_207_out !== 1))) begin $display("assertion((!(andOp_192_out === 1) || andOp_207_out !== 1)) failed: Overlapping state active transition for state 3"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_192_out === 1) || andOp_99_out !== 1))) begin $display("assertion((!(andOp_192_out === 1) || andOp_99_out !== 1)) failed: Overlapping state active transition for state 3"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_207_out === 1) || andOp_192_out !== 1))) begin $display("assertion((!(andOp_207_out === 1) || andOp_192_out !== 1)) failed: Overlapping state active transition for state 3"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_207_out === 1) || andOp_99_out !== 1))) begin $display("assertion((!(andOp_207_out === 1) || andOp_99_out !== 1)) failed: Overlapping state active transition for state 3"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_99_out === 1) || andOp_192_out !== 1))) begin $display("assertion((!(andOp_99_out === 1) || andOp_192_out !== 1)) failed: Overlapping state active transition for state 3"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_99_out === 1) || andOp_207_out !== 1))) begin $display("assertion((!(andOp_99_out === 1) || andOp_207_out !== 1)) failed: Overlapping state active transition for state 3"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_193_out === 1) || andOp_209_out !== 1))) begin $display("assertion((!(andOp_193_out === 1) || andOp_209_out !== 1)) failed: Overlapping state active transition for state 4"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_209_out === 1) || andOp_193_out !== 1))) begin $display("assertion((!(andOp_209_out === 1) || andOp_193_out !== 1)) failed: Overlapping state active transition for state 4"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_194_out === 1) || andOp_211_out !== 1))) begin $display("assertion((!(andOp_194_out === 1) || andOp_211_out !== 1)) failed: Overlapping state active transition for state 5"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_211_out === 1) || andOp_194_out !== 1))) begin $display("assertion((!(andOp_211_out === 1) || andOp_194_out !== 1)) failed: Overlapping state active transition for state 5"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_195_out === 1) || andOp_213_out !== 1))) begin $display("assertion((!(andOp_195_out === 1) || andOp_213_out !== 1)) failed: Overlapping state active transition for state 6"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_213_out === 1) || andOp_195_out !== 1))) begin $display("assertion((!(andOp_213_out === 1) || andOp_195_out !== 1)) failed: Overlapping state active transition for state 6"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_196_out === 1) || andOp_197_out !== 1))) begin $display("assertion((!(andOp_196_out === 1) || andOp_197_out !== 1)) failed: Overlapping state active transition for state 7"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_196_out === 1) || andOp_217_out !== 1))) begin $display("assertion((!(andOp_196_out === 1) || andOp_217_out !== 1)) failed: Overlapping state active transition for state 7"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_197_out === 1) || andOp_196_out !== 1))) begin $display("assertion((!(andOp_197_out === 1) || andOp_196_out !== 1)) failed: Overlapping state active transition for state 7"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_197_out === 1) || andOp_217_out !== 1))) begin $display("assertion((!(andOp_197_out === 1) || andOp_217_out !== 1)) failed: Overlapping state active transition for state 7"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_217_out === 1) || andOp_196_out !== 1))) begin $display("assertion((!(andOp_217_out === 1) || andOp_196_out !== 1)) failed: Overlapping state active transition for state 7"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_217_out === 1) || andOp_197_out !== 1))) begin $display("assertion((!(andOp_217_out === 1) || andOp_197_out !== 1)) failed: Overlapping state active transition for state 7"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_168_out) || !(andOp_177_out)))) begin $display("assertion((!(andOp_168_out) || !(andOp_177_out)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_177_out) || !(andOp_168_out)))) begin $display("assertion((!(andOp_177_out) || !(andOp_168_out)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_1_is_active) || !(1'd0)))) begin $display("assertion((!(state_1_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_2_is_active) || !(1'd0)))) begin $display("assertion((!(state_2_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_3_is_active) || !(1'd0)))) begin $display("assertion((!(state_3_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_4_is_active) || !(1'd0)))) begin $display("assertion((!(state_4_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_5_is_active) || !(1'd0)))) begin $display("assertion((!(state_5_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_6_is_active) || !(1'd0)))) begin $display("assertion((!(state_6_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_7_is_active) || !(1'd0)))) begin $display("assertion((!(state_7_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_0_is_active) || !(1'd0)))) begin $display("assertion((!(state_0_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_1_is_active) || !(1'd0)))) begin $display("assertion((!(state_1_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_2_is_active) || !(1'd0)))) begin $display("assertion((!(state_2_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_3_is_active) || !(1'd0)))) begin $display("assertion((!(state_3_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_4_is_active) || !(1'd0)))) begin $display("assertion((!(state_4_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_5_is_active) || !(1'd0)))) begin $display("assertion((!(state_5_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_6_is_active) || !(1'd0)))) begin $display("assertion((!(state_6_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_4_is_active) || !(1'd0)))) begin $display("assertion((!(state_4_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_5_is_active) || !(1'd0)))) begin $display("assertion((!(state_5_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_6_is_active) || !(1'd0)))) begin $display("assertion((!(state_6_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_7_is_active) || !(1'd0)))) begin $display("assertion((!(state_7_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_0_is_active) || !(1'd0)))) begin $display("assertion((!(state_0_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_1_is_active) || !(1'd0)))) begin $display("assertion((!(state_1_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_2_is_active) || !(1'd0)))) begin $display("assertion((!(state_2_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_3_is_active) || !(1'd0)))) begin $display("assertion((!(state_3_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_4_is_active) || !(1'd0)))) begin $display("assertion((!(state_4_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_5_is_active) || !(1'd0)))) begin $display("assertion((!(state_5_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_6_is_active) || !(1'd0)))) begin $display("assertion((!(state_6_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_0_is_active) || !(1'd0)))) begin $display("assertion((!(state_0_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_1_is_active) || !(1'd0)))) begin $display("assertion((!(state_1_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_2_is_active) || !(1'd0)))) begin $display("assertion((!(state_2_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_241_out) || add_add2_in0 !== 32'dx)) begin $display("assertion(!(andOp_241_out) || add_add2_in0 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_241_out) || add_add2_in1 !== 32'dx)) begin $display("assertion(!(andOp_241_out) || add_add2_in1 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_242_out) || add_add9_in0 !== 32'dx)) begin $display("assertion(!(andOp_242_out) || add_add9_in0 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_242_out) || add_add9_in1 !== 32'dx)) begin $display("assertion(!(andOp_242_out) || add_add9_in1 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_243_out) || add_add10_in0 !== 32'dx)) begin $display("assertion(!(andOp_243_out) || add_add10_in0 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_243_out) || add_add10_in1 !== 32'dx)) begin $display("assertion(!(andOp_243_out) || add_add10_in1 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_244_out) || add_add11_in0 !== 32'dx)) begin $display("assertion(!(andOp_244_out) || add_add11_in0 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_244_out) || add_add11_in1 !== 32'dx)) begin $display("assertion(!(andOp_244_out) || add_add11_in1 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_245_out) || add_add17_in0 !== 32'dx)) begin $display("assertion(!(andOp_245_out) || add_add17_in0 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_245_out) || add_add17_in1 !== 32'dx)) begin $display("assertion(!(andOp_245_out) || add_add17_in1 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_246_out) || add_add25_in0 !== 32'dx)) begin $display("assertion(!(andOp_246_out) || add_add25_in0 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_246_out) || add_add25_in1 !== 32'dx)) begin $display("assertion(!(andOp_246_out) || add_add25_in1 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_247_out) || mul_mul3_in0 !== 32'dx)) begin $display("assertion(!(andOp_247_out) || mul_mul3_in0 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_247_out) || mul_mul3_in1 !== 32'dx)) begin $display("assertion(!(andOp_247_out) || mul_mul3_in1 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_248_out) || mul_mul16_in0 !== 32'dx)) begin $display("assertion(!(andOp_248_out) || mul_mul16_in0 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_248_out) || mul_mul16_in1 !== 32'dx)) begin $display("assertion(!(andOp_248_out) || mul_mul16_in1 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_249_out) || phi_phi1_out !== 'dx))) begin $display("assertion((!(andOp_249_out) || phi_phi1_out !== 'dx))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_250_out) || phi_phi7_out !== 'dx))) begin $display("assertion((!(andOp_250_out) || phi_phi7_out !== 'dx))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_251_out) || add_add2_out !== 32'dx))) begin $display("assertion((!(andOp_251_out) || add_add2_out !== 32'dx))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_252_out) || data_in_4_41_out_data !== 32'dx))) begin $display("assertion((!(andOp_252_out) || data_in_4_41_out_data !== 32'dx))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_253_out) || 32'd0 !== 32'dx))) begin $display("assertion((!(andOp_253_out) || 32'd0 !== 32'dx))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_254_out) || add_add17_out !== 32'dx))) begin $display("assertion((!(andOp_254_out) || add_add17_out !== 32'dx))"); $finish(); end
	end




	// End debug wires and ports

	// Start Functional Units
	br_dummy br_unit();

	wire [63:0] phi_phi7_in;
	wire [31:0] phi_phi7_last_block;
	wire [63:0] phi_phi7_s;
	wire [31:0] phi_phi7_out;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_phi7(.in(phi_phi7_in), .last_block(phi_phi7_last_block), .out(phi_phi7_out), .s(phi_phi7_s));

	wire [63:0] phi_phi1_in;
	wire [31:0] phi_phi1_last_block;
	wire [63:0] phi_phi1_s;
	wire [31:0] phi_phi1_out;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_phi1(.in(phi_phi1_in), .last_block(phi_phi1_last_block), .out(phi_phi1_out), .s(phi_phi1_s));

	wire [31:0] add_add2_in0;
	wire [31:0] add_add2_in1;
	wire [31:0] add_add2_out;
	add #(.WIDTH(32)) add_add2(.in0(add_add2_in0), .in1(add_add2_in1), .out(add_add2_out));

	wire [31:0] mul_mul3_in0;
	wire [31:0] mul_mul3_in1;
	wire [31:0] mul_mul3_out;
	mul #(.WIDTH(32)) mul_mul3(.in0(mul_mul3_in0), .in1(mul_mul3_in1), .out(mul_mul3_out));

	wire [31:0] add_add25_in0;
	wire [31:0] add_add25_in1;
	wire [31:0] add_add25_out;
	add #(.WIDTH(32)) add_add25(.in0(add_add25_in0), .in1(add_add25_in1), .out(add_add25_out));

	wire [31:0] icmp_icmp26_in0;
	wire [31:0] icmp_icmp26_in1;
	wire [0:0] icmp_icmp26_out;
	eq #(.WIDTH(32)) icmp_icmp26(.in0(icmp_icmp26_in0), .in1(icmp_icmp26_in1), .out(icmp_icmp26_out));

	wire [31:0] add_add9_in0;
	wire [31:0] add_add9_in1;
	wire [31:0] add_add9_out;
	add #(.WIDTH(32)) add_add9(.in0(add_add9_in0), .in1(add_add9_in1), .out(add_add9_out));

	wire [31:0] add_add10_in0;
	wire [31:0] add_add10_in1;
	wire [31:0] add_add10_out;
	add #(.WIDTH(32)) add_add10(.in0(add_add10_in0), .in1(add_add10_in1), .out(add_add10_out));

	wire [31:0] mul_mul16_in0;
	wire [31:0] mul_mul16_in1;
	wire [31:0] mul_mul16_out;
	mul #(.WIDTH(32)) mul_mul16(.in0(mul_mul16_in0), .in1(mul_mul16_in1), .out(mul_mul16_out));

	wire [31:0] add_add17_in0;
	wire [31:0] add_add17_in1;
	wire [31:0] add_add17_out;
	add #(.WIDTH(32)) add_add17(.in0(add_add17_in0), .in1(add_add17_in1), .out(add_add17_out));

	wire [31:0] add_add11_in0;
	wire [31:0] add_add11_in1;
	wire [31:0] add_add11_out;
	add #(.WIDTH(32)) add_add11(.in0(add_add11_in0), .in1(add_add11_in1), .out(add_add11_out));

	wire [31:0] icmp_icmp12_in0;
	wire [31:0] icmp_icmp12_in1;
	wire [0:0] icmp_icmp12_out;
	eq #(.WIDTH(32)) icmp_icmp12(.in0(icmp_icmp12_in0), .in1(icmp_icmp12_in1), .out(icmp_icmp12_out));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] bb_2_active_in_state_0_in_data;
	wire [0:0] bb_2_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_0(.in_data(bb_2_active_in_state_0_in_data), .out_data(bb_2_active_in_state_0_out_data));

	reg [31:0] bb_2_predecessor_in_state_0_in_data;
	wire [31:0] bb_2_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_0(.in_data(bb_2_predecessor_in_state_0_in_data), .out_data(bb_2_predecessor_in_state_0_out_data));

	reg [0:0] br_2_happened_in_state_0_in_data;
	wire [0:0] br_2_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_2_happened_in_state_0(.in_data(br_2_happened_in_state_0_in_data), .out_data(br_2_happened_in_state_0_out_data));

	reg [0:0] bb_2_active_in_state_1_in_data;
	wire [0:0] bb_2_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_1(.in_data(bb_2_active_in_state_1_in_data), .out_data(bb_2_active_in_state_1_out_data));

	reg [31:0] bb_2_predecessor_in_state_1_in_data;
	wire [31:0] bb_2_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_1(.in_data(bb_2_predecessor_in_state_1_in_data), .out_data(bb_2_predecessor_in_state_1_out_data));

	reg [0:0] br_2_happened_in_state_1_in_data;
	wire [0:0] br_2_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_2_happened_in_state_1(.in_data(br_2_happened_in_state_1_in_data), .out_data(br_2_happened_in_state_1_out_data));

	reg [0:0] bb_2_active_in_state_2_in_data;
	wire [0:0] bb_2_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_2(.in_data(bb_2_active_in_state_2_in_data), .out_data(bb_2_active_in_state_2_out_data));

	reg [31:0] bb_2_predecessor_in_state_2_in_data;
	wire [31:0] bb_2_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_2(.in_data(bb_2_predecessor_in_state_2_in_data), .out_data(bb_2_predecessor_in_state_2_out_data));

	reg [0:0] br_2_happened_in_state_2_in_data;
	wire [0:0] br_2_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_2_happened_in_state_2(.in_data(br_2_happened_in_state_2_in_data), .out_data(br_2_happened_in_state_2_out_data));

	reg [0:0] bb_2_active_in_state_3_in_data;
	wire [0:0] bb_2_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_3(.in_data(bb_2_active_in_state_3_in_data), .out_data(bb_2_active_in_state_3_out_data));

	reg [31:0] bb_2_predecessor_in_state_3_in_data;
	wire [31:0] bb_2_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_3(.in_data(bb_2_predecessor_in_state_3_in_data), .out_data(bb_2_predecessor_in_state_3_out_data));

	reg [0:0] br_2_happened_in_state_3_in_data;
	wire [0:0] br_2_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_2_happened_in_state_3(.in_data(br_2_happened_in_state_3_in_data), .out_data(br_2_happened_in_state_3_out_data));

	reg [0:0] bb_4_active_in_state_3_in_data;
	wire [0:0] bb_4_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_3(.in_data(bb_4_active_in_state_3_in_data), .out_data(bb_4_active_in_state_3_out_data));

	reg [31:0] bb_4_predecessor_in_state_3_in_data;
	wire [31:0] bb_4_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_3(.in_data(bb_4_predecessor_in_state_3_in_data), .out_data(bb_4_predecessor_in_state_3_out_data));

	reg [0:0] br_4_happened_in_state_3_in_data;
	wire [0:0] br_4_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_3(.in_data(br_4_happened_in_state_3_in_data), .out_data(br_4_happened_in_state_3_out_data));

	reg [0:0] bb_4_active_in_state_4_in_data;
	wire [0:0] bb_4_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_4(.in_data(bb_4_active_in_state_4_in_data), .out_data(bb_4_active_in_state_4_out_data));

	reg [31:0] bb_4_predecessor_in_state_4_in_data;
	wire [31:0] bb_4_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_4(.in_data(bb_4_predecessor_in_state_4_in_data), .out_data(bb_4_predecessor_in_state_4_out_data));

	reg [0:0] br_4_happened_in_state_4_in_data;
	wire [0:0] br_4_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_4(.in_data(br_4_happened_in_state_4_in_data), .out_data(br_4_happened_in_state_4_out_data));

	reg [0:0] bb_4_active_in_state_5_in_data;
	wire [0:0] bb_4_active_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_5(.in_data(bb_4_active_in_state_5_in_data), .out_data(bb_4_active_in_state_5_out_data));

	reg [31:0] bb_4_predecessor_in_state_5_in_data;
	wire [31:0] bb_4_predecessor_in_state_5_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_5(.in_data(bb_4_predecessor_in_state_5_in_data), .out_data(bb_4_predecessor_in_state_5_out_data));

	reg [0:0] br_4_happened_in_state_5_in_data;
	wire [0:0] br_4_happened_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_5(.in_data(br_4_happened_in_state_5_in_data), .out_data(br_4_happened_in_state_5_out_data));

	reg [0:0] bb_4_active_in_state_6_in_data;
	wire [0:0] bb_4_active_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_6(.in_data(bb_4_active_in_state_6_in_data), .out_data(bb_4_active_in_state_6_out_data));

	reg [31:0] bb_4_predecessor_in_state_6_in_data;
	wire [31:0] bb_4_predecessor_in_state_6_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_6(.in_data(bb_4_predecessor_in_state_6_in_data), .out_data(bb_4_predecessor_in_state_6_out_data));

	reg [0:0] br_4_happened_in_state_6_in_data;
	wire [0:0] br_4_happened_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_6(.in_data(br_4_happened_in_state_6_in_data), .out_data(br_4_happened_in_state_6_out_data));

	reg [0:0] bb_1_active_in_state_7_in_data;
	wire [0:0] bb_1_active_in_state_7_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_7(.in_data(bb_1_active_in_state_7_in_data), .out_data(bb_1_active_in_state_7_out_data));

	reg [31:0] bb_1_predecessor_in_state_7_in_data;
	wire [31:0] bb_1_predecessor_in_state_7_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_7(.in_data(bb_1_predecessor_in_state_7_in_data), .out_data(bb_1_predecessor_in_state_7_out_data));

	reg [0:0] bb_3_active_in_state_7_in_data;
	wire [0:0] bb_3_active_in_state_7_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_7(.in_data(bb_3_active_in_state_7_in_data), .out_data(bb_3_active_in_state_7_out_data));

	reg [31:0] bb_3_predecessor_in_state_7_in_data;
	wire [31:0] bb_3_predecessor_in_state_7_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_7(.in_data(bb_3_predecessor_in_state_7_in_data), .out_data(bb_3_predecessor_in_state_7_out_data));

	reg [0:0] br_3_happened_in_state_7_in_data;
	wire [0:0] br_3_happened_in_state_7_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_7(.in_data(br_3_happened_in_state_7_in_data), .out_data(br_3_happened_in_state_7_out_data));

	reg [0:0] bb_4_active_in_state_7_in_data;
	wire [0:0] bb_4_active_in_state_7_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_7(.in_data(bb_4_active_in_state_7_in_data), .out_data(bb_4_active_in_state_7_out_data));

	reg [31:0] bb_4_predecessor_in_state_7_in_data;
	wire [31:0] bb_4_predecessor_in_state_7_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_7(.in_data(bb_4_predecessor_in_state_7_in_data), .out_data(bb_4_predecessor_in_state_7_out_data));

	reg [0:0] br_4_happened_in_state_7_in_data;
	wire [0:0] br_4_happened_in_state_7_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_7(.in_data(br_4_happened_in_state_7_in_data), .out_data(br_4_happened_in_state_7_out_data));

	reg [31:0] data_in_0_4_in_data;
	wire [31:0] data_in_0_4_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_4(.in_data(data_in_0_4_in_data), .out_data(data_in_0_4_out_data));

	reg [31:0] data_in_0_6_in_data;
	wire [31:0] data_in_0_6_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_6(.in_data(data_in_0_6_in_data), .out_data(data_in_0_6_out_data));

	reg [31:0] data_in_1_8_in_data;
	wire [31:0] data_in_1_8_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_8(.in_data(data_in_1_8_in_data), .out_data(data_in_1_8_out_data));

	reg [31:0] data_in_1_10_in_data;
	wire [31:0] data_in_1_10_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_10(.in_data(data_in_1_10_in_data), .out_data(data_in_1_10_out_data));

	reg [31:0] data_in_1_12_in_data;
	wire [31:0] data_in_1_12_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_12(.in_data(data_in_1_12_in_data), .out_data(data_in_1_12_out_data));

	reg [31:0] data_in_1_14_in_data;
	wire [31:0] data_in_1_14_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_14(.in_data(data_in_1_14_in_data), .out_data(data_in_1_14_out_data));

	reg [31:0] data_in_1_16_in_data;
	wire [31:0] data_in_1_16_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_16(.in_data(data_in_1_16_in_data), .out_data(data_in_1_16_out_data));

	reg [31:0] data_in_2_18_in_data;
	wire [31:0] data_in_2_18_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_18(.in_data(data_in_2_18_in_data), .out_data(data_in_2_18_out_data));

	reg [31:0] data_in_2_20_in_data;
	wire [31:0] data_in_2_20_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_20(.in_data(data_in_2_20_in_data), .out_data(data_in_2_20_out_data));

	reg [31:0] data_in_2_22_in_data;
	wire [31:0] data_in_2_22_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_22(.in_data(data_in_2_22_in_data), .out_data(data_in_2_22_out_data));

	reg [31:0] data_in_2_24_in_data;
	wire [31:0] data_in_2_24_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_24(.in_data(data_in_2_24_in_data), .out_data(data_in_2_24_out_data));

	reg [31:0] data_in_2_26_in_data;
	wire [31:0] data_in_2_26_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_26(.in_data(data_in_2_26_in_data), .out_data(data_in_2_26_out_data));

	reg [31:0] data_in_3_28_in_data;
	wire [31:0] data_in_3_28_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_28(.in_data(data_in_3_28_in_data), .out_data(data_in_3_28_out_data));

	reg [31:0] data_in_3_30_in_data;
	wire [31:0] data_in_3_30_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_30(.in_data(data_in_3_30_in_data), .out_data(data_in_3_30_out_data));

	reg [31:0] data_in_3_32_in_data;
	wire [31:0] data_in_3_32_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_32(.in_data(data_in_3_32_in_data), .out_data(data_in_3_32_out_data));

	reg [31:0] data_in_3_34_in_data;
	wire [31:0] data_in_3_34_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_34(.in_data(data_in_3_34_in_data), .out_data(data_in_3_34_out_data));

	reg [31:0] data_in_3_36_in_data;
	wire [31:0] data_in_3_36_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_36(.in_data(data_in_3_36_in_data), .out_data(data_in_3_36_out_data));

	reg [31:0] data_in_4_39_in_data;
	wire [31:0] data_in_4_39_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_39(.in_data(data_in_4_39_in_data), .out_data(data_in_4_39_out_data));

	reg [31:0] data_in_4_41_in_data;
	wire [31:0] data_in_4_41_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_41(.in_data(data_in_4_41_in_data), .out_data(data_in_4_41_out_data));

	reg [31:0] data_in_4_43_in_data;
	wire [31:0] data_in_4_43_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_43(.in_data(data_in_4_43_in_data), .out_data(data_in_4_43_out_data));

	reg [31:0] data_in_4_45_in_data;
	wire [31:0] data_in_4_45_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_45(.in_data(data_in_4_45_in_data), .out_data(data_in_4_45_out_data));

	reg [31:0] data_in_4_47_in_data;
	wire [31:0] data_in_4_47_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_47(.in_data(data_in_4_47_in_data), .out_data(data_in_4_47_out_data));

	reg [0:0] data_in_4_49_in_data;
	wire [0:0] data_in_4_49_out_data;
	hls_wire #(.WIDTH(1)) data_in_4_49(.in_data(data_in_4_49_in_data), .out_data(data_in_4_49_out_data));

	reg [31:0] data_in_5_51_in_data;
	wire [31:0] data_in_5_51_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_51(.in_data(data_in_5_51_in_data), .out_data(data_in_5_51_out_data));

	reg [31:0] data_in_5_53_in_data;
	wire [31:0] data_in_5_53_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_53(.in_data(data_in_5_53_in_data), .out_data(data_in_5_53_out_data));

	reg [31:0] data_in_5_55_in_data;
	wire [31:0] data_in_5_55_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_55(.in_data(data_in_5_55_in_data), .out_data(data_in_5_55_out_data));

	reg [31:0] data_in_5_57_in_data;
	wire [31:0] data_in_5_57_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_57(.in_data(data_in_5_57_in_data), .out_data(data_in_5_57_out_data));

	reg [31:0] data_in_5_59_in_data;
	wire [31:0] data_in_5_59_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_59(.in_data(data_in_5_59_in_data), .out_data(data_in_5_59_out_data));

	reg [0:0] data_in_5_61_in_data;
	wire [0:0] data_in_5_61_out_data;
	hls_wire #(.WIDTH(1)) data_in_5_61(.in_data(data_in_5_61_in_data), .out_data(data_in_5_61_out_data));

	reg [31:0] data_in_6_63_in_data;
	wire [31:0] data_in_6_63_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_63(.in_data(data_in_6_63_in_data), .out_data(data_in_6_63_out_data));

	reg [31:0] data_in_6_65_in_data;
	wire [31:0] data_in_6_65_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_65(.in_data(data_in_6_65_in_data), .out_data(data_in_6_65_out_data));

	reg [31:0] data_in_6_67_in_data;
	wire [31:0] data_in_6_67_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_67(.in_data(data_in_6_67_in_data), .out_data(data_in_6_67_out_data));

	reg [31:0] data_in_6_69_in_data;
	wire [31:0] data_in_6_69_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_69(.in_data(data_in_6_69_in_data), .out_data(data_in_6_69_out_data));

	reg [31:0] data_in_6_71_in_data;
	wire [31:0] data_in_6_71_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_71(.in_data(data_in_6_71_in_data), .out_data(data_in_6_71_out_data));

	reg [0:0] data_in_6_73_in_data;
	wire [0:0] data_in_6_73_out_data;
	hls_wire #(.WIDTH(1)) data_in_6_73(.in_data(data_in_6_73_in_data), .out_data(data_in_6_73_out_data));

	reg [31:0] data_in_7_75_in_data;
	wire [31:0] data_in_7_75_out_data;
	hls_wire #(.WIDTH(32)) data_in_7_75(.in_data(data_in_7_75_in_data), .out_data(data_in_7_75_out_data));

	reg [31:0] data_in_7_77_in_data;
	wire [31:0] data_in_7_77_out_data;
	hls_wire #(.WIDTH(32)) data_in_7_77(.in_data(data_in_7_77_in_data), .out_data(data_in_7_77_out_data));

	reg [31:0] data_in_7_79_in_data;
	wire [31:0] data_in_7_79_out_data;
	hls_wire #(.WIDTH(32)) data_in_7_79(.in_data(data_in_7_79_in_data), .out_data(data_in_7_79_out_data));

	reg [31:0] data_in_7_81_in_data;
	wire [31:0] data_in_7_81_out_data;
	hls_wire #(.WIDTH(32)) data_in_7_81(.in_data(data_in_7_81_in_data), .out_data(data_in_7_81_out_data));

	reg [31:0] data_in_7_83_in_data;
	wire [31:0] data_in_7_83_out_data;
	hls_wire #(.WIDTH(32)) data_in_7_83(.in_data(data_in_7_83_in_data), .out_data(data_in_7_83_out_data));

	reg [0:0] data_in_7_84_in_data;
	wire [0:0] data_in_7_84_out_data;
	hls_wire #(.WIDTH(1)) data_in_7_84(.in_data(data_in_7_84_in_data), .out_data(data_in_7_84_out_data));

	wire [0:0] andOp_85_in0;
	wire [0:0] andOp_85_in1;
	wire [0:0] andOp_85_out;
	andOp #(.WIDTH(1)) andOp_85(.in0(andOp_85_in0), .in1(andOp_85_in1), .out(andOp_85_out));

	wire [0:0] notOp_86_in0;
	wire [0:0] notOp_86_out;
	notOp #(.WIDTH(1)) notOp_86(.in(notOp_86_in0), .out(notOp_86_out));

	wire [0:0] andOp_87_in0;
	wire [0:0] andOp_87_in1;
	wire [0:0] andOp_87_out;
	andOp #(.WIDTH(1)) andOp_87(.in0(andOp_87_in0), .in1(andOp_87_in1), .out(andOp_87_out));

	wire [0:0] notOp_88_in0;
	wire [0:0] notOp_88_out;
	notOp #(.WIDTH(1)) notOp_88(.in(notOp_88_in0), .out(notOp_88_out));

	wire [0:0] andOp_89_in0;
	wire [0:0] andOp_89_in1;
	wire [0:0] andOp_89_out;
	andOp #(.WIDTH(1)) andOp_89(.in0(andOp_89_in0), .in1(andOp_89_in1), .out(andOp_89_out));

	wire [0:0] notOp_90_in0;
	wire [0:0] notOp_90_out;
	notOp #(.WIDTH(1)) notOp_90(.in(notOp_90_in0), .out(notOp_90_out));

	wire [0:0] andOp_91_in0;
	wire [0:0] andOp_91_in1;
	wire [0:0] andOp_91_out;
	andOp #(.WIDTH(1)) andOp_91(.in0(andOp_91_in0), .in1(andOp_91_in1), .out(andOp_91_out));

	wire [0:0] notOp_92_in0;
	wire [0:0] notOp_92_out;
	notOp #(.WIDTH(1)) notOp_92(.in(notOp_92_in0), .out(notOp_92_out));

	wire [0:0] andOp_93_in0;
	wire [0:0] andOp_93_in1;
	wire [0:0] andOp_93_out;
	andOp #(.WIDTH(1)) andOp_93(.in0(andOp_93_in0), .in1(andOp_93_in1), .out(andOp_93_out));

	wire [0:0] notOp_94_in0;
	wire [0:0] notOp_94_out;
	notOp #(.WIDTH(1)) notOp_94(.in(notOp_94_in0), .out(notOp_94_out));

	wire [0:0] andOp_95_in0;
	wire [0:0] andOp_95_in1;
	wire [0:0] andOp_95_out;
	andOp #(.WIDTH(1)) andOp_95(.in0(andOp_95_in0), .in1(andOp_95_in1), .out(andOp_95_out));

	wire [0:0] notOp_96_in0;
	wire [0:0] notOp_96_out;
	notOp #(.WIDTH(1)) notOp_96(.in(notOp_96_in0), .out(notOp_96_out));

	wire [0:0] andOp_97_in0;
	wire [0:0] andOp_97_in1;
	wire [0:0] andOp_97_out;
	andOp #(.WIDTH(1)) andOp_97(.in0(andOp_97_in0), .in1(andOp_97_in1), .out(andOp_97_out));

	wire [0:0] notOp_98_in0;
	wire [0:0] notOp_98_out;
	notOp #(.WIDTH(1)) notOp_98(.in(notOp_98_in0), .out(notOp_98_out));

	wire [0:0] andOp_99_in0;
	wire [0:0] andOp_99_in1;
	wire [0:0] andOp_99_out;
	andOp #(.WIDTH(1)) andOp_99(.in0(andOp_99_in0), .in1(andOp_99_in1), .out(andOp_99_out));

	wire [0:0] andOp_100_in0;
	wire [0:0] andOp_100_in1;
	wire [0:0] andOp_100_out;
	andOp #(.WIDTH(1)) andOp_100(.in0(andOp_100_in0), .in1(andOp_100_in1), .out(andOp_100_out));

	wire [0:0] notOp_101_in0;
	wire [0:0] notOp_101_out;
	notOp #(.WIDTH(1)) notOp_101(.in(notOp_101_in0), .out(notOp_101_out));

	wire [0:0] andOp_102_in0;
	wire [0:0] andOp_102_in1;
	wire [0:0] andOp_102_out;
	andOp #(.WIDTH(1)) andOp_102(.in0(andOp_102_in0), .in1(andOp_102_in1), .out(andOp_102_out));

	wire [0:0] notOp_103_in0;
	wire [0:0] notOp_103_out;
	notOp #(.WIDTH(1)) notOp_103(.in(notOp_103_in0), .out(notOp_103_out));

	wire [0:0] andOp_104_in0;
	wire [0:0] andOp_104_in1;
	wire [0:0] andOp_104_out;
	andOp #(.WIDTH(1)) andOp_104(.in0(andOp_104_in0), .in1(andOp_104_in1), .out(andOp_104_out));

	wire [0:0] andOp_105_in0;
	wire [0:0] andOp_105_in1;
	wire [0:0] andOp_105_out;
	andOp #(.WIDTH(1)) andOp_105(.in0(andOp_105_in0), .in1(andOp_105_in1), .out(andOp_105_out));

	wire [0:0] notOp_106_in0;
	wire [0:0] notOp_106_out;
	notOp #(.WIDTH(1)) notOp_106(.in(notOp_106_in0), .out(notOp_106_out));

	wire [0:0] andOp_107_in0;
	wire [0:0] andOp_107_in1;
	wire [0:0] andOp_107_out;
	andOp #(.WIDTH(1)) andOp_107(.in0(andOp_107_in0), .in1(andOp_107_in1), .out(andOp_107_out));

	wire [0:0] notOp_108_in0;
	wire [0:0] notOp_108_out;
	notOp #(.WIDTH(1)) notOp_108(.in(notOp_108_in0), .out(notOp_108_out));

	wire [0:0] andOp_109_in0;
	wire [0:0] andOp_109_in1;
	wire [0:0] andOp_109_out;
	andOp #(.WIDTH(1)) andOp_109(.in0(andOp_109_in0), .in1(andOp_109_in1), .out(andOp_109_out));

	wire [0:0] andOp_110_in0;
	wire [0:0] andOp_110_in1;
	wire [0:0] andOp_110_out;
	andOp #(.WIDTH(1)) andOp_110(.in0(andOp_110_in0), .in1(andOp_110_in1), .out(andOp_110_out));

	wire [0:0] notOp_111_in0;
	wire [0:0] notOp_111_out;
	notOp #(.WIDTH(1)) notOp_111(.in(notOp_111_in0), .out(notOp_111_out));

	wire [0:0] andOp_112_in0;
	wire [0:0] andOp_112_in1;
	wire [0:0] andOp_112_out;
	andOp #(.WIDTH(1)) andOp_112(.in0(andOp_112_in0), .in1(andOp_112_in1), .out(andOp_112_out));

	wire [0:0] notOp_113_in0;
	wire [0:0] notOp_113_out;
	notOp #(.WIDTH(1)) notOp_113(.in(notOp_113_in0), .out(notOp_113_out));

	wire [0:0] andOp_114_in0;
	wire [0:0] andOp_114_in1;
	wire [0:0] andOp_114_out;
	andOp #(.WIDTH(1)) andOp_114(.in0(andOp_114_in0), .in1(andOp_114_in1), .out(andOp_114_out));

	wire [0:0] andOp_115_in0;
	wire [0:0] andOp_115_in1;
	wire [0:0] andOp_115_out;
	andOp #(.WIDTH(1)) andOp_115(.in0(andOp_115_in0), .in1(andOp_115_in1), .out(andOp_115_out));

	wire [0:0] notOp_116_in0;
	wire [0:0] notOp_116_out;
	notOp #(.WIDTH(1)) notOp_116(.in(notOp_116_in0), .out(notOp_116_out));

	wire [0:0] andOp_117_in0;
	wire [0:0] andOp_117_in1;
	wire [0:0] andOp_117_out;
	andOp #(.WIDTH(1)) andOp_117(.in0(andOp_117_in0), .in1(andOp_117_in1), .out(andOp_117_out));

	wire [0:0] notOp_118_in0;
	wire [0:0] notOp_118_out;
	notOp #(.WIDTH(1)) notOp_118(.in(notOp_118_in0), .out(notOp_118_out));

	wire [0:0] andOp_119_in0;
	wire [0:0] andOp_119_in1;
	wire [0:0] andOp_119_out;
	andOp #(.WIDTH(1)) andOp_119(.in0(andOp_119_in0), .in1(andOp_119_in1), .out(andOp_119_out));

	wire [0:0] andOp_120_in0;
	wire [0:0] andOp_120_in1;
	wire [0:0] andOp_120_out;
	andOp #(.WIDTH(1)) andOp_120(.in0(andOp_120_in0), .in1(andOp_120_in1), .out(andOp_120_out));

	wire [0:0] notOp_121_in0;
	wire [0:0] notOp_121_out;
	notOp #(.WIDTH(1)) notOp_121(.in(notOp_121_in0), .out(notOp_121_out));

	wire [0:0] andOp_122_in0;
	wire [0:0] andOp_122_in1;
	wire [0:0] andOp_122_out;
	andOp #(.WIDTH(1)) andOp_122(.in0(andOp_122_in0), .in1(andOp_122_in1), .out(andOp_122_out));

	wire [0:0] notOp_123_in0;
	wire [0:0] notOp_123_out;
	notOp #(.WIDTH(1)) notOp_123(.in(notOp_123_in0), .out(notOp_123_out));

	wire [0:0] andOp_124_in0;
	wire [0:0] andOp_124_in1;
	wire [0:0] andOp_124_out;
	andOp #(.WIDTH(1)) andOp_124(.in0(andOp_124_in0), .in1(andOp_124_in1), .out(andOp_124_out));

	wire [31:0] eq_125_in0;
	wire [31:0] eq_125_in1;
	wire [0:0] eq_125_out;
	eq #(.WIDTH(32)) eq_125(.in0(eq_125_in0), .in1(eq_125_in1), .out(eq_125_out));

	wire [31:0] eq_126_in0;
	wire [31:0] eq_126_in1;
	wire [0:0] eq_126_out;
	eq #(.WIDTH(32)) eq_126(.in0(eq_126_in0), .in1(eq_126_in1), .out(eq_126_out));

	wire [0:0] orOp_127_in0;
	wire [0:0] orOp_127_in1;
	wire [0:0] orOp_127_out;
	orOp #(.WIDTH(1)) orOp_127(.in0(orOp_127_in0), .in1(orOp_127_in1), .out(orOp_127_out));

	wire [31:0] eq_128_in0;
	wire [31:0] eq_128_in1;
	wire [0:0] eq_128_out;
	eq #(.WIDTH(32)) eq_128(.in0(eq_128_in0), .in1(eq_128_in1), .out(eq_128_out));

	wire [31:0] eq_129_in0;
	wire [31:0] eq_129_in1;
	wire [0:0] eq_129_out;
	eq #(.WIDTH(32)) eq_129(.in0(eq_129_in0), .in1(eq_129_in1), .out(eq_129_out));

	wire [31:0] eq_130_in0;
	wire [31:0] eq_130_in1;
	wire [0:0] eq_130_out;
	eq #(.WIDTH(32)) eq_130(.in0(eq_130_in0), .in1(eq_130_in1), .out(eq_130_out));

	wire [31:0] eq_131_in0;
	wire [31:0] eq_131_in1;
	wire [0:0] eq_131_out;
	eq #(.WIDTH(32)) eq_131(.in0(eq_131_in0), .in1(eq_131_in1), .out(eq_131_out));

	wire [0:0] orOp_132_in0;
	wire [0:0] orOp_132_in1;
	wire [0:0] orOp_132_out;
	orOp #(.WIDTH(1)) orOp_132(.in0(orOp_132_in0), .in1(orOp_132_in1), .out(orOp_132_out));

	wire [31:0] eq_133_in0;
	wire [31:0] eq_133_in1;
	wire [0:0] eq_133_out;
	eq #(.WIDTH(32)) eq_133(.in0(eq_133_in0), .in1(eq_133_in1), .out(eq_133_out));

	wire [31:0] eq_134_in0;
	wire [31:0] eq_134_in1;
	wire [0:0] eq_134_out;
	eq #(.WIDTH(32)) eq_134(.in0(eq_134_in0), .in1(eq_134_in1), .out(eq_134_out));

	wire [31:0] eq_135_in0;
	wire [31:0] eq_135_in1;
	wire [0:0] eq_135_out;
	eq #(.WIDTH(32)) eq_135(.in0(eq_135_in0), .in1(eq_135_in1), .out(eq_135_out));

	wire [31:0] eq_136_in0;
	wire [31:0] eq_136_in1;
	wire [0:0] eq_136_out;
	eq #(.WIDTH(32)) eq_136(.in0(eq_136_in0), .in1(eq_136_in1), .out(eq_136_out));

	wire [0:0] orOp_137_in0;
	wire [0:0] orOp_137_in1;
	wire [0:0] orOp_137_out;
	orOp #(.WIDTH(1)) orOp_137(.in0(orOp_137_in0), .in1(orOp_137_in1), .out(orOp_137_out));

	wire [31:0] eq_138_in0;
	wire [31:0] eq_138_in1;
	wire [0:0] eq_138_out;
	eq #(.WIDTH(32)) eq_138(.in0(eq_138_in0), .in1(eq_138_in1), .out(eq_138_out));

	wire [0:0] orOp_139_in0;
	wire [0:0] orOp_139_in1;
	wire [0:0] orOp_139_out;
	orOp #(.WIDTH(1)) orOp_139(.in0(orOp_139_in0), .in1(orOp_139_in1), .out(orOp_139_out));

	wire [31:0] eq_140_in0;
	wire [31:0] eq_140_in1;
	wire [0:0] eq_140_out;
	eq #(.WIDTH(32)) eq_140(.in0(eq_140_in0), .in1(eq_140_in1), .out(eq_140_out));

	wire [31:0] eq_141_in0;
	wire [31:0] eq_141_in1;
	wire [0:0] eq_141_out;
	eq #(.WIDTH(32)) eq_141(.in0(eq_141_in0), .in1(eq_141_in1), .out(eq_141_out));

	wire [31:0] eq_142_in0;
	wire [31:0] eq_142_in1;
	wire [0:0] eq_142_out;
	eq #(.WIDTH(32)) eq_142(.in0(eq_142_in0), .in1(eq_142_in1), .out(eq_142_out));

	wire [0:0] notOp_143_in0;
	wire [0:0] notOp_143_out;
	notOp #(.WIDTH(1)) notOp_143(.in(notOp_143_in0), .out(notOp_143_out));

	wire [0:0] andOp_144_in0;
	wire [0:0] andOp_144_in1;
	wire [0:0] andOp_144_out;
	andOp #(.WIDTH(1)) andOp_144(.in0(andOp_144_in0), .in1(andOp_144_in1), .out(andOp_144_out));

	wire [31:0] eq_145_in0;
	wire [31:0] eq_145_in1;
	wire [0:0] eq_145_out;
	eq #(.WIDTH(32)) eq_145(.in0(eq_145_in0), .in1(eq_145_in1), .out(eq_145_out));

	wire [31:0] eq_146_in0;
	wire [31:0] eq_146_in1;
	wire [0:0] eq_146_out;
	eq #(.WIDTH(32)) eq_146(.in0(eq_146_in0), .in1(eq_146_in1), .out(eq_146_out));

	wire [31:0] eq_147_in0;
	wire [31:0] eq_147_in1;
	wire [0:0] eq_147_out;
	eq #(.WIDTH(32)) eq_147(.in0(eq_147_in0), .in1(eq_147_in1), .out(eq_147_out));

	wire [31:0] eq_148_in0;
	wire [31:0] eq_148_in1;
	wire [0:0] eq_148_out;
	eq #(.WIDTH(32)) eq_148(.in0(eq_148_in0), .in1(eq_148_in1), .out(eq_148_out));

	wire [0:0] notOp_149_in0;
	wire [0:0] notOp_149_out;
	notOp #(.WIDTH(1)) notOp_149(.in(notOp_149_in0), .out(notOp_149_out));

	wire [0:0] andOp_150_in0;
	wire [0:0] andOp_150_in1;
	wire [0:0] andOp_150_out;
	andOp #(.WIDTH(1)) andOp_150(.in0(andOp_150_in0), .in1(andOp_150_in1), .out(andOp_150_out));

	wire [31:0] eq_151_in0;
	wire [31:0] eq_151_in1;
	wire [0:0] eq_151_out;
	eq #(.WIDTH(32)) eq_151(.in0(eq_151_in0), .in1(eq_151_in1), .out(eq_151_out));

	wire [31:0] eq_152_in0;
	wire [31:0] eq_152_in1;
	wire [0:0] eq_152_out;
	eq #(.WIDTH(32)) eq_152(.in0(eq_152_in0), .in1(eq_152_in1), .out(eq_152_out));

	wire [31:0] eq_153_in0;
	wire [31:0] eq_153_in1;
	wire [0:0] eq_153_out;
	eq #(.WIDTH(32)) eq_153(.in0(eq_153_in0), .in1(eq_153_in1), .out(eq_153_out));

	wire [31:0] eq_154_in0;
	wire [31:0] eq_154_in1;
	wire [0:0] eq_154_out;
	eq #(.WIDTH(32)) eq_154(.in0(eq_154_in0), .in1(eq_154_in1), .out(eq_154_out));

	wire [0:0] notOp_155_in0;
	wire [0:0] notOp_155_out;
	notOp #(.WIDTH(1)) notOp_155(.in(notOp_155_in0), .out(notOp_155_out));

	wire [0:0] andOp_156_in0;
	wire [0:0] andOp_156_in1;
	wire [0:0] andOp_156_out;
	andOp #(.WIDTH(1)) andOp_156(.in0(andOp_156_in0), .in1(andOp_156_in1), .out(andOp_156_out));

	wire [31:0] eq_157_in0;
	wire [31:0] eq_157_in1;
	wire [0:0] eq_157_out;
	eq #(.WIDTH(32)) eq_157(.in0(eq_157_in0), .in1(eq_157_in1), .out(eq_157_out));

	wire [0:0] notOp_158_in0;
	wire [0:0] notOp_158_out;
	notOp #(.WIDTH(1)) notOp_158(.in(notOp_158_in0), .out(notOp_158_out));

	wire [0:0] andOp_159_in0;
	wire [0:0] andOp_159_in1;
	wire [0:0] andOp_159_out;
	andOp #(.WIDTH(1)) andOp_159(.in0(andOp_159_in0), .in1(andOp_159_in1), .out(andOp_159_out));

	wire [31:0] eq_160_in0;
	wire [31:0] eq_160_in1;
	wire [0:0] eq_160_out;
	eq #(.WIDTH(32)) eq_160(.in0(eq_160_in0), .in1(eq_160_in1), .out(eq_160_out));

	wire [0:0] andOp_161_in0;
	wire [0:0] andOp_161_in1;
	wire [0:0] andOp_161_out;
	andOp #(.WIDTH(1)) andOp_161(.in0(andOp_161_in0), .in1(andOp_161_in1), .out(andOp_161_out));

	wire [31:0] concat_162_in0;
	wire [31:0] concat_162_in1;
	wire [63:0] concat_162_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_162(.in0(concat_162_in0), .in1(concat_162_in1), .out(concat_162_out));

	wire [31:0] concat_163_in0;
	wire [31:0] concat_163_in1;
	wire [63:0] concat_163_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_163(.in0(concat_163_in0), .in1(concat_163_in1), .out(concat_163_out));

	wire [0:0] andOp_164_in0;
	wire [0:0] andOp_164_in1;
	wire [0:0] andOp_164_out;
	andOp #(.WIDTH(1)) andOp_164(.in0(andOp_164_in0), .in1(andOp_164_in1), .out(andOp_164_out));

	wire [0:0] andOp_165_in0;
	wire [0:0] andOp_165_in1;
	wire [0:0] andOp_165_out;
	andOp #(.WIDTH(1)) andOp_165(.in0(andOp_165_in0), .in1(andOp_165_in1), .out(andOp_165_out));

	wire [0:0] andOp_166_in0;
	wire [0:0] andOp_166_in1;
	wire [0:0] andOp_166_out;
	andOp #(.WIDTH(1)) andOp_166(.in0(andOp_166_in0), .in1(andOp_166_in1), .out(andOp_166_out));

	wire [0:0] andOp_167_in0;
	wire [0:0] andOp_167_in1;
	wire [0:0] andOp_167_out;
	andOp #(.WIDTH(1)) andOp_167(.in0(andOp_167_in0), .in1(andOp_167_in1), .out(andOp_167_out));

	wire [0:0] andOp_168_in0;
	wire [0:0] andOp_168_in1;
	wire [0:0] andOp_168_out;
	andOp #(.WIDTH(1)) andOp_168(.in0(andOp_168_in0), .in1(andOp_168_in1), .out(andOp_168_out));

	wire [0:0] andOp_169_in0;
	wire [0:0] andOp_169_in1;
	wire [0:0] andOp_169_out;
	andOp #(.WIDTH(1)) andOp_169(.in0(andOp_169_in0), .in1(andOp_169_in1), .out(andOp_169_out));

	wire [0:0] andOp_170_in0;
	wire [0:0] andOp_170_in1;
	wire [0:0] andOp_170_out;
	andOp #(.WIDTH(1)) andOp_170(.in0(andOp_170_in0), .in1(andOp_170_in1), .out(andOp_170_out));

	wire [0:0] andOp_171_in0;
	wire [0:0] andOp_171_in1;
	wire [0:0] andOp_171_out;
	andOp #(.WIDTH(1)) andOp_171(.in0(andOp_171_in0), .in1(andOp_171_in1), .out(andOp_171_out));

	wire [0:0] andOp_172_in0;
	wire [0:0] andOp_172_in1;
	wire [0:0] andOp_172_out;
	andOp #(.WIDTH(1)) andOp_172(.in0(andOp_172_in0), .in1(andOp_172_in1), .out(andOp_172_out));

	wire [0:0] andOp_173_in0;
	wire [0:0] andOp_173_in1;
	wire [0:0] andOp_173_out;
	andOp #(.WIDTH(1)) andOp_173(.in0(andOp_173_in0), .in1(andOp_173_in1), .out(andOp_173_out));

	wire [0:0] andOp_174_in0;
	wire [0:0] andOp_174_in1;
	wire [0:0] andOp_174_out;
	andOp #(.WIDTH(1)) andOp_174(.in0(andOp_174_in0), .in1(andOp_174_in1), .out(andOp_174_out));

	wire [0:0] andOp_175_in0;
	wire [0:0] andOp_175_in1;
	wire [0:0] andOp_175_out;
	andOp #(.WIDTH(1)) andOp_175(.in0(andOp_175_in0), .in1(andOp_175_in1), .out(andOp_175_out));

	wire [0:0] andOp_176_in0;
	wire [0:0] andOp_176_in1;
	wire [0:0] andOp_176_out;
	andOp #(.WIDTH(1)) andOp_176(.in0(andOp_176_in0), .in1(andOp_176_in1), .out(andOp_176_out));

	wire [0:0] andOp_177_in0;
	wire [0:0] andOp_177_in1;
	wire [0:0] andOp_177_out;
	andOp #(.WIDTH(1)) andOp_177(.in0(andOp_177_in0), .in1(andOp_177_in1), .out(andOp_177_out));

	wire [0:0] andOp_178_in0;
	wire [0:0] andOp_178_in1;
	wire [0:0] andOp_178_out;
	andOp #(.WIDTH(1)) andOp_178(.in0(andOp_178_in0), .in1(andOp_178_in1), .out(andOp_178_out));

	wire [31:0] concat_179_in0;
	wire [31:0] concat_179_in1;
	wire [63:0] concat_179_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_179(.in0(concat_179_in0), .in1(concat_179_in1), .out(concat_179_out));

	wire [31:0] concat_180_in0;
	wire [31:0] concat_180_in1;
	wire [63:0] concat_180_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_180(.in0(concat_180_in0), .in1(concat_180_in1), .out(concat_180_out));

	wire [0:0] andOp_181_in0;
	wire [0:0] andOp_181_in1;
	wire [0:0] andOp_181_out;
	andOp #(.WIDTH(1)) andOp_181(.in0(andOp_181_in0), .in1(andOp_181_in1), .out(andOp_181_out));

	wire [0:0] andOp_182_in0;
	wire [0:0] andOp_182_in1;
	wire [0:0] andOp_182_out;
	andOp #(.WIDTH(1)) andOp_182(.in0(andOp_182_in0), .in1(andOp_182_in1), .out(andOp_182_out));

	wire [0:0] andOp_183_in0;
	wire [0:0] andOp_183_in1;
	wire [0:0] andOp_183_out;
	andOp #(.WIDTH(1)) andOp_183(.in0(andOp_183_in0), .in1(andOp_183_in1), .out(andOp_183_out));

	wire [0:0] andOp_184_in0;
	wire [0:0] andOp_184_in1;
	wire [0:0] andOp_184_out;
	andOp #(.WIDTH(1)) andOp_184(.in0(andOp_184_in0), .in1(andOp_184_in1), .out(andOp_184_out));

	wire [0:0] andOp_185_in0;
	wire [0:0] andOp_185_in1;
	wire [0:0] andOp_185_out;
	andOp #(.WIDTH(1)) andOp_185(.in0(andOp_185_in0), .in1(andOp_185_in1), .out(andOp_185_out));

	wire [0:0] andOp_186_in0;
	wire [0:0] andOp_186_in1;
	wire [0:0] andOp_186_out;
	andOp #(.WIDTH(1)) andOp_186(.in0(andOp_186_in0), .in1(andOp_186_in1), .out(andOp_186_out));

	wire [0:0] andOp_187_in0;
	wire [0:0] andOp_187_in1;
	wire [0:0] andOp_187_out;
	andOp #(.WIDTH(1)) andOp_187(.in0(andOp_187_in0), .in1(andOp_187_in1), .out(andOp_187_out));

	wire [0:0] andOp_188_in0;
	wire [0:0] andOp_188_in1;
	wire [0:0] andOp_188_out;
	andOp #(.WIDTH(1)) andOp_188(.in0(andOp_188_in0), .in1(andOp_188_in1), .out(andOp_188_out));

	wire [0:0] andOp_189_in0;
	wire [0:0] andOp_189_in1;
	wire [0:0] andOp_189_out;
	andOp #(.WIDTH(1)) andOp_189(.in0(andOp_189_in0), .in1(andOp_189_in1), .out(andOp_189_out));

	wire [0:0] andOp_190_in0;
	wire [0:0] andOp_190_in1;
	wire [0:0] andOp_190_out;
	andOp #(.WIDTH(1)) andOp_190(.in0(andOp_190_in0), .in1(andOp_190_in1), .out(andOp_190_out));

	wire [0:0] andOp_191_in0;
	wire [0:0] andOp_191_in1;
	wire [0:0] andOp_191_out;
	andOp #(.WIDTH(1)) andOp_191(.in0(andOp_191_in0), .in1(andOp_191_in1), .out(andOp_191_out));

	wire [0:0] andOp_192_in0;
	wire [0:0] andOp_192_in1;
	wire [0:0] andOp_192_out;
	andOp #(.WIDTH(1)) andOp_192(.in0(andOp_192_in0), .in1(andOp_192_in1), .out(andOp_192_out));

	wire [0:0] andOp_193_in0;
	wire [0:0] andOp_193_in1;
	wire [0:0] andOp_193_out;
	andOp #(.WIDTH(1)) andOp_193(.in0(andOp_193_in0), .in1(andOp_193_in1), .out(andOp_193_out));

	wire [0:0] andOp_194_in0;
	wire [0:0] andOp_194_in1;
	wire [0:0] andOp_194_out;
	andOp #(.WIDTH(1)) andOp_194(.in0(andOp_194_in0), .in1(andOp_194_in1), .out(andOp_194_out));

	wire [0:0] andOp_195_in0;
	wire [0:0] andOp_195_in1;
	wire [0:0] andOp_195_out;
	andOp #(.WIDTH(1)) andOp_195(.in0(andOp_195_in0), .in1(andOp_195_in1), .out(andOp_195_out));

	wire [0:0] andOp_196_in0;
	wire [0:0] andOp_196_in1;
	wire [0:0] andOp_196_out;
	andOp #(.WIDTH(1)) andOp_196(.in0(andOp_196_in0), .in1(andOp_196_in1), .out(andOp_196_out));

	wire [0:0] andOp_197_in0;
	wire [0:0] andOp_197_in1;
	wire [0:0] andOp_197_out;
	andOp #(.WIDTH(1)) andOp_197(.in0(andOp_197_in0), .in1(andOp_197_in1), .out(andOp_197_out));

	wire [0:0] notOp_198_in0;
	wire [0:0] notOp_198_out;
	notOp #(.WIDTH(1)) notOp_198(.in(notOp_198_in0), .out(notOp_198_out));

	wire [0:0] andOp_199_in0;
	wire [0:0] andOp_199_in1;
	wire [0:0] andOp_199_out;
	andOp #(.WIDTH(1)) andOp_199(.in0(andOp_199_in0), .in1(andOp_199_in1), .out(andOp_199_out));

	wire [0:0] notOp_200_in0;
	wire [0:0] notOp_200_out;
	notOp #(.WIDTH(1)) notOp_200(.in(notOp_200_in0), .out(notOp_200_out));

	wire [0:0] andOp_201_in0;
	wire [0:0] andOp_201_in1;
	wire [0:0] andOp_201_out;
	andOp #(.WIDTH(1)) andOp_201(.in0(andOp_201_in0), .in1(andOp_201_in1), .out(andOp_201_out));

	wire [0:0] notOp_202_in0;
	wire [0:0] notOp_202_out;
	notOp #(.WIDTH(1)) notOp_202(.in(notOp_202_in0), .out(notOp_202_out));

	wire [0:0] andOp_203_in0;
	wire [0:0] andOp_203_in1;
	wire [0:0] andOp_203_out;
	andOp #(.WIDTH(1)) andOp_203(.in0(andOp_203_in0), .in1(andOp_203_in1), .out(andOp_203_out));

	wire [0:0] notOp_204_in0;
	wire [0:0] notOp_204_out;
	notOp #(.WIDTH(1)) notOp_204(.in(notOp_204_in0), .out(notOp_204_out));

	wire [0:0] andOp_205_in0;
	wire [0:0] andOp_205_in1;
	wire [0:0] andOp_205_out;
	andOp #(.WIDTH(1)) andOp_205(.in0(andOp_205_in0), .in1(andOp_205_in1), .out(andOp_205_out));

	wire [0:0] notOp_206_in0;
	wire [0:0] notOp_206_out;
	notOp #(.WIDTH(1)) notOp_206(.in(notOp_206_in0), .out(notOp_206_out));

	wire [0:0] andOp_207_in0;
	wire [0:0] andOp_207_in1;
	wire [0:0] andOp_207_out;
	andOp #(.WIDTH(1)) andOp_207(.in0(andOp_207_in0), .in1(andOp_207_in1), .out(andOp_207_out));

	wire [0:0] notOp_208_in0;
	wire [0:0] notOp_208_out;
	notOp #(.WIDTH(1)) notOp_208(.in(notOp_208_in0), .out(notOp_208_out));

	wire [0:0] andOp_209_in0;
	wire [0:0] andOp_209_in1;
	wire [0:0] andOp_209_out;
	andOp #(.WIDTH(1)) andOp_209(.in0(andOp_209_in0), .in1(andOp_209_in1), .out(andOp_209_out));

	wire [0:0] notOp_210_in0;
	wire [0:0] notOp_210_out;
	notOp #(.WIDTH(1)) notOp_210(.in(notOp_210_in0), .out(notOp_210_out));

	wire [0:0] andOp_211_in0;
	wire [0:0] andOp_211_in1;
	wire [0:0] andOp_211_out;
	andOp #(.WIDTH(1)) andOp_211(.in0(andOp_211_in0), .in1(andOp_211_in1), .out(andOp_211_out));

	wire [0:0] notOp_212_in0;
	wire [0:0] notOp_212_out;
	notOp #(.WIDTH(1)) notOp_212(.in(notOp_212_in0), .out(notOp_212_out));

	wire [0:0] andOp_213_in0;
	wire [0:0] andOp_213_in1;
	wire [0:0] andOp_213_out;
	andOp #(.WIDTH(1)) andOp_213(.in0(andOp_213_in0), .in1(andOp_213_in1), .out(andOp_213_out));

	wire [0:0] notOp_214_in0;
	wire [0:0] notOp_214_out;
	notOp #(.WIDTH(1)) notOp_214(.in(notOp_214_in0), .out(notOp_214_out));

	wire [0:0] andOp_215_in0;
	wire [0:0] andOp_215_in1;
	wire [0:0] andOp_215_out;
	andOp #(.WIDTH(1)) andOp_215(.in0(andOp_215_in0), .in1(andOp_215_in1), .out(andOp_215_out));

	wire [0:0] notOp_216_in0;
	wire [0:0] notOp_216_out;
	notOp #(.WIDTH(1)) notOp_216(.in(notOp_216_in0), .out(notOp_216_out));

	wire [0:0] andOp_217_in0;
	wire [0:0] andOp_217_in1;
	wire [0:0] andOp_217_out;
	andOp #(.WIDTH(1)) andOp_217(.in0(andOp_217_in0), .in1(andOp_217_in1), .out(andOp_217_out));

	wire [31:0] eq_218_in0;
	wire [31:0] eq_218_in1;
	wire [0:0] eq_218_out;
	eq #(.WIDTH(32)) eq_218(.in0(eq_218_in0), .in1(eq_218_in1), .out(eq_218_out));

	wire [31:0] eq_219_in0;
	wire [31:0] eq_219_in1;
	wire [0:0] eq_219_out;
	eq #(.WIDTH(32)) eq_219(.in0(eq_219_in0), .in1(eq_219_in1), .out(eq_219_out));

	wire [0:0] andOp_220_in0;
	wire [0:0] andOp_220_in1;
	wire [0:0] andOp_220_out;
	andOp #(.WIDTH(1)) andOp_220(.in0(andOp_220_in0), .in1(andOp_220_in1), .out(andOp_220_out));

	wire [0:0] andOp_221_in0;
	wire [0:0] andOp_221_in1;
	wire [0:0] andOp_221_out;
	andOp #(.WIDTH(1)) andOp_221(.in0(andOp_221_in0), .in1(andOp_221_in1), .out(andOp_221_out));

	wire [0:0] andOp_222_in0;
	wire [0:0] andOp_222_in1;
	wire [0:0] andOp_222_out;
	andOp #(.WIDTH(1)) andOp_222(.in0(andOp_222_in0), .in1(andOp_222_in1), .out(andOp_222_out));

	wire [31:0] eq_223_in0;
	wire [31:0] eq_223_in1;
	wire [0:0] eq_223_out;
	eq #(.WIDTH(32)) eq_223(.in0(eq_223_in0), .in1(eq_223_in1), .out(eq_223_out));

	wire [31:0] eq_224_in0;
	wire [31:0] eq_224_in1;
	wire [0:0] eq_224_out;
	eq #(.WIDTH(32)) eq_224(.in0(eq_224_in0), .in1(eq_224_in1), .out(eq_224_out));

	wire [31:0] eq_225_in0;
	wire [31:0] eq_225_in1;
	wire [0:0] eq_225_out;
	eq #(.WIDTH(32)) eq_225(.in0(eq_225_in0), .in1(eq_225_in1), .out(eq_225_out));

	wire [31:0] eq_226_in0;
	wire [31:0] eq_226_in1;
	wire [0:0] eq_226_out;
	eq #(.WIDTH(32)) eq_226(.in0(eq_226_in0), .in1(eq_226_in1), .out(eq_226_out));

	wire [31:0] eq_227_in0;
	wire [31:0] eq_227_in1;
	wire [0:0] eq_227_out;
	eq #(.WIDTH(32)) eq_227(.in0(eq_227_in0), .in1(eq_227_in1), .out(eq_227_out));

	wire [31:0] eq_228_in0;
	wire [31:0] eq_228_in1;
	wire [0:0] eq_228_out;
	eq #(.WIDTH(32)) eq_228(.in0(eq_228_in0), .in1(eq_228_in1), .out(eq_228_out));

	wire [31:0] eq_229_in0;
	wire [31:0] eq_229_in1;
	wire [0:0] eq_229_out;
	eq #(.WIDTH(32)) eq_229(.in0(eq_229_in0), .in1(eq_229_in1), .out(eq_229_out));

	wire [0:0] andOp_230_in0;
	wire [0:0] andOp_230_in1;
	wire [0:0] andOp_230_out;
	andOp #(.WIDTH(1)) andOp_230(.in0(andOp_230_in0), .in1(andOp_230_in1), .out(andOp_230_out));

	wire [0:0] andOp_231_in0;
	wire [0:0] andOp_231_in1;
	wire [0:0] andOp_231_out;
	andOp #(.WIDTH(1)) andOp_231(.in0(andOp_231_in0), .in1(andOp_231_in1), .out(andOp_231_out));

	wire [31:0] eq_232_in0;
	wire [31:0] eq_232_in1;
	wire [0:0] eq_232_out;
	eq #(.WIDTH(32)) eq_232(.in0(eq_232_in0), .in1(eq_232_in1), .out(eq_232_out));

	wire [31:0] eq_233_in0;
	wire [31:0] eq_233_in1;
	wire [0:0] eq_233_out;
	eq #(.WIDTH(32)) eq_233(.in0(eq_233_in0), .in1(eq_233_in1), .out(eq_233_out));

	wire [31:0] eq_234_in0;
	wire [31:0] eq_234_in1;
	wire [0:0] eq_234_out;
	eq #(.WIDTH(32)) eq_234(.in0(eq_234_in0), .in1(eq_234_in1), .out(eq_234_out));

	wire [31:0] eq_235_in0;
	wire [31:0] eq_235_in1;
	wire [0:0] eq_235_out;
	eq #(.WIDTH(32)) eq_235(.in0(eq_235_in0), .in1(eq_235_in1), .out(eq_235_out));

	wire [31:0] eq_236_in0;
	wire [31:0] eq_236_in1;
	wire [0:0] eq_236_out;
	eq #(.WIDTH(32)) eq_236(.in0(eq_236_in0), .in1(eq_236_in1), .out(eq_236_out));

	wire [31:0] eq_237_in0;
	wire [31:0] eq_237_in1;
	wire [0:0] eq_237_out;
	eq #(.WIDTH(32)) eq_237(.in0(eq_237_in0), .in1(eq_237_in1), .out(eq_237_out));

	wire [31:0] eq_238_in0;
	wire [31:0] eq_238_in1;
	wire [0:0] eq_238_out;
	eq #(.WIDTH(32)) eq_238(.in0(eq_238_in0), .in1(eq_238_in1), .out(eq_238_out));

	wire [31:0] eq_239_in0;
	wire [31:0] eq_239_in1;
	wire [0:0] eq_239_out;
	eq #(.WIDTH(32)) eq_239(.in0(eq_239_in0), .in1(eq_239_in1), .out(eq_239_out));

	wire [0:0] andOp_240_in0;
	wire [0:0] andOp_240_in1;
	wire [0:0] andOp_240_out;
	andOp #(.WIDTH(1)) andOp_240(.in0(andOp_240_in0), .in1(andOp_240_in1), .out(andOp_240_out));

	wire [0:0] andOp_241_in0;
	wire [0:0] andOp_241_in1;
	wire [0:0] andOp_241_out;
	andOp #(.WIDTH(1)) andOp_241(.in0(andOp_241_in0), .in1(andOp_241_in1), .out(andOp_241_out));

	wire [0:0] andOp_242_in0;
	wire [0:0] andOp_242_in1;
	wire [0:0] andOp_242_out;
	andOp #(.WIDTH(1)) andOp_242(.in0(andOp_242_in0), .in1(andOp_242_in1), .out(andOp_242_out));

	wire [0:0] andOp_243_in0;
	wire [0:0] andOp_243_in1;
	wire [0:0] andOp_243_out;
	andOp #(.WIDTH(1)) andOp_243(.in0(andOp_243_in0), .in1(andOp_243_in1), .out(andOp_243_out));

	wire [0:0] andOp_244_in0;
	wire [0:0] andOp_244_in1;
	wire [0:0] andOp_244_out;
	andOp #(.WIDTH(1)) andOp_244(.in0(andOp_244_in0), .in1(andOp_244_in1), .out(andOp_244_out));

	wire [0:0] andOp_245_in0;
	wire [0:0] andOp_245_in1;
	wire [0:0] andOp_245_out;
	andOp #(.WIDTH(1)) andOp_245(.in0(andOp_245_in0), .in1(andOp_245_in1), .out(andOp_245_out));

	wire [0:0] andOp_246_in0;
	wire [0:0] andOp_246_in1;
	wire [0:0] andOp_246_out;
	andOp #(.WIDTH(1)) andOp_246(.in0(andOp_246_in0), .in1(andOp_246_in1), .out(andOp_246_out));

	wire [0:0] andOp_247_in0;
	wire [0:0] andOp_247_in1;
	wire [0:0] andOp_247_out;
	andOp #(.WIDTH(1)) andOp_247(.in0(andOp_247_in0), .in1(andOp_247_in1), .out(andOp_247_out));

	wire [0:0] andOp_248_in0;
	wire [0:0] andOp_248_in1;
	wire [0:0] andOp_248_out;
	andOp #(.WIDTH(1)) andOp_248(.in0(andOp_248_in0), .in1(andOp_248_in1), .out(andOp_248_out));

	wire [0:0] andOp_249_in0;
	wire [0:0] andOp_249_in1;
	wire [0:0] andOp_249_out;
	andOp #(.WIDTH(1)) andOp_249(.in0(andOp_249_in0), .in1(andOp_249_in1), .out(andOp_249_out));

	wire [0:0] andOp_250_in0;
	wire [0:0] andOp_250_in1;
	wire [0:0] andOp_250_out;
	andOp #(.WIDTH(1)) andOp_250(.in0(andOp_250_in0), .in1(andOp_250_in1), .out(andOp_250_out));

	wire [0:0] andOp_251_in0;
	wire [0:0] andOp_251_in1;
	wire [0:0] andOp_251_out;
	andOp #(.WIDTH(1)) andOp_251(.in0(andOp_251_in0), .in1(andOp_251_in1), .out(andOp_251_out));

	wire [0:0] andOp_252_in0;
	wire [0:0] andOp_252_in1;
	wire [0:0] andOp_252_out;
	andOp #(.WIDTH(1)) andOp_252(.in0(andOp_252_in0), .in1(andOp_252_in1), .out(andOp_252_out));

	wire [0:0] andOp_253_in0;
	wire [0:0] andOp_253_in1;
	wire [0:0] andOp_253_out;
	andOp #(.WIDTH(1)) andOp_253(.in0(andOp_253_in0), .in1(andOp_253_in1), .out(andOp_253_out));

	wire [0:0] andOp_254_in0;
	wire [0:0] andOp_254_in1;
	wire [0:0] andOp_254_out;
	andOp #(.WIDTH(1)) andOp_254(.in0(andOp_254_in0), .in1(andOp_254_in1), .out(andOp_254_out));

	// End Functional Units

	reg [31:0] data_store_0_0;
	reg [31:0] data_store_0_1;
	reg [31:0] data_store_0_2;
	reg [31:0] data_store_0_3;
	reg [31:0] data_store_0_5;
	reg [31:0] data_store_1_11;
	reg [31:0] data_store_1_13;
	reg [31:0] data_store_1_15;
	reg [31:0] data_store_1_7;
	reg [31:0] data_store_1_9;
	reg [31:0] data_store_2_17;
	reg [31:0] data_store_2_19;
	reg [31:0] data_store_2_21;
	reg [31:0] data_store_2_23;
	reg [31:0] data_store_2_25;
	reg [31:0] data_store_3_27;
	reg [31:0] data_store_3_29;
	reg [31:0] data_store_3_31;
	reg [31:0] data_store_3_33;
	reg [31:0] data_store_3_35;
	reg [0:0] data_store_3_37;
	reg [31:0] data_store_4_38;
	reg [31:0] data_store_4_40;
	reg [31:0] data_store_4_42;
	reg [31:0] data_store_4_44;
	reg [31:0] data_store_4_46;
	reg [0:0] data_store_4_48;
	reg [31:0] data_store_5_50;
	reg [31:0] data_store_5_52;
	reg [31:0] data_store_5_54;
	reg [31:0] data_store_5_56;
	reg [31:0] data_store_5_58;
	reg [0:0] data_store_5_60;
	reg [31:0] data_store_6_62;
	reg [31:0] data_store_6_64;
	reg [31:0] data_store_6_66;
	reg [31:0] data_store_6_68;
	reg [31:0] data_store_6_70;
	reg [0:0] data_store_6_72;
	reg [31:0] data_store_7_74;
	reg [31:0] data_store_7_76;
	reg [31:0] data_store_7_78;
	reg [31:0] data_store_7_80;
	reg [31:0] data_store_7_82;
	reg [31:0] global_state;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_3_last_state;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;
	reg [31:0] state_4_last_state;
	reg [31:0] state_5_entry_BB_reg;
	reg [0:0] state_5_is_active;
	reg [31:0] state_5_last_BB_reg;
	reg [31:0] state_5_last_state;
	reg [31:0] state_6_entry_BB_reg;
	reg [0:0] state_6_is_active;
	reg [31:0] state_6_last_BB_reg;
	reg [31:0] state_6_last_state;
	reg [31:0] state_7_entry_BB_reg;
	reg [0:0] state_7_is_active;
	reg [31:0] state_7_last_BB_reg;
	reg [31:0] state_7_last_state;

	// controller for add_add10.add_add10_in0
	// controller for add_add10.add_add10_in1
	// Insensitive connections
	assign add_add10_in0 = phi_phi7_out;
	assign add_add10_in1 = 32'd9;
	// controller for add_add11.add_add11_in0
	// controller for add_add11.add_add11_in1
	// Insensitive connections
	assign add_add11_in0 = phi_phi7_out;
	assign add_add11_in1 = 32'd1;
	// controller for add_add17.add_add17_in0
	// controller for add_add17.add_add17_in1
	// Insensitive connections
	assign add_add17_in0 = mul_mul16_out;
	assign add_add17_in1 = ram_rdata_0;
	// controller for add_add2.add_add2_in0
	// controller for add_add2.add_add2_in1
	// Insensitive connections
	assign add_add2_in0 = phi_phi1_out;
	assign add_add2_in1 = 32'd12;
	// controller for add_add25.add_add25_in0
	// controller for add_add25.add_add25_in1
	// Insensitive connections
	assign add_add25_in0 = data_in_7_75_out_data;
	assign add_add25_in1 = 32'd1;
	// controller for add_add9.add_add9_in0
	// controller for add_add9.add_add9_in1
	// Insensitive connections
	assign add_add9_in0 = phi_phi7_out;
	assign add_add9_in1 = data_in_3_32_out_data;
	// controller for andOp_100.andOp_100_in0
	// controller for andOp_100.andOp_100_in1
	// Insensitive connections
	assign andOp_100_in0 = bb_4_active_in_state_7_out_data;
	assign andOp_100_in1 = state_7_is_active;
	// controller for andOp_102.andOp_102_in0
	// controller for andOp_102.andOp_102_in1
	// Insensitive connections
	assign andOp_102_in0 = andOp_100_out;
	assign andOp_102_in1 = data_in_7_84_out_data;
	// controller for andOp_104.andOp_104_in0
	// controller for andOp_104.andOp_104_in1
	// Insensitive connections
	assign andOp_104_in0 = andOp_100_out;
	assign andOp_104_in1 = notOp_103_out;
	// controller for andOp_105.andOp_105_in0
	// controller for andOp_105.andOp_105_in1
	// Insensitive connections
	assign andOp_105_in0 = bb_4_active_in_state_7_out_data;
	assign andOp_105_in1 = state_7_is_active;
	// controller for andOp_107.andOp_107_in0
	// controller for andOp_107.andOp_107_in1
	// Insensitive connections
	assign andOp_107_in0 = andOp_105_out;
	assign andOp_107_in1 = data_in_7_84_out_data;
	// controller for andOp_109.andOp_109_in0
	// controller for andOp_109.andOp_109_in1
	// Insensitive connections
	assign andOp_109_in0 = andOp_105_out;
	assign andOp_109_in1 = notOp_108_out;
	// controller for andOp_110.andOp_110_in0
	// controller for andOp_110.andOp_110_in1
	// Insensitive connections
	assign andOp_110_in0 = bb_4_active_in_state_7_out_data;
	assign andOp_110_in1 = state_7_is_active;
	// controller for andOp_112.andOp_112_in0
	// controller for andOp_112.andOp_112_in1
	// Insensitive connections
	assign andOp_112_in0 = andOp_110_out;
	assign andOp_112_in1 = data_in_7_84_out_data;
	// controller for andOp_114.andOp_114_in0
	// controller for andOp_114.andOp_114_in1
	// Insensitive connections
	assign andOp_114_in0 = andOp_110_out;
	assign andOp_114_in1 = notOp_113_out;
	// controller for andOp_115.andOp_115_in0
	// controller for andOp_115.andOp_115_in1
	// Insensitive connections
	assign andOp_115_in0 = bb_3_active_in_state_7_out_data;
	assign andOp_115_in1 = state_7_is_active;
	// controller for andOp_117.andOp_117_in0
	// controller for andOp_117.andOp_117_in1
	// Insensitive connections
	assign andOp_117_in0 = andOp_115_out;
	assign andOp_117_in1 = icmp_icmp26_out;
	// controller for andOp_119.andOp_119_in0
	// controller for andOp_119.andOp_119_in1
	// Insensitive connections
	assign andOp_119_in0 = andOp_115_out;
	assign andOp_119_in1 = notOp_118_out;
	// controller for andOp_120.andOp_120_in0
	// controller for andOp_120.andOp_120_in1
	// Insensitive connections
	assign andOp_120_in0 = bb_4_active_in_state_7_out_data;
	assign andOp_120_in1 = state_7_is_active;
	// controller for andOp_122.andOp_122_in0
	// controller for andOp_122.andOp_122_in1
	// Insensitive connections
	assign andOp_122_in0 = andOp_120_out;
	assign andOp_122_in1 = data_in_7_84_out_data;
	// controller for andOp_124.andOp_124_in0
	// controller for andOp_124.andOp_124_in1
	// Insensitive connections
	assign andOp_124_in0 = andOp_120_out;
	assign andOp_124_in1 = notOp_123_out;
	// controller for andOp_144.andOp_144_in0
	// controller for andOp_144.andOp_144_in1
	// Insensitive connections
	assign andOp_144_in0 = notOp_143_out;
	assign andOp_144_in1 = andOp_85_out;
	// controller for andOp_150.andOp_150_in0
	// controller for andOp_150.andOp_150_in1
	// Insensitive connections
	assign andOp_150_in0 = notOp_149_out;
	assign andOp_150_in1 = andOp_87_out;
	// controller for andOp_156.andOp_156_in0
	// controller for andOp_156.andOp_156_in1
	// Insensitive connections
	assign andOp_156_in0 = notOp_155_out;
	assign andOp_156_in1 = andOp_117_out;
	// controller for andOp_159.andOp_159_in0
	// controller for andOp_159.andOp_159_in1
	// Insensitive connections
	assign andOp_159_in0 = notOp_158_out;
	assign andOp_159_in1 = andOp_97_out;
	// controller for andOp_161.andOp_161_in0
	// controller for andOp_161.andOp_161_in1
	// Insensitive connections
	assign andOp_161_in0 = bb_2_active_in_state_0_out_data;
	assign andOp_161_in1 = state_0_is_active;
	// controller for andOp_164.andOp_164_in0
	// controller for andOp_164.andOp_164_in1
	// Insensitive connections
	assign andOp_164_in0 = bb_2_active_in_state_0_out_data;
	assign andOp_164_in1 = state_0_is_active;
	// controller for andOp_165.andOp_165_in0
	// controller for andOp_165.andOp_165_in1
	// Insensitive connections
	assign andOp_165_in0 = bb_2_active_in_state_0_out_data;
	assign andOp_165_in1 = state_0_is_active;
	// controller for andOp_166.andOp_166_in0
	// controller for andOp_166.andOp_166_in1
	// Insensitive connections
	assign andOp_166_in0 = bb_2_active_in_state_0_out_data;
	assign andOp_166_in1 = state_0_is_active;
	// controller for andOp_167.andOp_167_in0
	// controller for andOp_167.andOp_167_in1
	// Insensitive connections
	assign andOp_167_in0 = bb_2_active_in_state_0_out_data;
	assign andOp_167_in1 = state_0_is_active;
	// controller for andOp_168.andOp_168_in0
	// controller for andOp_168.andOp_168_in1
	// Insensitive connections
	assign andOp_168_in0 = bb_2_active_in_state_0_out_data;
	assign andOp_168_in1 = state_0_is_active;
	// controller for andOp_169.andOp_169_in0
	// controller for andOp_169.andOp_169_in1
	// Insensitive connections
	assign andOp_169_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_169_in1 = state_3_is_active;
	// controller for andOp_170.andOp_170_in0
	// controller for andOp_170.andOp_170_in1
	// Insensitive connections
	assign andOp_170_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_170_in1 = state_3_is_active;
	// controller for andOp_171.andOp_171_in0
	// controller for andOp_171.andOp_171_in1
	// Insensitive connections
	assign andOp_171_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_171_in1 = state_3_is_active;
	// controller for andOp_172.andOp_172_in0
	// controller for andOp_172.andOp_172_in1
	// Insensitive connections
	assign andOp_172_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_172_in1 = state_4_is_active;
	// controller for andOp_173.andOp_173_in0
	// controller for andOp_173.andOp_173_in1
	// Insensitive connections
	assign andOp_173_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_173_in1 = state_4_is_active;
	// controller for andOp_174.andOp_174_in0
	// controller for andOp_174.andOp_174_in1
	// Insensitive connections
	assign andOp_174_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_174_in1 = state_4_is_active;
	// controller for andOp_175.andOp_175_in0
	// controller for andOp_175.andOp_175_in1
	// Insensitive connections
	assign andOp_175_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_175_in1 = state_4_is_active;
	// controller for andOp_176.andOp_176_in0
	// controller for andOp_176.andOp_176_in1
	// Insensitive connections
	assign andOp_176_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_176_in1 = state_4_is_active;
	// controller for andOp_177.andOp_177_in0
	// controller for andOp_177.andOp_177_in1
	// Insensitive connections
	assign andOp_177_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_177_in1 = state_4_is_active;
	// controller for andOp_178.andOp_178_in0
	// controller for andOp_178.andOp_178_in1
	// Insensitive connections
	assign andOp_178_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_178_in1 = state_3_is_active;
	// controller for andOp_181.andOp_181_in0
	// controller for andOp_181.andOp_181_in1
	// Insensitive connections
	assign andOp_181_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_181_in1 = state_3_is_active;
	// controller for andOp_182.andOp_182_in0
	// controller for andOp_182.andOp_182_in1
	// Insensitive connections
	assign andOp_182_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_182_in1 = state_3_is_active;
	// controller for andOp_183.andOp_183_in0
	// controller for andOp_183.andOp_183_in1
	// Insensitive connections
	assign andOp_183_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_183_in1 = state_3_is_active;
	// controller for andOp_184.andOp_184_in0
	// controller for andOp_184.andOp_184_in1
	// Insensitive connections
	assign andOp_184_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_184_in1 = state_3_is_active;
	// controller for andOp_185.andOp_185_in0
	// controller for andOp_185.andOp_185_in1
	// Insensitive connections
	assign andOp_185_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_185_in1 = state_4_is_active;
	// controller for andOp_186.andOp_186_in0
	// controller for andOp_186.andOp_186_in1
	// Insensitive connections
	assign andOp_186_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_186_in1 = state_4_is_active;
	// controller for andOp_187.andOp_187_in0
	// controller for andOp_187.andOp_187_in1
	// Insensitive connections
	assign andOp_187_in0 = bb_1_active_in_state_7_out_data;
	assign andOp_187_in1 = state_7_is_active;
	// controller for andOp_188.andOp_188_in0
	// controller for andOp_188.andOp_188_in1
	// Insensitive connections
	assign andOp_188_in0 = bb_3_active_in_state_7_out_data;
	assign andOp_188_in1 = state_7_is_active;
	// controller for andOp_189.andOp_189_in0
	// controller for andOp_189.andOp_189_in1
	// Insensitive connections
	assign andOp_189_in0 = bb_3_active_in_state_7_out_data;
	assign andOp_189_in1 = state_7_is_active;
	// controller for andOp_190.andOp_190_in0
	// controller for andOp_190.andOp_190_in1
	// Insensitive connections
	assign andOp_190_in0 = bb_2_active_in_state_0_out_data;
	assign andOp_190_in1 = state_0_is_active;
	// controller for andOp_191.andOp_191_in0
	// controller for andOp_191.andOp_191_in1
	// Insensitive connections
	assign andOp_191_in0 = bb_2_active_in_state_1_out_data;
	assign andOp_191_in1 = state_1_is_active;
	// controller for andOp_192.andOp_192_in0
	// controller for andOp_192.andOp_192_in1
	// Insensitive connections
	assign andOp_192_in0 = bb_2_active_in_state_2_out_data;
	assign andOp_192_in1 = state_2_is_active;
	// controller for andOp_193.andOp_193_in0
	// controller for andOp_193.andOp_193_in1
	// Insensitive connections
	assign andOp_193_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_193_in1 = state_3_is_active;
	// controller for andOp_194.andOp_194_in0
	// controller for andOp_194.andOp_194_in1
	// Insensitive connections
	assign andOp_194_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_194_in1 = state_4_is_active;
	// controller for andOp_195.andOp_195_in0
	// controller for andOp_195.andOp_195_in1
	// Insensitive connections
	assign andOp_195_in0 = bb_4_active_in_state_5_out_data;
	assign andOp_195_in1 = state_5_is_active;
	// controller for andOp_196.andOp_196_in0
	// controller for andOp_196.andOp_196_in1
	// Insensitive connections
	assign andOp_196_in0 = bb_4_active_in_state_6_out_data;
	assign andOp_196_in1 = state_6_is_active;
	// controller for andOp_197.andOp_197_in0
	// controller for andOp_197.andOp_197_in1
	// Insensitive connections
	assign andOp_197_in0 = bb_1_active_in_state_7_out_data;
	assign andOp_197_in1 = state_7_is_active;
	// controller for andOp_199.andOp_199_in0
	// controller for andOp_199.andOp_199_in1
	// Insensitive connections
	assign andOp_199_in0 = notOp_198_out;
	assign andOp_199_in1 = 1'd1;
	// controller for andOp_201.andOp_201_in0
	// controller for andOp_201.andOp_201_in1
	// Insensitive connections
	assign andOp_201_in0 = notOp_200_out;
	assign andOp_201_in1 = 1'd1;
	// controller for andOp_203.andOp_203_in0
	// controller for andOp_203.andOp_203_in1
	// Insensitive connections
	assign andOp_203_in0 = notOp_202_out;
	assign andOp_203_in1 = 1'd1;
	// controller for andOp_205.andOp_205_in0
	// controller for andOp_205.andOp_205_in1
	// Insensitive connections
	assign andOp_205_in0 = notOp_204_out;
	assign andOp_205_in1 = 1'd1;
	// controller for andOp_207.andOp_207_in0
	// controller for andOp_207.andOp_207_in1
	// Insensitive connections
	assign andOp_207_in0 = notOp_206_out;
	assign andOp_207_in1 = andOp_205_out;
	// controller for andOp_209.andOp_209_in0
	// controller for andOp_209.andOp_209_in1
	// Insensitive connections
	assign andOp_209_in0 = notOp_208_out;
	assign andOp_209_in1 = 1'd1;
	// controller for andOp_211.andOp_211_in0
	// controller for andOp_211.andOp_211_in1
	// Insensitive connections
	assign andOp_211_in0 = notOp_210_out;
	assign andOp_211_in1 = 1'd1;
	// controller for andOp_213.andOp_213_in0
	// controller for andOp_213.andOp_213_in1
	// Insensitive connections
	assign andOp_213_in0 = notOp_212_out;
	assign andOp_213_in1 = 1'd1;
	// controller for andOp_215.andOp_215_in0
	// controller for andOp_215.andOp_215_in1
	// Insensitive connections
	assign andOp_215_in0 = notOp_214_out;
	assign andOp_215_in1 = 1'd1;
	// controller for andOp_217.andOp_217_in0
	// controller for andOp_217.andOp_217_in1
	// Insensitive connections
	assign andOp_217_in0 = notOp_216_out;
	assign andOp_217_in1 = andOp_215_out;
	// controller for andOp_220.andOp_220_in0
	// controller for andOp_220.andOp_220_in1
	// Insensitive connections
	assign andOp_220_in0 = bb_2_active_in_state_0_out_data;
	assign andOp_220_in1 = state_0_is_active;
	// controller for andOp_221.andOp_221_in0
	// controller for andOp_221.andOp_221_in1
	// Insensitive connections
	assign andOp_221_in0 = bb_2_active_in_state_0_out_data;
	assign andOp_221_in1 = state_0_is_active;
	// controller for andOp_222.andOp_222_in0
	// controller for andOp_222.andOp_222_in1
	// Insensitive connections
	assign andOp_222_in0 = bb_2_active_in_state_0_out_data;
	assign andOp_222_in1 = state_0_is_active;
	// controller for andOp_230.andOp_230_in0
	// controller for andOp_230.andOp_230_in1
	// Insensitive connections
	assign andOp_230_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_230_in1 = state_3_is_active;
	// controller for andOp_231.andOp_231_in0
	// controller for andOp_231.andOp_231_in1
	// Insensitive connections
	assign andOp_231_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_231_in1 = state_3_is_active;
	// controller for andOp_240.andOp_240_in0
	// controller for andOp_240.andOp_240_in1
	// Insensitive connections
	assign andOp_240_in0 = bb_3_active_in_state_7_out_data;
	assign andOp_240_in1 = state_7_is_active;
	// controller for andOp_241.andOp_241_in0
	// controller for andOp_241.andOp_241_in1
	// Insensitive connections
	assign andOp_241_in0 = bb_2_active_in_state_0_out_data;
	assign andOp_241_in1 = state_0_is_active;
	// controller for andOp_242.andOp_242_in0
	// controller for andOp_242.andOp_242_in1
	// Insensitive connections
	assign andOp_242_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_242_in1 = state_3_is_active;
	// controller for andOp_243.andOp_243_in0
	// controller for andOp_243.andOp_243_in1
	// Insensitive connections
	assign andOp_243_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_243_in1 = state_3_is_active;
	// controller for andOp_244.andOp_244_in0
	// controller for andOp_244.andOp_244_in1
	// Insensitive connections
	assign andOp_244_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_244_in1 = state_3_is_active;
	// controller for andOp_245.andOp_245_in0
	// controller for andOp_245.andOp_245_in1
	// Insensitive connections
	assign andOp_245_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_245_in1 = state_4_is_active;
	// controller for andOp_246.andOp_246_in0
	// controller for andOp_246.andOp_246_in1
	// Insensitive connections
	assign andOp_246_in0 = bb_3_active_in_state_7_out_data;
	assign andOp_246_in1 = state_7_is_active;
	// controller for andOp_247.andOp_247_in0
	// controller for andOp_247.andOp_247_in1
	// Insensitive connections
	assign andOp_247_in0 = bb_2_active_in_state_0_out_data;
	assign andOp_247_in1 = state_0_is_active;
	// controller for andOp_248.andOp_248_in0
	// controller for andOp_248.andOp_248_in1
	// Insensitive connections
	assign andOp_248_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_248_in1 = state_4_is_active;
	// controller for andOp_249.andOp_249_in0
	// controller for andOp_249.andOp_249_in1
	// Insensitive connections
	assign andOp_249_in0 = bb_2_active_in_state_0_out_data;
	assign andOp_249_in1 = state_0_is_active;
	// controller for andOp_250.andOp_250_in0
	// controller for andOp_250.andOp_250_in1
	// Insensitive connections
	assign andOp_250_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_250_in1 = state_3_is_active;
	// controller for andOp_251.andOp_251_in0
	// controller for andOp_251.andOp_251_in1
	// Insensitive connections
	assign andOp_251_in0 = bb_2_active_in_state_0_out_data;
	assign andOp_251_in1 = state_0_is_active;
	// controller for andOp_252.andOp_252_in0
	// controller for andOp_252.andOp_252_in1
	// Insensitive connections
	assign andOp_252_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_252_in1 = state_4_is_active;
	// controller for andOp_253.andOp_253_in0
	// controller for andOp_253.andOp_253_in1
	// Insensitive connections
	assign andOp_253_in0 = bb_2_active_in_state_0_out_data;
	assign andOp_253_in1 = state_0_is_active;
	// controller for andOp_254.andOp_254_in0
	// controller for andOp_254.andOp_254_in1
	// Insensitive connections
	assign andOp_254_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_254_in1 = state_4_is_active;
	// controller for andOp_85.andOp_85_in0
	// controller for andOp_85.andOp_85_in1
	// Insensitive connections
	assign andOp_85_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_85_in1 = state_0_is_active;
	// controller for andOp_87.andOp_87_in0
	// controller for andOp_87.andOp_87_in1
	// Insensitive connections
	assign andOp_87_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_87_in1 = state_3_is_active;
	// controller for andOp_89.andOp_89_in0
	// controller for andOp_89.andOp_89_in1
	// Insensitive connections
	assign andOp_89_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_89_in1 = state_3_is_active;
	// controller for andOp_91.andOp_91_in0
	// controller for andOp_91.andOp_91_in1
	// Insensitive connections
	assign andOp_91_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_91_in1 = state_3_is_active;
	// controller for andOp_93.andOp_93_in0
	// controller for andOp_93.andOp_93_in1
	// Insensitive connections
	assign andOp_93_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_93_in1 = state_3_is_active;
	// controller for andOp_95.andOp_95_in0
	// controller for andOp_95.andOp_95_in1
	// Insensitive connections
	assign andOp_95_in0 = bb_4_active_in_state_7_out_data;
	assign andOp_95_in1 = state_7_is_active;
	// controller for andOp_97.andOp_97_in0
	// controller for andOp_97.andOp_97_in1
	// Insensitive connections
	assign andOp_97_in0 = andOp_95_out;
	assign andOp_97_in1 = data_in_7_84_out_data;
	// controller for andOp_99.andOp_99_in0
	// controller for andOp_99.andOp_99_in1
	// Insensitive connections
	assign andOp_99_in0 = andOp_95_out;
	assign andOp_99_in1 = notOp_98_out;
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_125_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_141_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_7.bb_1_active_in_state_7_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_7_in_data = orOp_137_out;
		end else begin
			bb_1_active_in_state_7_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_7.bb_1_predecessor_in_state_7_in_data
	always @(*) begin
		if (andOp_156_out) begin 
			bb_1_predecessor_in_state_7_in_data = 32'd3;
		end else if (eq_154_out) begin 
			bb_1_predecessor_in_state_7_in_data = state_7_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_7_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_0.bb_2_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_0_in_data = orOp_127_out;
		end else begin
			bb_2_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_1.bb_2_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_1_in_data = eq_128_out;
		end else begin
			bb_2_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_2.bb_2_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_2_in_data = eq_129_out;
		end else begin
			bb_2_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_3.bb_2_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_3_in_data = eq_130_out;
		end else begin
			bb_2_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_0.bb_2_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_144_out) begin 
			bb_2_predecessor_in_state_0_in_data = 32'd0;
		end else if (eq_142_out) begin 
			bb_2_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_1.bb_2_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_145_out) begin 
			bb_2_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_2.bb_2_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_146_out) begin 
			bb_2_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_3.bb_2_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_147_out) begin 
			bb_2_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_7.bb_3_active_in_state_7_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_7_in_data = orOp_139_out;
		end else begin
			bb_3_active_in_state_7_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_7.bb_3_predecessor_in_state_7_in_data
	always @(*) begin
		if (andOp_159_out) begin 
			bb_3_predecessor_in_state_7_in_data = 32'd4;
		end else if (eq_157_out) begin 
			bb_3_predecessor_in_state_7_in_data = state_7_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_7_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_3.bb_4_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_3_in_data = orOp_132_out;
		end else begin
			bb_4_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_4.bb_4_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_4_in_data = eq_133_out;
		end else begin
			bb_4_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_5.bb_4_active_in_state_5_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_5_in_data = eq_134_out;
		end else begin
			bb_4_active_in_state_5_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_6.bb_4_active_in_state_6_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_6_in_data = eq_135_out;
		end else begin
			bb_4_active_in_state_6_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_7.bb_4_active_in_state_7_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_7_in_data = eq_140_out;
		end else begin
			bb_4_active_in_state_7_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_3.bb_4_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_150_out) begin 
			bb_4_predecessor_in_state_3_in_data = 32'd2;
		end else if (eq_148_out) begin 
			bb_4_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_4.bb_4_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_151_out) begin 
			bb_4_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_5.bb_4_predecessor_in_state_5_in_data
	always @(*) begin
		if (eq_152_out) begin 
			bb_4_predecessor_in_state_5_in_data = state_5_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_5_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_6.bb_4_predecessor_in_state_6_in_data
	always @(*) begin
		if (eq_153_out) begin 
			bb_4_predecessor_in_state_6_in_data = state_6_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_6_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_7.bb_4_predecessor_in_state_7_in_data
	always @(*) begin
		if (eq_160_out) begin 
			bb_4_predecessor_in_state_7_in_data = state_7_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_7_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_85_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_86_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_2_happened_in_state_0.br_2_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_87_out) begin 
			br_2_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_88_out) begin 
			br_2_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_2_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_2_happened_in_state_1.br_2_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_89_out) begin 
			br_2_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_90_out) begin 
			br_2_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_2_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_2_happened_in_state_2.br_2_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_91_out) begin 
			br_2_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_92_out) begin 
			br_2_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_2_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_2_happened_in_state_3.br_2_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_93_out) begin 
			br_2_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_94_out) begin 
			br_2_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_2_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_7.br_3_happened_in_state_7_in_data
	always @(*) begin
		if (andOp_115_out) begin 
			br_3_happened_in_state_7_in_data = 1'd1;
		end else if (notOp_116_out) begin 
			br_3_happened_in_state_7_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_7_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_3.br_4_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_95_out) begin 
			br_4_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_96_out) begin 
			br_4_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_4.br_4_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_100_out) begin 
			br_4_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_101_out) begin 
			br_4_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_5.br_4_happened_in_state_5_in_data
	always @(*) begin
		if (andOp_105_out) begin 
			br_4_happened_in_state_5_in_data = 1'd1;
		end else if (notOp_106_out) begin 
			br_4_happened_in_state_5_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_5_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_6.br_4_happened_in_state_6_in_data
	always @(*) begin
		if (andOp_110_out) begin 
			br_4_happened_in_state_6_in_data = 1'd1;
		end else if (notOp_111_out) begin 
			br_4_happened_in_state_6_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_6_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_7.br_4_happened_in_state_7_in_data
	always @(*) begin
		if (andOp_120_out) begin 
			br_4_happened_in_state_7_in_data = 1'd1;
		end else if (notOp_121_out) begin 
			br_4_happened_in_state_7_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_7_in_data = 0;
		end
	end
	// controller for concat_162.concat_162_in0
	// controller for concat_162.concat_162_in1
	// Insensitive connections
	assign concat_162_in0 = data_in_0_4_out_data;
	assign concat_162_in1 = 32'd0;
	// controller for concat_163.concat_163_in0
	// controller for concat_163.concat_163_in1
	// Insensitive connections
	assign concat_163_in0 = 32'd3;
	assign concat_163_in1 = 32'd0;
	// controller for concat_179.concat_179_in0
	// controller for concat_179.concat_179_in1
	// Insensitive connections
	assign concat_179_in0 = data_in_3_36_out_data;
	assign concat_179_in1 = 32'd0;
	// controller for concat_180.concat_180_in0
	// controller for concat_180.concat_180_in1
	// Insensitive connections
	assign concat_180_in0 = 32'd4;
	assign concat_180_in1 = 32'd2;
	// controller for data_in_0_4.data_in_0_4_in_data
	always @(*) begin
		if (eq_218_out) begin 
			data_in_0_4_in_data = data_store_0_3;
		end else if (eq_219_out) begin 
			data_in_0_4_in_data = data_store_7_80;
		end else begin
			data_in_0_4_in_data = 0;
		end
	end
	// controller for data_in_0_6.data_in_0_6_in_data
	always @(*) begin
		if (eq_218_out) begin 
			data_in_0_6_in_data = data_store_0_5;
		end else if (eq_219_out) begin 
			data_in_0_6_in_data = data_store_7_82;
		end else begin
			data_in_0_6_in_data = 0;
		end
	end
	// controller for data_in_1_10.data_in_1_10_in_data
	always @(*) begin
		if (eq_223_out) begin 
			data_in_1_10_in_data = data_store_0_1;
		end else if (eq_224_out) begin 
			data_in_1_10_in_data = data_store_1_9;
		end else begin
			data_in_1_10_in_data = 0;
		end
	end
	// controller for data_in_1_12.data_in_1_12_in_data
	always @(*) begin
		if (eq_223_out) begin 
			data_in_1_12_in_data = data_store_0_2;
		end else if (eq_224_out) begin 
			data_in_1_12_in_data = data_store_1_11;
		end else begin
			data_in_1_12_in_data = 0;
		end
	end
	// controller for data_in_1_14.data_in_1_14_in_data
	always @(*) begin
		if (eq_223_out) begin 
			data_in_1_14_in_data = data_store_0_3;
		end else if (eq_224_out) begin 
			data_in_1_14_in_data = data_store_1_13;
		end else begin
			data_in_1_14_in_data = 0;
		end
	end
	// controller for data_in_1_16.data_in_1_16_in_data
	always @(*) begin
		if (eq_223_out) begin 
			data_in_1_16_in_data = data_store_0_5;
		end else if (eq_224_out) begin 
			data_in_1_16_in_data = data_store_1_15;
		end else begin
			data_in_1_16_in_data = 0;
		end
	end
	// controller for data_in_1_8.data_in_1_8_in_data
	always @(*) begin
		if (eq_223_out) begin 
			data_in_1_8_in_data = data_store_0_0;
		end else if (eq_224_out) begin 
			data_in_1_8_in_data = data_store_1_7;
		end else begin
			data_in_1_8_in_data = 0;
		end
	end
	// controller for data_in_2_18.data_in_2_18_in_data
	always @(*) begin
		if (eq_225_out) begin 
			data_in_2_18_in_data = data_store_1_7;
		end else if (eq_226_out) begin 
			data_in_2_18_in_data = data_store_2_17;
		end else begin
			data_in_2_18_in_data = 0;
		end
	end
	// controller for data_in_2_20.data_in_2_20_in_data
	always @(*) begin
		if (eq_225_out) begin 
			data_in_2_20_in_data = data_store_1_9;
		end else if (eq_226_out) begin 
			data_in_2_20_in_data = data_store_2_19;
		end else begin
			data_in_2_20_in_data = 0;
		end
	end
	// controller for data_in_2_22.data_in_2_22_in_data
	always @(*) begin
		if (eq_225_out) begin 
			data_in_2_22_in_data = data_store_1_11;
		end else if (eq_226_out) begin 
			data_in_2_22_in_data = data_store_2_21;
		end else begin
			data_in_2_22_in_data = 0;
		end
	end
	// controller for data_in_2_24.data_in_2_24_in_data
	always @(*) begin
		if (eq_225_out) begin 
			data_in_2_24_in_data = data_store_1_13;
		end else if (eq_226_out) begin 
			data_in_2_24_in_data = data_store_2_23;
		end else begin
			data_in_2_24_in_data = 0;
		end
	end
	// controller for data_in_2_26.data_in_2_26_in_data
	always @(*) begin
		if (eq_225_out) begin 
			data_in_2_26_in_data = data_store_1_15;
		end else if (eq_226_out) begin 
			data_in_2_26_in_data = data_store_2_25;
		end else begin
			data_in_2_26_in_data = 0;
		end
	end
	// controller for data_in_3_28.data_in_3_28_in_data
	always @(*) begin
		if (eq_227_out) begin 
			data_in_3_28_in_data = data_store_2_17;
		end else if (eq_228_out) begin 
			data_in_3_28_in_data = data_store_3_27;
		end else if (eq_229_out) begin 
			data_in_3_28_in_data = data_store_7_74;
		end else begin
			data_in_3_28_in_data = 0;
		end
	end
	// controller for data_in_3_30.data_in_3_30_in_data
	always @(*) begin
		if (eq_227_out) begin 
			data_in_3_30_in_data = data_store_2_19;
		end else if (eq_228_out) begin 
			data_in_3_30_in_data = data_store_3_29;
		end else if (eq_229_out) begin 
			data_in_3_30_in_data = data_store_7_76;
		end else begin
			data_in_3_30_in_data = 0;
		end
	end
	// controller for data_in_3_32.data_in_3_32_in_data
	always @(*) begin
		if (eq_227_out) begin 
			data_in_3_32_in_data = data_store_2_21;
		end else if (eq_228_out) begin 
			data_in_3_32_in_data = data_store_3_31;
		end else if (eq_229_out) begin 
			data_in_3_32_in_data = data_store_7_78;
		end else begin
			data_in_3_32_in_data = 0;
		end
	end
	// controller for data_in_3_34.data_in_3_34_in_data
	always @(*) begin
		if (eq_227_out) begin 
			data_in_3_34_in_data = data_store_2_23;
		end else if (eq_228_out) begin 
			data_in_3_34_in_data = data_store_3_33;
		end else if (eq_229_out) begin 
			data_in_3_34_in_data = data_store_7_80;
		end else begin
			data_in_3_34_in_data = 0;
		end
	end
	// controller for data_in_3_36.data_in_3_36_in_data
	always @(*) begin
		if (eq_227_out) begin 
			data_in_3_36_in_data = data_store_2_25;
		end else if (eq_228_out) begin 
			data_in_3_36_in_data = data_store_3_35;
		end else if (eq_229_out) begin 
			data_in_3_36_in_data = data_store_7_82;
		end else begin
			data_in_3_36_in_data = 0;
		end
	end
	// controller for data_in_4_39.data_in_4_39_in_data
	always @(*) begin
		if (eq_232_out) begin 
			data_in_4_39_in_data = data_store_3_27;
		end else if (eq_233_out) begin 
			data_in_4_39_in_data = data_store_4_38;
		end else begin
			data_in_4_39_in_data = 0;
		end
	end
	// controller for data_in_4_41.data_in_4_41_in_data
	always @(*) begin
		if (eq_232_out) begin 
			data_in_4_41_in_data = data_store_3_29;
		end else if (eq_233_out) begin 
			data_in_4_41_in_data = data_store_4_40;
		end else begin
			data_in_4_41_in_data = 0;
		end
	end
	// controller for data_in_4_43.data_in_4_43_in_data
	always @(*) begin
		if (eq_232_out) begin 
			data_in_4_43_in_data = data_store_3_31;
		end else if (eq_233_out) begin 
			data_in_4_43_in_data = data_store_4_42;
		end else begin
			data_in_4_43_in_data = 0;
		end
	end
	// controller for data_in_4_45.data_in_4_45_in_data
	always @(*) begin
		if (eq_232_out) begin 
			data_in_4_45_in_data = data_store_3_33;
		end else if (eq_233_out) begin 
			data_in_4_45_in_data = data_store_4_44;
		end else begin
			data_in_4_45_in_data = 0;
		end
	end
	// controller for data_in_4_47.data_in_4_47_in_data
	always @(*) begin
		if (eq_232_out) begin 
			data_in_4_47_in_data = data_store_3_35;
		end else if (eq_233_out) begin 
			data_in_4_47_in_data = data_store_4_46;
		end else begin
			data_in_4_47_in_data = 0;
		end
	end
	// controller for data_in_4_49.data_in_4_49_in_data
	always @(*) begin
		if (eq_232_out) begin 
			data_in_4_49_in_data = data_store_3_37;
		end else if (eq_233_out) begin 
			data_in_4_49_in_data = data_store_4_48;
		end else begin
			data_in_4_49_in_data = 0;
		end
	end
	// controller for data_in_5_51.data_in_5_51_in_data
	always @(*) begin
		if (eq_234_out) begin 
			data_in_5_51_in_data = data_store_4_38;
		end else if (eq_235_out) begin 
			data_in_5_51_in_data = data_store_5_50;
		end else begin
			data_in_5_51_in_data = 0;
		end
	end
	// controller for data_in_5_53.data_in_5_53_in_data
	always @(*) begin
		if (eq_234_out) begin 
			data_in_5_53_in_data = data_store_4_40;
		end else if (eq_235_out) begin 
			data_in_5_53_in_data = data_store_5_52;
		end else begin
			data_in_5_53_in_data = 0;
		end
	end
	// controller for data_in_5_55.data_in_5_55_in_data
	always @(*) begin
		if (eq_234_out) begin 
			data_in_5_55_in_data = data_store_4_42;
		end else if (eq_235_out) begin 
			data_in_5_55_in_data = data_store_5_54;
		end else begin
			data_in_5_55_in_data = 0;
		end
	end
	// controller for data_in_5_57.data_in_5_57_in_data
	always @(*) begin
		if (eq_234_out) begin 
			data_in_5_57_in_data = data_store_4_44;
		end else if (eq_235_out) begin 
			data_in_5_57_in_data = data_store_5_56;
		end else begin
			data_in_5_57_in_data = 0;
		end
	end
	// controller for data_in_5_59.data_in_5_59_in_data
	always @(*) begin
		if (eq_234_out) begin 
			data_in_5_59_in_data = data_store_4_46;
		end else if (eq_235_out) begin 
			data_in_5_59_in_data = data_store_5_58;
		end else begin
			data_in_5_59_in_data = 0;
		end
	end
	// controller for data_in_5_61.data_in_5_61_in_data
	always @(*) begin
		if (eq_234_out) begin 
			data_in_5_61_in_data = data_store_4_48;
		end else if (eq_235_out) begin 
			data_in_5_61_in_data = data_store_5_60;
		end else begin
			data_in_5_61_in_data = 0;
		end
	end
	// controller for data_in_6_63.data_in_6_63_in_data
	always @(*) begin
		if (eq_236_out) begin 
			data_in_6_63_in_data = data_store_5_50;
		end else if (eq_237_out) begin 
			data_in_6_63_in_data = data_store_6_62;
		end else begin
			data_in_6_63_in_data = 0;
		end
	end
	// controller for data_in_6_65.data_in_6_65_in_data
	always @(*) begin
		if (eq_236_out) begin 
			data_in_6_65_in_data = data_store_5_52;
		end else if (eq_237_out) begin 
			data_in_6_65_in_data = data_store_6_64;
		end else begin
			data_in_6_65_in_data = 0;
		end
	end
	// controller for data_in_6_67.data_in_6_67_in_data
	always @(*) begin
		if (eq_236_out) begin 
			data_in_6_67_in_data = data_store_5_54;
		end else if (eq_237_out) begin 
			data_in_6_67_in_data = data_store_6_66;
		end else begin
			data_in_6_67_in_data = 0;
		end
	end
	// controller for data_in_6_69.data_in_6_69_in_data
	always @(*) begin
		if (eq_236_out) begin 
			data_in_6_69_in_data = data_store_5_56;
		end else if (eq_237_out) begin 
			data_in_6_69_in_data = data_store_6_68;
		end else begin
			data_in_6_69_in_data = 0;
		end
	end
	// controller for data_in_6_71.data_in_6_71_in_data
	always @(*) begin
		if (eq_236_out) begin 
			data_in_6_71_in_data = data_store_5_58;
		end else if (eq_237_out) begin 
			data_in_6_71_in_data = data_store_6_70;
		end else begin
			data_in_6_71_in_data = 0;
		end
	end
	// controller for data_in_6_73.data_in_6_73_in_data
	always @(*) begin
		if (eq_236_out) begin 
			data_in_6_73_in_data = data_store_5_60;
		end else if (eq_237_out) begin 
			data_in_6_73_in_data = data_store_6_72;
		end else begin
			data_in_6_73_in_data = 0;
		end
	end
	// controller for data_in_7_75.data_in_7_75_in_data
	always @(*) begin
		if (eq_238_out) begin 
			data_in_7_75_in_data = data_store_6_62;
		end else if (eq_239_out) begin 
			data_in_7_75_in_data = data_store_7_74;
		end else begin
			data_in_7_75_in_data = 0;
		end
	end
	// controller for data_in_7_77.data_in_7_77_in_data
	always @(*) begin
		if (eq_238_out) begin 
			data_in_7_77_in_data = data_store_6_64;
		end else if (eq_239_out) begin 
			data_in_7_77_in_data = data_store_7_76;
		end else begin
			data_in_7_77_in_data = 0;
		end
	end
	// controller for data_in_7_79.data_in_7_79_in_data
	always @(*) begin
		if (eq_238_out) begin 
			data_in_7_79_in_data = data_store_6_66;
		end else if (eq_239_out) begin 
			data_in_7_79_in_data = data_store_7_78;
		end else begin
			data_in_7_79_in_data = 0;
		end
	end
	// controller for data_in_7_81.data_in_7_81_in_data
	always @(*) begin
		if (eq_238_out) begin 
			data_in_7_81_in_data = data_store_6_68;
		end else if (eq_239_out) begin 
			data_in_7_81_in_data = data_store_7_80;
		end else begin
			data_in_7_81_in_data = 0;
		end
	end
	// controller for data_in_7_83.data_in_7_83_in_data
	always @(*) begin
		if (eq_238_out) begin 
			data_in_7_83_in_data = data_store_6_70;
		end else if (eq_239_out) begin 
			data_in_7_83_in_data = data_store_7_82;
		end else begin
			data_in_7_83_in_data = 0;
		end
	end
	// controller for data_in_7_84.data_in_7_84_in_data
	always @(*) begin
		if (eq_238_out) begin 
			data_in_7_84_in_data = data_store_6_72;
		end else if (eq_239_out) begin 
			data_in_7_84_in_data = 1'd0;
		end else begin
			data_in_7_84_in_data = 0;
		end
	end
	// controller for eq_125.eq_125_in0
	// controller for eq_125.eq_125_in1
	// Insensitive connections
	assign eq_125_in0 = 32'd0;
	assign eq_125_in1 = state_0_entry_BB_reg;
	// controller for eq_126.eq_126_in0
	// controller for eq_126.eq_126_in1
	// Insensitive connections
	assign eq_126_in0 = 32'd2;
	assign eq_126_in1 = state_0_entry_BB_reg;
	// controller for eq_128.eq_128_in0
	// controller for eq_128.eq_128_in1
	// Insensitive connections
	assign eq_128_in0 = 32'd2;
	assign eq_128_in1 = state_1_entry_BB_reg;
	// controller for eq_129.eq_129_in0
	// controller for eq_129.eq_129_in1
	// Insensitive connections
	assign eq_129_in0 = 32'd2;
	assign eq_129_in1 = state_2_entry_BB_reg;
	// controller for eq_130.eq_130_in0
	// controller for eq_130.eq_130_in1
	// Insensitive connections
	assign eq_130_in0 = 32'd2;
	assign eq_130_in1 = state_3_entry_BB_reg;
	// controller for eq_131.eq_131_in0
	// controller for eq_131.eq_131_in1
	// Insensitive connections
	assign eq_131_in0 = 32'd4;
	assign eq_131_in1 = state_3_entry_BB_reg;
	// controller for eq_133.eq_133_in0
	// controller for eq_133.eq_133_in1
	// Insensitive connections
	assign eq_133_in0 = 32'd4;
	assign eq_133_in1 = state_4_entry_BB_reg;
	// controller for eq_134.eq_134_in0
	// controller for eq_134.eq_134_in1
	// Insensitive connections
	assign eq_134_in0 = 32'd4;
	assign eq_134_in1 = state_5_entry_BB_reg;
	// controller for eq_135.eq_135_in0
	// controller for eq_135.eq_135_in1
	// Insensitive connections
	assign eq_135_in0 = 32'd4;
	assign eq_135_in1 = state_6_entry_BB_reg;
	// controller for eq_136.eq_136_in0
	// controller for eq_136.eq_136_in1
	// Insensitive connections
	assign eq_136_in0 = 32'd1;
	assign eq_136_in1 = state_7_entry_BB_reg;
	// controller for eq_138.eq_138_in0
	// controller for eq_138.eq_138_in1
	// Insensitive connections
	assign eq_138_in0 = 32'd3;
	assign eq_138_in1 = state_7_entry_BB_reg;
	// controller for eq_140.eq_140_in0
	// controller for eq_140.eq_140_in1
	// Insensitive connections
	assign eq_140_in0 = 32'd4;
	assign eq_140_in1 = state_7_entry_BB_reg;
	// controller for eq_141.eq_141_in0
	// controller for eq_141.eq_141_in1
	// Insensitive connections
	assign eq_141_in0 = 32'd0;
	assign eq_141_in1 = state_0_entry_BB_reg;
	// controller for eq_142.eq_142_in0
	// controller for eq_142.eq_142_in1
	// Insensitive connections
	assign eq_142_in0 = 32'd2;
	assign eq_142_in1 = state_0_entry_BB_reg;
	// controller for eq_145.eq_145_in0
	// controller for eq_145.eq_145_in1
	// Insensitive connections
	assign eq_145_in0 = 32'd2;
	assign eq_145_in1 = state_1_entry_BB_reg;
	// controller for eq_146.eq_146_in0
	// controller for eq_146.eq_146_in1
	// Insensitive connections
	assign eq_146_in0 = 32'd2;
	assign eq_146_in1 = state_2_entry_BB_reg;
	// controller for eq_147.eq_147_in0
	// controller for eq_147.eq_147_in1
	// Insensitive connections
	assign eq_147_in0 = 32'd2;
	assign eq_147_in1 = state_3_entry_BB_reg;
	// controller for eq_148.eq_148_in0
	// controller for eq_148.eq_148_in1
	// Insensitive connections
	assign eq_148_in0 = 32'd4;
	assign eq_148_in1 = state_3_entry_BB_reg;
	// controller for eq_151.eq_151_in0
	// controller for eq_151.eq_151_in1
	// Insensitive connections
	assign eq_151_in0 = 32'd4;
	assign eq_151_in1 = state_4_entry_BB_reg;
	// controller for eq_152.eq_152_in0
	// controller for eq_152.eq_152_in1
	// Insensitive connections
	assign eq_152_in0 = 32'd4;
	assign eq_152_in1 = state_5_entry_BB_reg;
	// controller for eq_153.eq_153_in0
	// controller for eq_153.eq_153_in1
	// Insensitive connections
	assign eq_153_in0 = 32'd4;
	assign eq_153_in1 = state_6_entry_BB_reg;
	// controller for eq_154.eq_154_in0
	// controller for eq_154.eq_154_in1
	// Insensitive connections
	assign eq_154_in0 = 32'd1;
	assign eq_154_in1 = state_7_entry_BB_reg;
	// controller for eq_157.eq_157_in0
	// controller for eq_157.eq_157_in1
	// Insensitive connections
	assign eq_157_in0 = 32'd3;
	assign eq_157_in1 = state_7_entry_BB_reg;
	// controller for eq_160.eq_160_in0
	// controller for eq_160.eq_160_in1
	// Insensitive connections
	assign eq_160_in0 = 32'd4;
	assign eq_160_in1 = state_7_entry_BB_reg;
	// controller for eq_218.eq_218_in0
	// controller for eq_218.eq_218_in1
	// Insensitive connections
	assign eq_218_in0 = 32'd0;
	assign eq_218_in1 = state_0_last_state;
	// controller for eq_219.eq_219_in0
	// controller for eq_219.eq_219_in1
	// Insensitive connections
	assign eq_219_in0 = 32'd7;
	assign eq_219_in1 = state_0_last_state;
	// controller for eq_223.eq_223_in0
	// controller for eq_223.eq_223_in1
	// Insensitive connections
	assign eq_223_in0 = 32'd0;
	assign eq_223_in1 = state_1_last_state;
	// controller for eq_224.eq_224_in0
	// controller for eq_224.eq_224_in1
	// Insensitive connections
	assign eq_224_in0 = 32'd1;
	assign eq_224_in1 = state_1_last_state;
	// controller for eq_225.eq_225_in0
	// controller for eq_225.eq_225_in1
	// Insensitive connections
	assign eq_225_in0 = 32'd1;
	assign eq_225_in1 = state_2_last_state;
	// controller for eq_226.eq_226_in0
	// controller for eq_226.eq_226_in1
	// Insensitive connections
	assign eq_226_in0 = 32'd2;
	assign eq_226_in1 = state_2_last_state;
	// controller for eq_227.eq_227_in0
	// controller for eq_227.eq_227_in1
	// Insensitive connections
	assign eq_227_in0 = 32'd2;
	assign eq_227_in1 = state_3_last_state;
	// controller for eq_228.eq_228_in0
	// controller for eq_228.eq_228_in1
	// Insensitive connections
	assign eq_228_in0 = 32'd3;
	assign eq_228_in1 = state_3_last_state;
	// controller for eq_229.eq_229_in0
	// controller for eq_229.eq_229_in1
	// Insensitive connections
	assign eq_229_in0 = 32'd7;
	assign eq_229_in1 = state_3_last_state;
	// controller for eq_232.eq_232_in0
	// controller for eq_232.eq_232_in1
	// Insensitive connections
	assign eq_232_in0 = 32'd3;
	assign eq_232_in1 = state_4_last_state;
	// controller for eq_233.eq_233_in0
	// controller for eq_233.eq_233_in1
	// Insensitive connections
	assign eq_233_in0 = 32'd4;
	assign eq_233_in1 = state_4_last_state;
	// controller for eq_234.eq_234_in0
	// controller for eq_234.eq_234_in1
	// Insensitive connections
	assign eq_234_in0 = 32'd4;
	assign eq_234_in1 = state_5_last_state;
	// controller for eq_235.eq_235_in0
	// controller for eq_235.eq_235_in1
	// Insensitive connections
	assign eq_235_in0 = 32'd5;
	assign eq_235_in1 = state_5_last_state;
	// controller for eq_236.eq_236_in0
	// controller for eq_236.eq_236_in1
	// Insensitive connections
	assign eq_236_in0 = 32'd5;
	assign eq_236_in1 = state_6_last_state;
	// controller for eq_237.eq_237_in0
	// controller for eq_237.eq_237_in1
	// Insensitive connections
	assign eq_237_in0 = 32'd6;
	assign eq_237_in1 = state_6_last_state;
	// controller for eq_238.eq_238_in0
	// controller for eq_238.eq_238_in1
	// Insensitive connections
	assign eq_238_in0 = 32'd6;
	assign eq_238_in1 = state_7_last_state;
	// controller for eq_239.eq_239_in0
	// controller for eq_239.eq_239_in1
	// Insensitive connections
	assign eq_239_in0 = 32'd7;
	assign eq_239_in1 = state_7_last_state;
	// controller for icmp_icmp12.icmp_icmp12_in0
	// controller for icmp_icmp12.icmp_icmp12_in1
	// Insensitive connections
	assign icmp_icmp12_in0 = add_add11_out;
	assign icmp_icmp12_in1 = 32'd3;
	// controller for icmp_icmp26.icmp_icmp26_in0
	// controller for icmp_icmp26.icmp_icmp26_in1
	// Insensitive connections
	assign icmp_icmp26_in0 = add_add25_out;
	assign icmp_icmp26_in1 = 32'd3;
	// controller for mul_mul16.mul_mul16_in0
	// controller for mul_mul16.mul_mul16_in1
	// Insensitive connections
	assign mul_mul16_in0 = ram_rdata_2;
	assign mul_mul16_in1 = ram_rdata_1;
	// controller for mul_mul3.mul_mul3_in0
	// controller for mul_mul3.mul_mul3_in1
	// Insensitive connections
	assign mul_mul3_in0 = phi_phi1_out;
	assign mul_mul3_in1 = 32'd3;
	// controller for notOp_101.notOp_101_in0
	// Insensitive connections
	assign notOp_101_in0 = andOp_100_out;
	// controller for notOp_103.notOp_103_in0
	// Insensitive connections
	assign notOp_103_in0 = data_in_7_84_out_data;
	// controller for notOp_106.notOp_106_in0
	// Insensitive connections
	assign notOp_106_in0 = andOp_105_out;
	// controller for notOp_108.notOp_108_in0
	// Insensitive connections
	assign notOp_108_in0 = data_in_7_84_out_data;
	// controller for notOp_111.notOp_111_in0
	// Insensitive connections
	assign notOp_111_in0 = andOp_110_out;
	// controller for notOp_113.notOp_113_in0
	// Insensitive connections
	assign notOp_113_in0 = data_in_7_84_out_data;
	// controller for notOp_116.notOp_116_in0
	// Insensitive connections
	assign notOp_116_in0 = andOp_115_out;
	// controller for notOp_118.notOp_118_in0
	// Insensitive connections
	assign notOp_118_in0 = icmp_icmp26_out;
	// controller for notOp_121.notOp_121_in0
	// Insensitive connections
	assign notOp_121_in0 = andOp_120_out;
	// controller for notOp_123.notOp_123_in0
	// Insensitive connections
	assign notOp_123_in0 = data_in_7_84_out_data;
	// controller for notOp_143.notOp_143_in0
	// Insensitive connections
	assign notOp_143_in0 = eq_142_out;
	// controller for notOp_149.notOp_149_in0
	// Insensitive connections
	assign notOp_149_in0 = eq_148_out;
	// controller for notOp_155.notOp_155_in0
	// Insensitive connections
	assign notOp_155_in0 = eq_154_out;
	// controller for notOp_158.notOp_158_in0
	// Insensitive connections
	assign notOp_158_in0 = eq_157_out;
	// controller for notOp_198.notOp_198_in0
	// Insensitive connections
	assign notOp_198_in0 = andOp_119_out;
	// controller for notOp_200.notOp_200_in0
	// Insensitive connections
	assign notOp_200_in0 = andOp_190_out;
	// controller for notOp_202.notOp_202_in0
	// Insensitive connections
	assign notOp_202_in0 = andOp_191_out;
	// controller for notOp_204.notOp_204_in0
	// Insensitive connections
	assign notOp_204_in0 = andOp_192_out;
	// controller for notOp_206.notOp_206_in0
	// Insensitive connections
	assign notOp_206_in0 = andOp_99_out;
	// controller for notOp_208.notOp_208_in0
	// Insensitive connections
	assign notOp_208_in0 = andOp_193_out;
	// controller for notOp_210.notOp_210_in0
	// Insensitive connections
	assign notOp_210_in0 = andOp_194_out;
	// controller for notOp_212.notOp_212_in0
	// Insensitive connections
	assign notOp_212_in0 = andOp_195_out;
	// controller for notOp_214.notOp_214_in0
	// Insensitive connections
	assign notOp_214_in0 = andOp_196_out;
	// controller for notOp_216.notOp_216_in0
	// Insensitive connections
	assign notOp_216_in0 = andOp_197_out;
	// controller for notOp_86.notOp_86_in0
	// Insensitive connections
	assign notOp_86_in0 = andOp_85_out;
	// controller for notOp_88.notOp_88_in0
	// Insensitive connections
	assign notOp_88_in0 = andOp_87_out;
	// controller for notOp_90.notOp_90_in0
	// Insensitive connections
	assign notOp_90_in0 = andOp_89_out;
	// controller for notOp_92.notOp_92_in0
	// Insensitive connections
	assign notOp_92_in0 = andOp_91_out;
	// controller for notOp_94.notOp_94_in0
	// Insensitive connections
	assign notOp_94_in0 = andOp_93_out;
	// controller for notOp_96.notOp_96_in0
	// Insensitive connections
	assign notOp_96_in0 = andOp_95_out;
	// controller for notOp_98.notOp_98_in0
	// Insensitive connections
	assign notOp_98_in0 = data_in_7_84_out_data;
	// controller for orOp_127.orOp_127_in0
	// controller for orOp_127.orOp_127_in1
	// Insensitive connections
	assign orOp_127_in0 = eq_126_out;
	assign orOp_127_in1 = andOp_85_out;
	// controller for orOp_132.orOp_132_in0
	// controller for orOp_132.orOp_132_in1
	// Insensitive connections
	assign orOp_132_in0 = eq_131_out;
	assign orOp_132_in1 = andOp_87_out;
	// controller for orOp_137.orOp_137_in0
	// controller for orOp_137.orOp_137_in1
	// Insensitive connections
	assign orOp_137_in0 = eq_136_out;
	assign orOp_137_in1 = andOp_117_out;
	// controller for orOp_139.orOp_139_in0
	// controller for orOp_139.orOp_139_in1
	// Insensitive connections
	assign orOp_139_in0 = eq_138_out;
	assign orOp_139_in1 = andOp_97_out;
	// controller for phi_phi1.phi_phi1_in
	// controller for phi_phi1.phi_phi1_last_block
	// controller for phi_phi1.phi_phi1_s
	// Insensitive connections
	assign phi_phi1_in = concat_162_out;
	assign phi_phi1_last_block = bb_2_predecessor_in_state_0_out_data;
	assign phi_phi1_s = concat_163_out;
	// controller for phi_phi7.phi_phi7_in
	// controller for phi_phi7.phi_phi7_last_block
	// controller for phi_phi7.phi_phi7_s
	// Insensitive connections
	assign phi_phi7_in = concat_179_out;
	assign phi_phi7_last_block = bb_4_predecessor_in_state_3_out_data;
	assign phi_phi7_s = concat_180_out;
	// controller for ram.ram_raddr_0_reg
	always @(*) begin
		if (andOp_170_out) begin 
			ram_raddr_0_reg = data_in_3_30_out_data;
		end else begin
			ram_raddr_0_reg = 0;
		end
	end
	// controller for ram.ram_raddr_1_reg
	always @(*) begin
		if (andOp_171_out) begin 
			ram_raddr_1_reg = add_add9_out;
		end else begin
			ram_raddr_1_reg = 0;
		end
	end
	// controller for ram.ram_raddr_2_reg
	always @(*) begin
		if (andOp_169_out) begin 
			ram_raddr_2_reg = add_add10_out;
		end else begin
			ram_raddr_2_reg = 0;
		end
	end
	// controller for ram.ram_waddr_0_reg
	always @(*) begin
		if (andOp_166_out) begin 
			ram_waddr_0_reg = add_add2_out;
		end else if (andOp_175_out) begin 
			ram_waddr_0_reg = data_in_4_41_out_data;
		end else begin
			ram_waddr_0_reg = 0;
		end
	end
	// controller for ram.ram_wdata_0_reg
	always @(*) begin
		if (andOp_167_out) begin 
			ram_wdata_0_reg = 32'd0;
		end else if (andOp_176_out) begin 
			ram_wdata_0_reg = add_add17_out;
		end else begin
			ram_wdata_0_reg = 0;
		end
	end
	// controller for ram.ram_wen_0_reg
	always @(*) begin
		if (andOp_168_out) begin 
			ram_wen_0_reg = -(1'd1);
		end else if (andOp_177_out) begin 
			ram_wen_0_reg = -(1'd1);
		end else begin
			ram_wen_0_reg = 0;
		end
	end
	// controller for ret24.valid_reg
	always @(*) begin
		if (andOp_187_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			data_store_0_0 <= 0;
		end else begin
			if (andOp_220_out) begin
				data_store_0_0 <= phi_phi1_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_1 <= 0;
		end else begin
			if (andOp_221_out) begin
				data_store_0_1 <= add_add2_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_2 <= 0;
		end else begin
			if (andOp_222_out) begin
				data_store_0_2 <= mul_mul3_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_3 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_3 <= data_in_0_4_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_5 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_5 <= data_in_0_6_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_11 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_11 <= data_in_1_12_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_13 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_13 <= data_in_1_14_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_15 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_15 <= data_in_1_16_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_7 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_7 <= data_in_1_8_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_9 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_9 <= data_in_1_10_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_17 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_17 <= data_in_2_18_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_19 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_19 <= data_in_2_20_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_21 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_21 <= data_in_2_22_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_23 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_23 <= data_in_2_24_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_25 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_25 <= data_in_2_26_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_27 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_27 <= data_in_3_28_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_29 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_29 <= data_in_3_30_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_31 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_31 <= data_in_3_32_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_33 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_33 <= data_in_3_34_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_35 <= 0;
		end else begin
			if (andOp_230_out) begin
				data_store_3_35 <= add_add11_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_37 <= 0;
		end else begin
			if (andOp_231_out) begin
				data_store_3_37 <= icmp_icmp12_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_38 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_38 <= data_in_4_39_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_40 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_40 <= data_in_4_41_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_42 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_42 <= data_in_4_43_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_44 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_44 <= data_in_4_45_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_46 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_46 <= data_in_4_47_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_48 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_48 <= data_in_4_49_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_50 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_50 <= data_in_5_51_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_52 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_52 <= data_in_5_53_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_54 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_54 <= data_in_5_55_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_56 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_56 <= data_in_5_57_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_58 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_58 <= data_in_5_59_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_60 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_60 <= data_in_5_61_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_62 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_62 <= data_in_6_63_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_64 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_64 <= data_in_6_65_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_66 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_66 <= data_in_6_67_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_68 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_68 <= data_in_6_69_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_70 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_70 <= data_in_6_71_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_72 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_72 <= data_in_6_73_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_7_74 <= 0;
		end else begin
			if (state_7_is_active) begin
				data_store_7_74 <= data_in_7_75_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_7_76 <= 0;
		end else begin
			if (state_7_is_active) begin
				data_store_7_76 <= data_in_7_77_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_7_78 <= 0;
		end else begin
			if (state_7_is_active) begin
				data_store_7_78 <= data_in_7_79_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_7_80 <= 0;
		end else begin
			if (andOp_240_out) begin
				data_store_7_80 <= add_add25_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_7_82 <= 0;
		end else begin
			if (state_7_is_active) begin
				data_store_7_82 <= data_in_7_83_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_119_out) begin
				global_state <= 32'd0;
			end
			if (andOp_190_out) begin
				global_state <= 32'd1;
			end
			if (andOp_191_out) begin
				global_state <= 32'd2;
			end
			if (andOp_192_out) begin
				global_state <= 32'd3;
			end
			if (andOp_193_out) begin
				global_state <= 32'd4;
			end
			if (andOp_194_out) begin
				global_state <= 32'd5;
			end
			if (andOp_195_out) begin
				global_state <= 32'd6;
			end
			if (andOp_196_out) begin
				global_state <= 32'd7;
			end
			if (andOp_197_out) begin
				global_state <= 32'd7;
			end
			if (andOp_99_out) begin
				global_state <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
			if (andOp_119_out) begin
				state_0_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (andOp_119_out) begin
				state_0_is_active <= 1'd1;
			end
			if (andOp_199_out) begin
				state_0_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
			if (andOp_119_out) begin
				state_0_last_BB_reg <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
			if (andOp_119_out) begin
				state_0_last_state <= 32'd7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_190_out) begin
				state_1_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_190_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_201_out) begin
				state_1_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_190_out) begin
				state_1_last_BB_reg <= bb_2_predecessor_in_state_0_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_190_out) begin
				state_1_last_state <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_191_out) begin
				state_2_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_191_out) begin
				state_2_is_active <= 1'd1;
			end
			if (andOp_203_out) begin
				state_2_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_191_out) begin
				state_2_last_BB_reg <= bb_2_predecessor_in_state_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_191_out) begin
				state_2_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_192_out) begin
				state_3_entry_BB_reg <= 32'd2;
			end
			if (andOp_99_out) begin
				state_3_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_192_out) begin
				state_3_is_active <= 1'd1;
			end
			if (andOp_207_out) begin
				state_3_is_active <= 1'd0;
			end
			if (andOp_99_out) begin
				state_3_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_192_out) begin
				state_3_last_BB_reg <= bb_2_predecessor_in_state_2_out_data;
			end
			if (andOp_99_out) begin
				state_3_last_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_state <= 0;
		end else begin
			if (andOp_192_out) begin
				state_3_last_state <= 32'd2;
			end
			if (andOp_99_out) begin
				state_3_last_state <= 32'd7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_193_out) begin
				state_4_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_193_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_209_out) begin
				state_4_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_193_out) begin
				state_4_last_BB_reg <= bb_4_predecessor_in_state_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_state <= 0;
		end else begin
			if (andOp_193_out) begin
				state_4_last_state <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_entry_BB_reg <= 0;
		end else begin
			if (andOp_194_out) begin
				state_5_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_is_active <= 0;
		end else begin
			if (andOp_194_out) begin
				state_5_is_active <= 1'd1;
			end
			if (andOp_211_out) begin
				state_5_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_last_BB_reg <= 0;
		end else begin
			if (andOp_194_out) begin
				state_5_last_BB_reg <= bb_4_predecessor_in_state_4_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_last_state <= 0;
		end else begin
			if (andOp_194_out) begin
				state_5_last_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_entry_BB_reg <= 0;
		end else begin
			if (andOp_195_out) begin
				state_6_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_is_active <= 0;
		end else begin
			if (andOp_195_out) begin
				state_6_is_active <= 1'd1;
			end
			if (andOp_213_out) begin
				state_6_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_last_BB_reg <= 0;
		end else begin
			if (andOp_195_out) begin
				state_6_last_BB_reg <= bb_4_predecessor_in_state_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_last_state <= 0;
		end else begin
			if (andOp_195_out) begin
				state_6_last_state <= 32'd5;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_entry_BB_reg <= 0;
		end else begin
			if (andOp_196_out) begin
				state_7_entry_BB_reg <= 32'd4;
			end
			if (andOp_197_out) begin
				state_7_entry_BB_reg <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_is_active <= 0;
		end else begin
			if (andOp_196_out) begin
				state_7_is_active <= 1'd1;
			end
			if (andOp_197_out) begin
				state_7_is_active <= 1'd1;
			end
			if (andOp_217_out) begin
				state_7_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_last_BB_reg <= 0;
		end else begin
			if (andOp_196_out) begin
				state_7_last_BB_reg <= bb_4_predecessor_in_state_6_out_data;
			end
			if (andOp_197_out) begin
				state_7_last_BB_reg <= bb_1_predecessor_in_state_7_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_last_state <= 0;
		end else begin
			if (andOp_196_out) begin
				state_7_last_state <= 32'd6;
			end
			if (andOp_197_out) begin
				state_7_last_state <= 32'd7;
			end
		end
	end

endmodule

