module median_filter(input [0:0] clk, input [0:0] rst, output [0:0] valid, output [31:0] in0_in_data, input [31:0] in0_out_data, output [31:0] in1_in_data, input [31:0] in1_out_data, output [31:0] in2_in_data, input [31:0] in2_out_data, output [31:0] out_in_data, input [31:0] out_out_data);

	reg [0:0] valid_reg;
	reg [31:0] in0_in_data_reg;
	reg [31:0] in1_in_data_reg;
	reg [31:0] in2_in_data_reg;
	reg [31:0] out_in_data_reg;

	assign valid = valid_reg;
	assign in0_in_data = in0_in_data_reg;
	assign in1_in_data = in1_in_data_reg;
	assign in2_in_data = in2_in_data_reg;
	assign out_in_data = out_in_data_reg;

	// Start debug wires and ports

	initial begin
	end





	// End debug wires and ports

	// Start Functional Units
	reg [0:0] m_rst_n;
	reg [31:0] m_word0;
	reg [31:0] m_word1;
	reg [31:0] m_word2;
	wire [31:0] m_median_word;
	median m(.clk(clk), .median_word(m_median_word), .rst_n(m_rst_n), .word0(m_word0), .word1(m_word1), .word2(m_word2));

	br_dummy br_unit();

	reg [63:0] phi_in_phi_8;
	reg [31:0] phi_last_block_phi_8;
	reg [63:0] phi_s_phi_8;
	wire [31:0] phi_out_phi_8;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_8(.in(phi_in_phi_8), .last_block(phi_last_block_phi_8), .out(phi_out_phi_8), .s(phi_s_phi_8));

	reg [31:0] add_in0_add_9;
	reg [31:0] add_in1_add_9;
	wire [31:0] add_out_add_9;
	add #(.WIDTH(32)) add_add_9(.in0(add_in0_add_9), .in1(add_in1_add_9), .out(add_out_add_9));

	reg [31:0] cmp_in0_icmp_18;
	reg [31:0] cmp_in1_icmp_18;
	wire [0:0] cmp_out_icmp_18;
	ne #(.WIDTH(32)) icmp_18(.in0(cmp_in0_icmp_18), .in1(cmp_in1_icmp_18), .out(cmp_out_icmp_18));

	reg [31:0] data_in_0_1_in_data;
	wire [31:0] data_in_0_1_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_1(.in_data(data_in_0_1_in_data), .out_data(data_in_0_1_out_data));

	reg [31:0] data_in_0_3_in_data;
	wire [31:0] data_in_0_3_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_3(.in_data(data_in_0_3_in_data), .out_data(data_in_0_3_out_data));

	reg [31:0] data_in_0_5_in_data;
	wire [31:0] data_in_0_5_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_5(.in_data(data_in_0_5_in_data), .out_data(data_in_0_5_out_data));

	reg [31:0] data_in_0_7_in_data;
	wire [31:0] data_in_0_7_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_7(.in_data(data_in_0_7_in_data), .out_data(data_in_0_7_out_data));

	reg [31:0] data_in_0_9_in_data;
	wire [31:0] data_in_0_9_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_9(.in_data(data_in_0_9_in_data), .out_data(data_in_0_9_out_data));

	reg [31:0] data_in_0_11_in_data;
	wire [31:0] data_in_0_11_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_11(.in_data(data_in_0_11_in_data), .out_data(data_in_0_11_out_data));

	reg [0:0] data_in_0_13_in_data;
	wire [0:0] data_in_0_13_out_data;
	hls_wire #(.WIDTH(1)) data_in_0_13(.in_data(data_in_0_13_in_data), .out_data(data_in_0_13_out_data));

	reg [31:0] data_in_1_15_in_data;
	wire [31:0] data_in_1_15_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_15(.in_data(data_in_1_15_in_data), .out_data(data_in_1_15_out_data));

	reg [31:0] data_in_1_17_in_data;
	wire [31:0] data_in_1_17_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_17(.in_data(data_in_1_17_in_data), .out_data(data_in_1_17_out_data));

	reg [31:0] data_in_1_19_in_data;
	wire [31:0] data_in_1_19_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_19(.in_data(data_in_1_19_in_data), .out_data(data_in_1_19_out_data));

	reg [31:0] data_in_1_21_in_data;
	wire [31:0] data_in_1_21_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_21(.in_data(data_in_1_21_in_data), .out_data(data_in_1_21_out_data));

	reg [31:0] data_in_1_23_in_data;
	wire [31:0] data_in_1_23_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_23(.in_data(data_in_1_23_in_data), .out_data(data_in_1_23_out_data));

	reg [31:0] data_in_1_25_in_data;
	wire [31:0] data_in_1_25_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_25(.in_data(data_in_1_25_in_data), .out_data(data_in_1_25_out_data));

	reg [0:0] data_in_1_27_in_data;
	wire [0:0] data_in_1_27_out_data;
	hls_wire #(.WIDTH(1)) data_in_1_27(.in_data(data_in_1_27_in_data), .out_data(data_in_1_27_out_data));

	reg [31:0] data_in_2_29_in_data;
	wire [31:0] data_in_2_29_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_29(.in_data(data_in_2_29_in_data), .out_data(data_in_2_29_out_data));

	reg [31:0] data_in_2_31_in_data;
	wire [31:0] data_in_2_31_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_31(.in_data(data_in_2_31_in_data), .out_data(data_in_2_31_out_data));

	reg [31:0] data_in_2_33_in_data;
	wire [31:0] data_in_2_33_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_33(.in_data(data_in_2_33_in_data), .out_data(data_in_2_33_out_data));

	reg [31:0] data_in_2_35_in_data;
	wire [31:0] data_in_2_35_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_35(.in_data(data_in_2_35_in_data), .out_data(data_in_2_35_out_data));

	reg [31:0] data_in_2_37_in_data;
	wire [31:0] data_in_2_37_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_37(.in_data(data_in_2_37_in_data), .out_data(data_in_2_37_out_data));

	reg [31:0] data_in_2_39_in_data;
	wire [31:0] data_in_2_39_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_39(.in_data(data_in_2_39_in_data), .out_data(data_in_2_39_out_data));

	reg [0:0] data_in_2_41_in_data;
	wire [0:0] data_in_2_41_out_data;
	hls_wire #(.WIDTH(1)) data_in_2_41(.in_data(data_in_2_41_in_data), .out_data(data_in_2_41_out_data));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] bb_2_active_in_state_0_in_data;
	wire [0:0] bb_2_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_0(.in_data(bb_2_active_in_state_0_in_data), .out_data(bb_2_active_in_state_0_out_data));

	reg [31:0] bb_2_predecessor_in_state_0_in_data;
	wire [31:0] bb_2_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_0(.in_data(bb_2_predecessor_in_state_0_in_data), .out_data(bb_2_predecessor_in_state_0_out_data));

	reg [0:0] bb_2_active_in_state_1_in_data;
	wire [0:0] bb_2_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_1(.in_data(bb_2_active_in_state_1_in_data), .out_data(bb_2_active_in_state_1_out_data));

	reg [31:0] bb_2_predecessor_in_state_1_in_data;
	wire [31:0] bb_2_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_1(.in_data(bb_2_predecessor_in_state_1_in_data), .out_data(bb_2_predecessor_in_state_1_out_data));

	reg [0:0] bb_1_active_in_state_2_in_data;
	wire [0:0] bb_1_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_2(.in_data(bb_1_active_in_state_2_in_data), .out_data(bb_1_active_in_state_2_out_data));

	reg [31:0] bb_1_predecessor_in_state_2_in_data;
	wire [31:0] bb_1_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_2(.in_data(bb_1_predecessor_in_state_2_in_data), .out_data(bb_1_predecessor_in_state_2_out_data));

	reg [0:0] bb_2_active_in_state_2_in_data;
	wire [0:0] bb_2_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_2(.in_data(bb_2_active_in_state_2_in_data), .out_data(bb_2_active_in_state_2_out_data));

	reg [31:0] bb_2_predecessor_in_state_2_in_data;
	wire [31:0] bb_2_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_2(.in_data(bb_2_predecessor_in_state_2_in_data), .out_data(bb_2_predecessor_in_state_2_out_data));

	reg [0:0] bb_3_active_in_state_2_in_data;
	wire [0:0] bb_3_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_2(.in_data(bb_3_active_in_state_2_in_data), .out_data(bb_3_active_in_state_2_out_data));

	reg [31:0] bb_3_predecessor_in_state_2_in_data;
	wire [31:0] bb_3_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_2(.in_data(bb_3_predecessor_in_state_2_in_data), .out_data(bb_3_predecessor_in_state_2_out_data));

	reg [0:0] bb_4_active_in_state_2_in_data;
	wire [0:0] bb_4_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_2(.in_data(bb_4_active_in_state_2_in_data), .out_data(bb_4_active_in_state_2_out_data));

	reg [31:0] bb_4_predecessor_in_state_2_in_data;
	wire [31:0] bb_4_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_2(.in_data(bb_4_predecessor_in_state_2_in_data), .out_data(bb_4_predecessor_in_state_2_out_data));

	reg [0:0] andOp_42_in0;
	reg [0:0] andOp_42_in1;
	wire [0:0] andOp_42_out;
	andOp #(.WIDTH(1)) andOp_42(.in0(andOp_42_in0), .in1(andOp_42_in1), .out(andOp_42_out));

	reg [0:0] andOp_43_in0;
	reg [0:0] andOp_43_in1;
	wire [0:0] andOp_43_out;
	andOp #(.WIDTH(1)) andOp_43(.in0(andOp_43_in0), .in1(andOp_43_in1), .out(andOp_43_out));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] notOp_44_in0;
	wire [0:0] notOp_44_out;
	notOp #(.WIDTH(1)) notOp_44(.in(notOp_44_in0), .out(notOp_44_out));

	reg [0:0] andOp_45_in0;
	reg [0:0] andOp_45_in1;
	wire [0:0] andOp_45_out;
	andOp #(.WIDTH(1)) andOp_45(.in0(andOp_45_in0), .in1(andOp_45_in1), .out(andOp_45_out));

	reg [0:0] andOp_46_in0;
	reg [0:0] andOp_46_in1;
	wire [0:0] andOp_46_out;
	andOp #(.WIDTH(1)) andOp_46(.in0(andOp_46_in0), .in1(andOp_46_in1), .out(andOp_46_out));

	reg [0:0] br_2_happened_in_state_0_in_data;
	wire [0:0] br_2_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_2_happened_in_state_0(.in_data(br_2_happened_in_state_0_in_data), .out_data(br_2_happened_in_state_0_out_data));

	reg [0:0] notOp_47_in0;
	wire [0:0] notOp_47_out;
	notOp #(.WIDTH(1)) notOp_47(.in(notOp_47_in0), .out(notOp_47_out));

	reg [0:0] andOp_48_in0;
	reg [0:0] andOp_48_in1;
	wire [0:0] andOp_48_out;
	andOp #(.WIDTH(1)) andOp_48(.in0(andOp_48_in0), .in1(andOp_48_in1), .out(andOp_48_out));

	reg [0:0] andOp_49_in0;
	reg [0:0] andOp_49_in1;
	wire [0:0] andOp_49_out;
	andOp #(.WIDTH(1)) andOp_49(.in0(andOp_49_in0), .in1(andOp_49_in1), .out(andOp_49_out));

	reg [0:0] br_2_happened_in_state_1_in_data;
	wire [0:0] br_2_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_2_happened_in_state_1(.in_data(br_2_happened_in_state_1_in_data), .out_data(br_2_happened_in_state_1_out_data));

	reg [0:0] notOp_50_in0;
	wire [0:0] notOp_50_out;
	notOp #(.WIDTH(1)) notOp_50(.in(notOp_50_in0), .out(notOp_50_out));

	reg [0:0] andOp_51_in0;
	reg [0:0] andOp_51_in1;
	wire [0:0] andOp_51_out;
	andOp #(.WIDTH(1)) andOp_51(.in0(andOp_51_in0), .in1(andOp_51_in1), .out(andOp_51_out));

	reg [0:0] andOp_52_in0;
	reg [0:0] andOp_52_in1;
	wire [0:0] andOp_52_out;
	andOp #(.WIDTH(1)) andOp_52(.in0(andOp_52_in0), .in1(andOp_52_in1), .out(andOp_52_out));

	reg [0:0] br_2_happened_in_state_2_in_data;
	wire [0:0] br_2_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_2_happened_in_state_2(.in_data(br_2_happened_in_state_2_in_data), .out_data(br_2_happened_in_state_2_out_data));

	reg [0:0] notOp_53_in0;
	wire [0:0] notOp_53_out;
	notOp #(.WIDTH(1)) notOp_53(.in(notOp_53_in0), .out(notOp_53_out));

	reg [0:0] andOp_54_in0;
	reg [0:0] andOp_54_in1;
	wire [0:0] andOp_54_out;
	andOp #(.WIDTH(1)) andOp_54(.in0(andOp_54_in0), .in1(andOp_54_in1), .out(andOp_54_out));

	reg [0:0] andOp_55_in0;
	reg [0:0] andOp_55_in1;
	wire [0:0] andOp_55_out;
	andOp #(.WIDTH(1)) andOp_55(.in0(andOp_55_in0), .in1(andOp_55_in1), .out(andOp_55_out));

	reg [0:0] br_3_happened_in_state_2_in_data;
	wire [0:0] br_3_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_2(.in_data(br_3_happened_in_state_2_in_data), .out_data(br_3_happened_in_state_2_out_data));

	reg [0:0] notOp_56_in0;
	wire [0:0] notOp_56_out;
	notOp #(.WIDTH(1)) notOp_56(.in(notOp_56_in0), .out(notOp_56_out));

	reg [0:0] andOp_57_in0;
	reg [0:0] andOp_57_in1;
	wire [0:0] andOp_57_out;
	andOp #(.WIDTH(1)) andOp_57(.in0(andOp_57_in0), .in1(andOp_57_in1), .out(andOp_57_out));

	reg [0:0] andOp_58_in0;
	reg [0:0] andOp_58_in1;
	wire [0:0] andOp_58_out;
	andOp #(.WIDTH(1)) andOp_58(.in0(andOp_58_in0), .in1(andOp_58_in1), .out(andOp_58_out));

	reg [0:0] br_4_happened_in_state_2_in_data;
	wire [0:0] br_4_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_2(.in_data(br_4_happened_in_state_2_in_data), .out_data(br_4_happened_in_state_2_out_data));

	reg [0:0] notOp_59_in0;
	wire [0:0] notOp_59_out;
	notOp #(.WIDTH(1)) notOp_59(.in(notOp_59_in0), .out(notOp_59_out));

	reg [0:0] andOp_60_in0;
	reg [0:0] andOp_60_in1;
	wire [0:0] andOp_60_out;
	andOp #(.WIDTH(1)) andOp_60(.in0(andOp_60_in0), .in1(andOp_60_in1), .out(andOp_60_out));

	reg [0:0] notOp_61_in0;
	wire [0:0] notOp_61_out;
	notOp #(.WIDTH(1)) notOp_61(.in(notOp_61_in0), .out(notOp_61_out));

	reg [0:0] andOp_62_in0;
	reg [0:0] andOp_62_in1;
	wire [0:0] andOp_62_out;
	andOp #(.WIDTH(1)) andOp_62(.in0(andOp_62_in0), .in1(andOp_62_in1), .out(andOp_62_out));

	reg [31:0] eq_63_in0;
	reg [31:0] eq_63_in1;
	wire [0:0] eq_63_out;
	eq #(.WIDTH(32)) eq_63(.in0(eq_63_in0), .in1(eq_63_in1), .out(eq_63_out));

	reg [31:0] eq_64_in0;
	reg [31:0] eq_64_in1;
	wire [0:0] eq_64_out;
	eq #(.WIDTH(32)) eq_64(.in0(eq_64_in0), .in1(eq_64_in1), .out(eq_64_out));

	reg [0:0] orOp_65_in0;
	reg [0:0] orOp_65_in1;
	wire [0:0] orOp_65_out;
	orOp #(.WIDTH(1)) orOp_65(.in0(orOp_65_in0), .in1(orOp_65_in1), .out(orOp_65_out));

	reg [31:0] eq_66_in0;
	reg [31:0] eq_66_in1;
	wire [0:0] eq_66_out;
	eq #(.WIDTH(32)) eq_66(.in0(eq_66_in0), .in1(eq_66_in1), .out(eq_66_out));

	reg [31:0] eq_67_in0;
	reg [31:0] eq_67_in1;
	wire [0:0] eq_67_out;
	eq #(.WIDTH(32)) eq_67(.in0(eq_67_in0), .in1(eq_67_in1), .out(eq_67_out));

	reg [0:0] orOp_68_in0;
	reg [0:0] orOp_68_in1;
	wire [0:0] orOp_68_out;
	orOp #(.WIDTH(1)) orOp_68(.in0(orOp_68_in0), .in1(orOp_68_in1), .out(orOp_68_out));

	reg [31:0] eq_69_in0;
	reg [31:0] eq_69_in1;
	wire [0:0] eq_69_out;
	eq #(.WIDTH(32)) eq_69(.in0(eq_69_in0), .in1(eq_69_in1), .out(eq_69_out));

	reg [31:0] eq_70_in0;
	reg [31:0] eq_70_in1;
	wire [0:0] eq_70_out;
	eq #(.WIDTH(32)) eq_70(.in0(eq_70_in0), .in1(eq_70_in1), .out(eq_70_out));

	reg [0:0] orOp_71_in0;
	reg [0:0] orOp_71_in1;
	wire [0:0] orOp_71_out;
	orOp #(.WIDTH(1)) orOp_71(.in0(orOp_71_in0), .in1(orOp_71_in1), .out(orOp_71_out));

	reg [31:0] eq_72_in0;
	reg [31:0] eq_72_in1;
	wire [0:0] eq_72_out;
	eq #(.WIDTH(32)) eq_72(.in0(eq_72_in0), .in1(eq_72_in1), .out(eq_72_out));

	reg [0:0] orOp_73_in0;
	reg [0:0] orOp_73_in1;
	wire [0:0] orOp_73_out;
	orOp #(.WIDTH(1)) orOp_73(.in0(orOp_73_in0), .in1(orOp_73_in1), .out(orOp_73_out));

	reg [31:0] eq_74_in0;
	reg [31:0] eq_74_in1;
	wire [0:0] eq_74_out;
	eq #(.WIDTH(32)) eq_74(.in0(eq_74_in0), .in1(eq_74_in1), .out(eq_74_out));

	reg [31:0] eq_75_in0;
	reg [31:0] eq_75_in1;
	wire [0:0] eq_75_out;
	eq #(.WIDTH(32)) eq_75(.in0(eq_75_in0), .in1(eq_75_in1), .out(eq_75_out));

	reg [0:0] notOp_76_in0;
	wire [0:0] notOp_76_out;
	notOp #(.WIDTH(1)) notOp_76(.in(notOp_76_in0), .out(notOp_76_out));

	reg [0:0] andOp_77_in0;
	reg [0:0] andOp_77_in1;
	wire [0:0] andOp_77_out;
	andOp #(.WIDTH(1)) andOp_77(.in0(andOp_77_in0), .in1(andOp_77_in1), .out(andOp_77_out));

	reg [31:0] eq_78_in0;
	reg [31:0] eq_78_in1;
	wire [0:0] eq_78_out;
	eq #(.WIDTH(32)) eq_78(.in0(eq_78_in0), .in1(eq_78_in1), .out(eq_78_out));

	reg [31:0] eq_79_in0;
	reg [31:0] eq_79_in1;
	wire [0:0] eq_79_out;
	eq #(.WIDTH(32)) eq_79(.in0(eq_79_in0), .in1(eq_79_in1), .out(eq_79_out));

	reg [0:0] notOp_80_in0;
	wire [0:0] notOp_80_out;
	notOp #(.WIDTH(1)) notOp_80(.in(notOp_80_in0), .out(notOp_80_out));

	reg [0:0] andOp_81_in0;
	reg [0:0] andOp_81_in1;
	wire [0:0] andOp_81_out;
	andOp #(.WIDTH(1)) andOp_81(.in0(andOp_81_in0), .in1(andOp_81_in1), .out(andOp_81_out));

	reg [31:0] eq_82_in0;
	reg [31:0] eq_82_in1;
	wire [0:0] eq_82_out;
	eq #(.WIDTH(32)) eq_82(.in0(eq_82_in0), .in1(eq_82_in1), .out(eq_82_out));

	reg [31:0] eq_83_in0;
	reg [31:0] eq_83_in1;
	wire [0:0] eq_83_out;
	eq #(.WIDTH(32)) eq_83(.in0(eq_83_in0), .in1(eq_83_in1), .out(eq_83_out));

	reg [0:0] notOp_84_in0;
	wire [0:0] notOp_84_out;
	notOp #(.WIDTH(1)) notOp_84(.in(notOp_84_in0), .out(notOp_84_out));

	reg [0:0] andOp_85_in0;
	reg [0:0] andOp_85_in1;
	wire [0:0] andOp_85_out;
	andOp #(.WIDTH(1)) andOp_85(.in0(andOp_85_in0), .in1(andOp_85_in1), .out(andOp_85_out));

	reg [31:0] eq_86_in0;
	reg [31:0] eq_86_in1;
	wire [0:0] eq_86_out;
	eq #(.WIDTH(32)) eq_86(.in0(eq_86_in0), .in1(eq_86_in1), .out(eq_86_out));

	reg [0:0] notOp_87_in0;
	wire [0:0] notOp_87_out;
	notOp #(.WIDTH(1)) notOp_87(.in(notOp_87_in0), .out(notOp_87_out));

	reg [0:0] andOp_88_in0;
	reg [0:0] andOp_88_in1;
	wire [0:0] andOp_88_out;
	andOp #(.WIDTH(1)) andOp_88(.in0(andOp_88_in0), .in1(andOp_88_in1), .out(andOp_88_out));

	reg [0:0] andOp_89_in0;
	reg [0:0] andOp_89_in1;
	wire [0:0] andOp_89_out;
	andOp #(.WIDTH(1)) andOp_89(.in0(andOp_89_in0), .in1(andOp_89_in1), .out(andOp_89_out));

	reg [0:0] andOp_90_in0;
	reg [0:0] andOp_90_in1;
	wire [0:0] andOp_90_out;
	andOp #(.WIDTH(1)) andOp_90(.in0(andOp_90_in0), .in1(andOp_90_in1), .out(andOp_90_out));

	reg [0:0] andOp_91_in0;
	reg [0:0] andOp_91_in1;
	wire [0:0] andOp_91_out;
	andOp #(.WIDTH(1)) andOp_91(.in0(andOp_91_in0), .in1(andOp_91_in1), .out(andOp_91_out));

	reg [0:0] andOp_92_in0;
	reg [0:0] andOp_92_in1;
	wire [0:0] andOp_92_out;
	andOp #(.WIDTH(1)) andOp_92(.in0(andOp_92_in0), .in1(andOp_92_in1), .out(andOp_92_out));

	reg [0:0] andOp_93_in0;
	reg [0:0] andOp_93_in1;
	wire [0:0] andOp_93_out;
	andOp #(.WIDTH(1)) andOp_93(.in0(andOp_93_in0), .in1(andOp_93_in1), .out(andOp_93_out));

	reg [0:0] andOp_94_in0;
	reg [0:0] andOp_94_in1;
	wire [0:0] andOp_94_out;
	andOp #(.WIDTH(1)) andOp_94(.in0(andOp_94_in0), .in1(andOp_94_in1), .out(andOp_94_out));

	reg [0:0] andOp_95_in0;
	reg [0:0] andOp_95_in1;
	wire [0:0] andOp_95_out;
	andOp #(.WIDTH(1)) andOp_95(.in0(andOp_95_in0), .in1(andOp_95_in1), .out(andOp_95_out));

	reg [0:0] andOp_96_in0;
	reg [0:0] andOp_96_in1;
	wire [0:0] andOp_96_out;
	andOp #(.WIDTH(1)) andOp_96(.in0(andOp_96_in0), .in1(andOp_96_in1), .out(andOp_96_out));

	reg [0:0] andOp_97_in0;
	reg [0:0] andOp_97_in1;
	wire [0:0] andOp_97_out;
	andOp #(.WIDTH(1)) andOp_97(.in0(andOp_97_in0), .in1(andOp_97_in1), .out(andOp_97_out));

	reg [0:0] andOp_98_in0;
	reg [0:0] andOp_98_in1;
	wire [0:0] andOp_98_out;
	andOp #(.WIDTH(1)) andOp_98(.in0(andOp_98_in0), .in1(andOp_98_in1), .out(andOp_98_out));

	reg [31:0] concat_99_in0;
	reg [31:0] concat_99_in1;
	wire [63:0] concat_99_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_99(.in0(concat_99_in0), .in1(concat_99_in1), .out(concat_99_out));

	reg [31:0] concat_100_in0;
	reg [31:0] concat_100_in1;
	wire [63:0] concat_100_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_100(.in0(concat_100_in0), .in1(concat_100_in1), .out(concat_100_out));

	reg [0:0] andOp_101_in0;
	reg [0:0] andOp_101_in1;
	wire [0:0] andOp_101_out;
	andOp #(.WIDTH(1)) andOp_101(.in0(andOp_101_in0), .in1(andOp_101_in1), .out(andOp_101_out));

	reg [0:0] andOp_102_in0;
	reg [0:0] andOp_102_in1;
	wire [0:0] andOp_102_out;
	andOp #(.WIDTH(1)) andOp_102(.in0(andOp_102_in0), .in1(andOp_102_in1), .out(andOp_102_out));

	reg [0:0] andOp_103_in0;
	reg [0:0] andOp_103_in1;
	wire [0:0] andOp_103_out;
	andOp #(.WIDTH(1)) andOp_103(.in0(andOp_103_in0), .in1(andOp_103_in1), .out(andOp_103_out));

	reg [0:0] andOp_104_in0;
	reg [0:0] andOp_104_in1;
	wire [0:0] andOp_104_out;
	andOp #(.WIDTH(1)) andOp_104(.in0(andOp_104_in0), .in1(andOp_104_in1), .out(andOp_104_out));

	reg [0:0] andOp_105_in0;
	reg [0:0] andOp_105_in1;
	wire [0:0] andOp_105_out;
	andOp #(.WIDTH(1)) andOp_105(.in0(andOp_105_in0), .in1(andOp_105_in1), .out(andOp_105_out));

	reg [0:0] andOp_106_in0;
	reg [0:0] andOp_106_in1;
	wire [0:0] andOp_106_out;
	andOp #(.WIDTH(1)) andOp_106(.in0(andOp_106_in0), .in1(andOp_106_in1), .out(andOp_106_out));

	reg [0:0] andOp_107_in0;
	reg [0:0] andOp_107_in1;
	wire [0:0] andOp_107_out;
	andOp #(.WIDTH(1)) andOp_107(.in0(andOp_107_in0), .in1(andOp_107_in1), .out(andOp_107_out));

	reg [0:0] andOp_108_in0;
	reg [0:0] andOp_108_in1;
	wire [0:0] andOp_108_out;
	andOp #(.WIDTH(1)) andOp_108(.in0(andOp_108_in0), .in1(andOp_108_in1), .out(andOp_108_out));

	reg [0:0] andOp_109_in0;
	reg [0:0] andOp_109_in1;
	wire [0:0] andOp_109_out;
	andOp #(.WIDTH(1)) andOp_109(.in0(andOp_109_in0), .in1(andOp_109_in1), .out(andOp_109_out));

	reg [0:0] notOp_110_in0;
	wire [0:0] notOp_110_out;
	notOp #(.WIDTH(1)) notOp_110(.in(notOp_110_in0), .out(notOp_110_out));

	reg [0:0] andOp_111_in0;
	reg [0:0] andOp_111_in1;
	wire [0:0] andOp_111_out;
	andOp #(.WIDTH(1)) andOp_111(.in0(andOp_111_in0), .in1(andOp_111_in1), .out(andOp_111_out));

	reg [0:0] notOp_112_in0;
	wire [0:0] notOp_112_out;
	notOp #(.WIDTH(1)) notOp_112(.in(notOp_112_in0), .out(notOp_112_out));

	reg [0:0] andOp_113_in0;
	reg [0:0] andOp_113_in1;
	wire [0:0] andOp_113_out;
	andOp #(.WIDTH(1)) andOp_113(.in0(andOp_113_in0), .in1(andOp_113_in1), .out(andOp_113_out));

	reg [0:0] notOp_114_in0;
	wire [0:0] notOp_114_out;
	notOp #(.WIDTH(1)) notOp_114(.in(notOp_114_in0), .out(notOp_114_out));

	reg [0:0] andOp_115_in0;
	reg [0:0] andOp_115_in1;
	wire [0:0] andOp_115_out;
	andOp #(.WIDTH(1)) andOp_115(.in0(andOp_115_in0), .in1(andOp_115_in1), .out(andOp_115_out));

	reg [0:0] notOp_116_in0;
	wire [0:0] notOp_116_out;
	notOp #(.WIDTH(1)) notOp_116(.in(notOp_116_in0), .out(notOp_116_out));

	reg [0:0] andOp_117_in0;
	reg [0:0] andOp_117_in1;
	wire [0:0] andOp_117_out;
	andOp #(.WIDTH(1)) andOp_117(.in0(andOp_117_in0), .in1(andOp_117_in1), .out(andOp_117_out));

	reg [0:0] andOp_118_in0;
	reg [0:0] andOp_118_in1;
	wire [0:0] andOp_118_out;
	andOp #(.WIDTH(1)) andOp_118(.in0(andOp_118_in0), .in1(andOp_118_in1), .out(andOp_118_out));

	reg [31:0] eq_119_in0;
	reg [31:0] eq_119_in1;
	wire [0:0] eq_119_out;
	eq #(.WIDTH(32)) eq_119(.in0(eq_119_in0), .in1(eq_119_in1), .out(eq_119_out));

	reg [0:0] andOp_120_in0;
	reg [0:0] andOp_120_in1;
	wire [0:0] andOp_120_out;
	andOp #(.WIDTH(1)) andOp_120(.in0(andOp_120_in0), .in1(andOp_120_in1), .out(andOp_120_out));

	reg [31:0] eq_121_in0;
	reg [31:0] eq_121_in1;
	wire [0:0] eq_121_out;
	eq #(.WIDTH(32)) eq_121(.in0(eq_121_in0), .in1(eq_121_in1), .out(eq_121_out));

	reg [0:0] andOp_122_in0;
	reg [0:0] andOp_122_in1;
	wire [0:0] andOp_122_out;
	andOp #(.WIDTH(1)) andOp_122(.in0(andOp_122_in0), .in1(andOp_122_in1), .out(andOp_122_out));

	reg [31:0] eq_123_in0;
	reg [31:0] eq_123_in1;
	wire [0:0] eq_123_out;
	eq #(.WIDTH(32)) eq_123(.in0(eq_123_in0), .in1(eq_123_in1), .out(eq_123_out));

	reg [0:0] andOp_124_in0;
	reg [0:0] andOp_124_in1;
	wire [0:0] andOp_124_out;
	andOp #(.WIDTH(1)) andOp_124(.in0(andOp_124_in0), .in1(andOp_124_in1), .out(andOp_124_out));

	reg [0:0] andOp_125_in0;
	reg [0:0] andOp_125_in1;
	wire [0:0] andOp_125_out;
	andOp #(.WIDTH(1)) andOp_125(.in0(andOp_125_in0), .in1(andOp_125_in1), .out(andOp_125_out));

	reg [31:0] eq_126_in0;
	reg [31:0] eq_126_in1;
	wire [0:0] eq_126_out;
	eq #(.WIDTH(32)) eq_126(.in0(eq_126_in0), .in1(eq_126_in1), .out(eq_126_out));

	reg [0:0] andOp_127_in0;
	reg [0:0] andOp_127_in1;
	wire [0:0] andOp_127_out;
	andOp #(.WIDTH(1)) andOp_127(.in0(andOp_127_in0), .in1(andOp_127_in1), .out(andOp_127_out));

	reg [0:0] notOp_128_in0;
	wire [0:0] notOp_128_out;
	notOp #(.WIDTH(1)) notOp_128(.in(notOp_128_in0), .out(notOp_128_out));

	reg [0:0] andOp_129_in0;
	reg [0:0] andOp_129_in1;
	wire [0:0] andOp_129_out;
	andOp #(.WIDTH(1)) andOp_129(.in0(andOp_129_in0), .in1(andOp_129_in1), .out(andOp_129_out));

	reg [0:0] notOp_130_in0;
	wire [0:0] notOp_130_out;
	notOp #(.WIDTH(1)) notOp_130(.in(notOp_130_in0), .out(notOp_130_out));

	reg [0:0] andOp_131_in0;
	reg [0:0] andOp_131_in1;
	wire [0:0] andOp_131_out;
	andOp #(.WIDTH(1)) andOp_131(.in0(andOp_131_in0), .in1(andOp_131_in1), .out(andOp_131_out));

	reg [0:0] notOp_132_in0;
	wire [0:0] notOp_132_out;
	notOp #(.WIDTH(1)) notOp_132(.in(notOp_132_in0), .out(notOp_132_out));

	reg [0:0] andOp_133_in0;
	reg [0:0] andOp_133_in1;
	wire [0:0] andOp_133_out;
	andOp #(.WIDTH(1)) andOp_133(.in0(andOp_133_in0), .in1(andOp_133_in1), .out(andOp_133_out));

	reg [0:0] andOp_134_in0;
	reg [0:0] andOp_134_in1;
	wire [0:0] andOp_134_out;
	andOp #(.WIDTH(1)) andOp_134(.in0(andOp_134_in0), .in1(andOp_134_in1), .out(andOp_134_out));

	reg [31:0] eq_135_in0;
	reg [31:0] eq_135_in1;
	wire [0:0] eq_135_out;
	eq #(.WIDTH(32)) eq_135(.in0(eq_135_in0), .in1(eq_135_in1), .out(eq_135_out));

	reg [0:0] andOp_136_in0;
	reg [0:0] andOp_136_in1;
	wire [0:0] andOp_136_out;
	andOp #(.WIDTH(1)) andOp_136(.in0(andOp_136_in0), .in1(andOp_136_in1), .out(andOp_136_out));

	reg [0:0] notOp_137_in0;
	wire [0:0] notOp_137_out;
	notOp #(.WIDTH(1)) notOp_137(.in(notOp_137_in0), .out(notOp_137_out));

	reg [0:0] andOp_138_in0;
	reg [0:0] andOp_138_in1;
	wire [0:0] andOp_138_out;
	andOp #(.WIDTH(1)) andOp_138(.in0(andOp_138_in0), .in1(andOp_138_in1), .out(andOp_138_out));

	reg [0:0] notOp_139_in0;
	wire [0:0] notOp_139_out;
	notOp #(.WIDTH(1)) notOp_139(.in(notOp_139_in0), .out(notOp_139_out));

	reg [0:0] andOp_140_in0;
	reg [0:0] andOp_140_in1;
	wire [0:0] andOp_140_out;
	andOp #(.WIDTH(1)) andOp_140(.in0(andOp_140_in0), .in1(andOp_140_in1), .out(andOp_140_out));

	reg [0:0] notOp_141_in0;
	wire [0:0] notOp_141_out;
	notOp #(.WIDTH(1)) notOp_141(.in(notOp_141_in0), .out(notOp_141_out));

	reg [0:0] andOp_142_in0;
	reg [0:0] andOp_142_in1;
	wire [0:0] andOp_142_out;
	andOp #(.WIDTH(1)) andOp_142(.in0(andOp_142_in0), .in1(andOp_142_in1), .out(andOp_142_out));

	reg [0:0] andOp_143_in0;
	reg [0:0] andOp_143_in1;
	wire [0:0] andOp_143_out;
	andOp #(.WIDTH(1)) andOp_143(.in0(andOp_143_in0), .in1(andOp_143_in1), .out(andOp_143_out));

	reg [31:0] eq_144_in0;
	reg [31:0] eq_144_in1;
	wire [0:0] eq_144_out;
	eq #(.WIDTH(32)) eq_144(.in0(eq_144_in0), .in1(eq_144_in1), .out(eq_144_out));

	reg [0:0] andOp_145_in0;
	reg [0:0] andOp_145_in1;
	wire [0:0] andOp_145_out;
	andOp #(.WIDTH(1)) andOp_145(.in0(andOp_145_in0), .in1(andOp_145_in1), .out(andOp_145_out));

	reg [0:0] notOp_146_in0;
	wire [0:0] notOp_146_out;
	notOp #(.WIDTH(1)) notOp_146(.in(notOp_146_in0), .out(notOp_146_out));

	reg [0:0] andOp_147_in0;
	reg [0:0] andOp_147_in1;
	wire [0:0] andOp_147_out;
	andOp #(.WIDTH(1)) andOp_147(.in0(andOp_147_in0), .in1(andOp_147_in1), .out(andOp_147_out));

	reg [0:0] notOp_148_in0;
	wire [0:0] notOp_148_out;
	notOp #(.WIDTH(1)) notOp_148(.in(notOp_148_in0), .out(notOp_148_out));

	reg [0:0] andOp_149_in0;
	reg [0:0] andOp_149_in1;
	wire [0:0] andOp_149_out;
	andOp #(.WIDTH(1)) andOp_149(.in0(andOp_149_in0), .in1(andOp_149_in1), .out(andOp_149_out));

	reg [0:0] notOp_150_in0;
	wire [0:0] notOp_150_out;
	notOp #(.WIDTH(1)) notOp_150(.in(notOp_150_in0), .out(notOp_150_out));

	reg [0:0] andOp_151_in0;
	reg [0:0] andOp_151_in1;
	wire [0:0] andOp_151_out;
	andOp #(.WIDTH(1)) andOp_151(.in0(andOp_151_in0), .in1(andOp_151_in1), .out(andOp_151_out));

	reg [0:0] andOp_152_in0;
	reg [0:0] andOp_152_in1;
	wire [0:0] andOp_152_out;
	andOp #(.WIDTH(1)) andOp_152(.in0(andOp_152_in0), .in1(andOp_152_in1), .out(andOp_152_out));

	reg [31:0] eq_153_in0;
	reg [31:0] eq_153_in1;
	wire [0:0] eq_153_out;
	eq #(.WIDTH(32)) eq_153(.in0(eq_153_in0), .in1(eq_153_in1), .out(eq_153_out));

	reg [0:0] andOp_154_in0;
	reg [0:0] andOp_154_in1;
	wire [0:0] andOp_154_out;
	andOp #(.WIDTH(1)) andOp_154(.in0(andOp_154_in0), .in1(andOp_154_in1), .out(andOp_154_out));

	reg [0:0] notOp_155_in0;
	wire [0:0] notOp_155_out;
	notOp #(.WIDTH(1)) notOp_155(.in(notOp_155_in0), .out(notOp_155_out));

	reg [0:0] andOp_156_in0;
	reg [0:0] andOp_156_in1;
	wire [0:0] andOp_156_out;
	andOp #(.WIDTH(1)) andOp_156(.in0(andOp_156_in0), .in1(andOp_156_in1), .out(andOp_156_out));

	reg [0:0] notOp_157_in0;
	wire [0:0] notOp_157_out;
	notOp #(.WIDTH(1)) notOp_157(.in(notOp_157_in0), .out(notOp_157_out));

	reg [0:0] andOp_158_in0;
	reg [0:0] andOp_158_in1;
	wire [0:0] andOp_158_out;
	andOp #(.WIDTH(1)) andOp_158(.in0(andOp_158_in0), .in1(andOp_158_in1), .out(andOp_158_out));

	reg [0:0] notOp_159_in0;
	wire [0:0] notOp_159_out;
	notOp #(.WIDTH(1)) notOp_159(.in(notOp_159_in0), .out(notOp_159_out));

	reg [0:0] andOp_160_in0;
	reg [0:0] andOp_160_in1;
	wire [0:0] andOp_160_out;
	andOp #(.WIDTH(1)) andOp_160(.in0(andOp_160_in0), .in1(andOp_160_in1), .out(andOp_160_out));

	reg [0:0] andOp_161_in0;
	reg [0:0] andOp_161_in1;
	wire [0:0] andOp_161_out;
	andOp #(.WIDTH(1)) andOp_161(.in0(andOp_161_in0), .in1(andOp_161_in1), .out(andOp_161_out));

	reg [31:0] eq_162_in0;
	reg [31:0] eq_162_in1;
	wire [0:0] eq_162_out;
	eq #(.WIDTH(32)) eq_162(.in0(eq_162_in0), .in1(eq_162_in1), .out(eq_162_out));

	reg [0:0] andOp_163_in0;
	reg [0:0] andOp_163_in1;
	wire [0:0] andOp_163_out;
	andOp #(.WIDTH(1)) andOp_163(.in0(andOp_163_in0), .in1(andOp_163_in1), .out(andOp_163_out));

	reg [0:0] notOp_164_in0;
	wire [0:0] notOp_164_out;
	notOp #(.WIDTH(1)) notOp_164(.in(notOp_164_in0), .out(notOp_164_out));

	reg [0:0] andOp_165_in0;
	reg [0:0] andOp_165_in1;
	wire [0:0] andOp_165_out;
	andOp #(.WIDTH(1)) andOp_165(.in0(andOp_165_in0), .in1(andOp_165_in1), .out(andOp_165_out));

	reg [0:0] notOp_166_in0;
	wire [0:0] notOp_166_out;
	notOp #(.WIDTH(1)) notOp_166(.in(notOp_166_in0), .out(notOp_166_out));

	reg [0:0] andOp_167_in0;
	reg [0:0] andOp_167_in1;
	wire [0:0] andOp_167_out;
	andOp #(.WIDTH(1)) andOp_167(.in0(andOp_167_in0), .in1(andOp_167_in1), .out(andOp_167_out));

	reg [0:0] notOp_168_in0;
	wire [0:0] notOp_168_out;
	notOp #(.WIDTH(1)) notOp_168(.in(notOp_168_in0), .out(notOp_168_out));

	reg [0:0] andOp_169_in0;
	reg [0:0] andOp_169_in1;
	wire [0:0] andOp_169_out;
	andOp #(.WIDTH(1)) andOp_169(.in0(andOp_169_in0), .in1(andOp_169_in1), .out(andOp_169_out));

	reg [0:0] andOp_170_in0;
	reg [0:0] andOp_170_in1;
	wire [0:0] andOp_170_out;
	andOp #(.WIDTH(1)) andOp_170(.in0(andOp_170_in0), .in1(andOp_170_in1), .out(andOp_170_out));

	reg [31:0] eq_171_in0;
	reg [31:0] eq_171_in1;
	wire [0:0] eq_171_out;
	eq #(.WIDTH(32)) eq_171(.in0(eq_171_in0), .in1(eq_171_in1), .out(eq_171_out));

	reg [0:0] andOp_172_in0;
	reg [0:0] andOp_172_in1;
	wire [0:0] andOp_172_out;
	andOp #(.WIDTH(1)) andOp_172(.in0(andOp_172_in0), .in1(andOp_172_in1), .out(andOp_172_out));

	reg [0:0] notOp_173_in0;
	wire [0:0] notOp_173_out;
	notOp #(.WIDTH(1)) notOp_173(.in(notOp_173_in0), .out(notOp_173_out));

	reg [0:0] andOp_174_in0;
	reg [0:0] andOp_174_in1;
	wire [0:0] andOp_174_out;
	andOp #(.WIDTH(1)) andOp_174(.in0(andOp_174_in0), .in1(andOp_174_in1), .out(andOp_174_out));

	reg [0:0] notOp_175_in0;
	wire [0:0] notOp_175_out;
	notOp #(.WIDTH(1)) notOp_175(.in(notOp_175_in0), .out(notOp_175_out));

	reg [0:0] andOp_176_in0;
	reg [0:0] andOp_176_in1;
	wire [0:0] andOp_176_out;
	andOp #(.WIDTH(1)) andOp_176(.in0(andOp_176_in0), .in1(andOp_176_in1), .out(andOp_176_out));

	reg [0:0] notOp_177_in0;
	wire [0:0] notOp_177_out;
	notOp #(.WIDTH(1)) notOp_177(.in(notOp_177_in0), .out(notOp_177_out));

	reg [0:0] andOp_178_in0;
	reg [0:0] andOp_178_in1;
	wire [0:0] andOp_178_out;
	andOp #(.WIDTH(1)) andOp_178(.in0(andOp_178_in0), .in1(andOp_178_in1), .out(andOp_178_out));

	reg [0:0] andOp_179_in0;
	reg [0:0] andOp_179_in1;
	wire [0:0] andOp_179_out;
	andOp #(.WIDTH(1)) andOp_179(.in0(andOp_179_in0), .in1(andOp_179_in1), .out(andOp_179_out));

	reg [31:0] eq_180_in0;
	reg [31:0] eq_180_in1;
	wire [0:0] eq_180_out;
	eq #(.WIDTH(32)) eq_180(.in0(eq_180_in0), .in1(eq_180_in1), .out(eq_180_out));

	reg [0:0] andOp_181_in0;
	reg [0:0] andOp_181_in1;
	wire [0:0] andOp_181_out;
	andOp #(.WIDTH(1)) andOp_181(.in0(andOp_181_in0), .in1(andOp_181_in1), .out(andOp_181_out));

	reg [0:0] notOp_182_in0;
	wire [0:0] notOp_182_out;
	notOp #(.WIDTH(1)) notOp_182(.in(notOp_182_in0), .out(notOp_182_out));

	reg [0:0] andOp_183_in0;
	reg [0:0] andOp_183_in1;
	wire [0:0] andOp_183_out;
	andOp #(.WIDTH(1)) andOp_183(.in0(andOp_183_in0), .in1(andOp_183_in1), .out(andOp_183_out));

	reg [0:0] notOp_184_in0;
	wire [0:0] notOp_184_out;
	notOp #(.WIDTH(1)) notOp_184(.in(notOp_184_in0), .out(notOp_184_out));

	reg [0:0] andOp_185_in0;
	reg [0:0] andOp_185_in1;
	wire [0:0] andOp_185_out;
	andOp #(.WIDTH(1)) andOp_185(.in0(andOp_185_in0), .in1(andOp_185_in1), .out(andOp_185_out));

	reg [0:0] notOp_186_in0;
	wire [0:0] notOp_186_out;
	notOp #(.WIDTH(1)) notOp_186(.in(notOp_186_in0), .out(notOp_186_out));

	reg [0:0] andOp_187_in0;
	reg [0:0] andOp_187_in1;
	wire [0:0] andOp_187_out;
	andOp #(.WIDTH(1)) andOp_187(.in0(andOp_187_in0), .in1(andOp_187_in1), .out(andOp_187_out));

	reg [31:0] eq_188_in0;
	reg [31:0] eq_188_in1;
	wire [0:0] eq_188_out;
	eq #(.WIDTH(32)) eq_188(.in0(eq_188_in0), .in1(eq_188_in1), .out(eq_188_out));

	reg [0:0] andOp_189_in0;
	reg [0:0] andOp_189_in1;
	wire [0:0] andOp_189_out;
	andOp #(.WIDTH(1)) andOp_189(.in0(andOp_189_in0), .in1(andOp_189_in1), .out(andOp_189_out));

	reg [31:0] eq_190_in0;
	reg [31:0] eq_190_in1;
	wire [0:0] eq_190_out;
	eq #(.WIDTH(32)) eq_190(.in0(eq_190_in0), .in1(eq_190_in1), .out(eq_190_out));

	reg [0:0] andOp_191_in0;
	reg [0:0] andOp_191_in1;
	wire [0:0] andOp_191_out;
	andOp #(.WIDTH(1)) andOp_191(.in0(andOp_191_in0), .in1(andOp_191_in1), .out(andOp_191_out));

	reg [31:0] eq_192_in0;
	reg [31:0] eq_192_in1;
	wire [0:0] eq_192_out;
	eq #(.WIDTH(32)) eq_192(.in0(eq_192_in0), .in1(eq_192_in1), .out(eq_192_out));

	reg [0:0] andOp_193_in0;
	reg [0:0] andOp_193_in1;
	wire [0:0] andOp_193_out;
	andOp #(.WIDTH(1)) andOp_193(.in0(andOp_193_in0), .in1(andOp_193_in1), .out(andOp_193_out));

	reg [0:0] andOp_194_in0;
	reg [0:0] andOp_194_in1;
	wire [0:0] andOp_194_out;
	andOp #(.WIDTH(1)) andOp_194(.in0(andOp_194_in0), .in1(andOp_194_in1), .out(andOp_194_out));

	reg [31:0] eq_195_in0;
	reg [31:0] eq_195_in1;
	wire [0:0] eq_195_out;
	eq #(.WIDTH(32)) eq_195(.in0(eq_195_in0), .in1(eq_195_in1), .out(eq_195_out));

	reg [0:0] andOp_196_in0;
	reg [0:0] andOp_196_in1;
	wire [0:0] andOp_196_out;
	andOp #(.WIDTH(1)) andOp_196(.in0(andOp_196_in0), .in1(andOp_196_in1), .out(andOp_196_out));

	reg [0:0] notOp_197_in0;
	wire [0:0] notOp_197_out;
	notOp #(.WIDTH(1)) notOp_197(.in(notOp_197_in0), .out(notOp_197_out));

	reg [0:0] andOp_198_in0;
	reg [0:0] andOp_198_in1;
	wire [0:0] andOp_198_out;
	andOp #(.WIDTH(1)) andOp_198(.in0(andOp_198_in0), .in1(andOp_198_in1), .out(andOp_198_out));

	reg [0:0] notOp_199_in0;
	wire [0:0] notOp_199_out;
	notOp #(.WIDTH(1)) notOp_199(.in(notOp_199_in0), .out(notOp_199_out));

	reg [0:0] andOp_200_in0;
	reg [0:0] andOp_200_in1;
	wire [0:0] andOp_200_out;
	andOp #(.WIDTH(1)) andOp_200(.in0(andOp_200_in0), .in1(andOp_200_in1), .out(andOp_200_out));

	reg [0:0] notOp_201_in0;
	wire [0:0] notOp_201_out;
	notOp #(.WIDTH(1)) notOp_201(.in(notOp_201_in0), .out(notOp_201_out));

	reg [0:0] andOp_202_in0;
	reg [0:0] andOp_202_in1;
	wire [0:0] andOp_202_out;
	andOp #(.WIDTH(1)) andOp_202(.in0(andOp_202_in0), .in1(andOp_202_in1), .out(andOp_202_out));

	reg [0:0] andOp_203_in0;
	reg [0:0] andOp_203_in1;
	wire [0:0] andOp_203_out;
	andOp #(.WIDTH(1)) andOp_203(.in0(andOp_203_in0), .in1(andOp_203_in1), .out(andOp_203_out));

	reg [31:0] eq_204_in0;
	reg [31:0] eq_204_in1;
	wire [0:0] eq_204_out;
	eq #(.WIDTH(32)) eq_204(.in0(eq_204_in0), .in1(eq_204_in1), .out(eq_204_out));

	reg [0:0] andOp_205_in0;
	reg [0:0] andOp_205_in1;
	wire [0:0] andOp_205_out;
	andOp #(.WIDTH(1)) andOp_205(.in0(andOp_205_in0), .in1(andOp_205_in1), .out(andOp_205_out));

	reg [0:0] notOp_206_in0;
	wire [0:0] notOp_206_out;
	notOp #(.WIDTH(1)) notOp_206(.in(notOp_206_in0), .out(notOp_206_out));

	reg [0:0] andOp_207_in0;
	reg [0:0] andOp_207_in1;
	wire [0:0] andOp_207_out;
	andOp #(.WIDTH(1)) andOp_207(.in0(andOp_207_in0), .in1(andOp_207_in1), .out(andOp_207_out));

	reg [0:0] notOp_208_in0;
	wire [0:0] notOp_208_out;
	notOp #(.WIDTH(1)) notOp_208(.in(notOp_208_in0), .out(notOp_208_out));

	reg [0:0] andOp_209_in0;
	reg [0:0] andOp_209_in1;
	wire [0:0] andOp_209_out;
	andOp #(.WIDTH(1)) andOp_209(.in0(andOp_209_in0), .in1(andOp_209_in1), .out(andOp_209_out));

	reg [0:0] notOp_210_in0;
	wire [0:0] notOp_210_out;
	notOp #(.WIDTH(1)) notOp_210(.in(notOp_210_in0), .out(notOp_210_out));

	reg [0:0] andOp_211_in0;
	reg [0:0] andOp_211_in1;
	wire [0:0] andOp_211_out;
	andOp #(.WIDTH(1)) andOp_211(.in0(andOp_211_in0), .in1(andOp_211_in1), .out(andOp_211_out));

	reg [0:0] andOp_212_in0;
	reg [0:0] andOp_212_in1;
	wire [0:0] andOp_212_out;
	andOp #(.WIDTH(1)) andOp_212(.in0(andOp_212_in0), .in1(andOp_212_in1), .out(andOp_212_out));

	reg [31:0] eq_213_in0;
	reg [31:0] eq_213_in1;
	wire [0:0] eq_213_out;
	eq #(.WIDTH(32)) eq_213(.in0(eq_213_in0), .in1(eq_213_in1), .out(eq_213_out));

	reg [0:0] andOp_214_in0;
	reg [0:0] andOp_214_in1;
	wire [0:0] andOp_214_out;
	andOp #(.WIDTH(1)) andOp_214(.in0(andOp_214_in0), .in1(andOp_214_in1), .out(andOp_214_out));

	reg [0:0] notOp_215_in0;
	wire [0:0] notOp_215_out;
	notOp #(.WIDTH(1)) notOp_215(.in(notOp_215_in0), .out(notOp_215_out));

	reg [0:0] andOp_216_in0;
	reg [0:0] andOp_216_in1;
	wire [0:0] andOp_216_out;
	andOp #(.WIDTH(1)) andOp_216(.in0(andOp_216_in0), .in1(andOp_216_in1), .out(andOp_216_out));

	reg [0:0] notOp_217_in0;
	wire [0:0] notOp_217_out;
	notOp #(.WIDTH(1)) notOp_217(.in(notOp_217_in0), .out(notOp_217_out));

	reg [0:0] andOp_218_in0;
	reg [0:0] andOp_218_in1;
	wire [0:0] andOp_218_out;
	andOp #(.WIDTH(1)) andOp_218(.in0(andOp_218_in0), .in1(andOp_218_in1), .out(andOp_218_out));

	reg [0:0] notOp_219_in0;
	wire [0:0] notOp_219_out;
	notOp #(.WIDTH(1)) notOp_219(.in(notOp_219_in0), .out(notOp_219_out));

	reg [0:0] andOp_220_in0;
	reg [0:0] andOp_220_in1;
	wire [0:0] andOp_220_out;
	andOp #(.WIDTH(1)) andOp_220(.in0(andOp_220_in0), .in1(andOp_220_in1), .out(andOp_220_out));

	reg [0:0] andOp_221_in0;
	reg [0:0] andOp_221_in1;
	wire [0:0] andOp_221_out;
	andOp #(.WIDTH(1)) andOp_221(.in0(andOp_221_in0), .in1(andOp_221_in1), .out(andOp_221_out));

	reg [31:0] eq_222_in0;
	reg [31:0] eq_222_in1;
	wire [0:0] eq_222_out;
	eq #(.WIDTH(32)) eq_222(.in0(eq_222_in0), .in1(eq_222_in1), .out(eq_222_out));

	reg [0:0] andOp_223_in0;
	reg [0:0] andOp_223_in1;
	wire [0:0] andOp_223_out;
	andOp #(.WIDTH(1)) andOp_223(.in0(andOp_223_in0), .in1(andOp_223_in1), .out(andOp_223_out));

	reg [0:0] notOp_224_in0;
	wire [0:0] notOp_224_out;
	notOp #(.WIDTH(1)) notOp_224(.in(notOp_224_in0), .out(notOp_224_out));

	reg [0:0] andOp_225_in0;
	reg [0:0] andOp_225_in1;
	wire [0:0] andOp_225_out;
	andOp #(.WIDTH(1)) andOp_225(.in0(andOp_225_in0), .in1(andOp_225_in1), .out(andOp_225_out));

	reg [0:0] notOp_226_in0;
	wire [0:0] notOp_226_out;
	notOp #(.WIDTH(1)) notOp_226(.in(notOp_226_in0), .out(notOp_226_out));

	reg [0:0] andOp_227_in0;
	reg [0:0] andOp_227_in1;
	wire [0:0] andOp_227_out;
	andOp #(.WIDTH(1)) andOp_227(.in0(andOp_227_in0), .in1(andOp_227_in1), .out(andOp_227_out));

	reg [0:0] notOp_228_in0;
	wire [0:0] notOp_228_out;
	notOp #(.WIDTH(1)) notOp_228(.in(notOp_228_in0), .out(notOp_228_out));

	reg [0:0] andOp_229_in0;
	reg [0:0] andOp_229_in1;
	wire [0:0] andOp_229_out;
	andOp #(.WIDTH(1)) andOp_229(.in0(andOp_229_in0), .in1(andOp_229_in1), .out(andOp_229_out));

	reg [0:0] andOp_230_in0;
	reg [0:0] andOp_230_in1;
	wire [0:0] andOp_230_out;
	andOp #(.WIDTH(1)) andOp_230(.in0(andOp_230_in0), .in1(andOp_230_in1), .out(andOp_230_out));

	reg [31:0] eq_231_in0;
	reg [31:0] eq_231_in1;
	wire [0:0] eq_231_out;
	eq #(.WIDTH(32)) eq_231(.in0(eq_231_in0), .in1(eq_231_in1), .out(eq_231_out));

	reg [0:0] andOp_232_in0;
	reg [0:0] andOp_232_in1;
	wire [0:0] andOp_232_out;
	andOp #(.WIDTH(1)) andOp_232(.in0(andOp_232_in0), .in1(andOp_232_in1), .out(andOp_232_out));

	reg [0:0] notOp_233_in0;
	wire [0:0] notOp_233_out;
	notOp #(.WIDTH(1)) notOp_233(.in(notOp_233_in0), .out(notOp_233_out));

	reg [0:0] andOp_234_in0;
	reg [0:0] andOp_234_in1;
	wire [0:0] andOp_234_out;
	andOp #(.WIDTH(1)) andOp_234(.in0(andOp_234_in0), .in1(andOp_234_in1), .out(andOp_234_out));

	reg [0:0] notOp_235_in0;
	wire [0:0] notOp_235_out;
	notOp #(.WIDTH(1)) notOp_235(.in(notOp_235_in0), .out(notOp_235_out));

	reg [0:0] andOp_236_in0;
	reg [0:0] andOp_236_in1;
	wire [0:0] andOp_236_out;
	andOp #(.WIDTH(1)) andOp_236(.in0(andOp_236_in0), .in1(andOp_236_in1), .out(andOp_236_out));

	reg [0:0] notOp_237_in0;
	wire [0:0] notOp_237_out;
	notOp #(.WIDTH(1)) notOp_237(.in(notOp_237_in0), .out(notOp_237_out));

	reg [0:0] andOp_238_in0;
	reg [0:0] andOp_238_in1;
	wire [0:0] andOp_238_out;
	andOp #(.WIDTH(1)) andOp_238(.in0(andOp_238_in0), .in1(andOp_238_in1), .out(andOp_238_out));

	reg [0:0] andOp_239_in0;
	reg [0:0] andOp_239_in1;
	wire [0:0] andOp_239_out;
	andOp #(.WIDTH(1)) andOp_239(.in0(andOp_239_in0), .in1(andOp_239_in1), .out(andOp_239_out));

	reg [31:0] eq_240_in0;
	reg [31:0] eq_240_in1;
	wire [0:0] eq_240_out;
	eq #(.WIDTH(32)) eq_240(.in0(eq_240_in0), .in1(eq_240_in1), .out(eq_240_out));

	reg [0:0] andOp_241_in0;
	reg [0:0] andOp_241_in1;
	wire [0:0] andOp_241_out;
	andOp #(.WIDTH(1)) andOp_241(.in0(andOp_241_in0), .in1(andOp_241_in1), .out(andOp_241_out));

	reg [0:0] notOp_242_in0;
	wire [0:0] notOp_242_out;
	notOp #(.WIDTH(1)) notOp_242(.in(notOp_242_in0), .out(notOp_242_out));

	reg [0:0] andOp_243_in0;
	reg [0:0] andOp_243_in1;
	wire [0:0] andOp_243_out;
	andOp #(.WIDTH(1)) andOp_243(.in0(andOp_243_in0), .in1(andOp_243_in1), .out(andOp_243_out));

	reg [0:0] notOp_244_in0;
	wire [0:0] notOp_244_out;
	notOp #(.WIDTH(1)) notOp_244(.in(notOp_244_in0), .out(notOp_244_out));

	reg [0:0] andOp_245_in0;
	reg [0:0] andOp_245_in1;
	wire [0:0] andOp_245_out;
	andOp #(.WIDTH(1)) andOp_245(.in0(andOp_245_in0), .in1(andOp_245_in1), .out(andOp_245_out));

	reg [0:0] notOp_246_in0;
	wire [0:0] notOp_246_out;
	notOp #(.WIDTH(1)) notOp_246(.in(notOp_246_in0), .out(notOp_246_out));

	reg [0:0] andOp_247_in0;
	reg [0:0] andOp_247_in1;
	wire [0:0] andOp_247_out;
	andOp #(.WIDTH(1)) andOp_247(.in0(andOp_247_in0), .in1(andOp_247_in1), .out(andOp_247_out));

	reg [0:0] andOp_248_in0;
	reg [0:0] andOp_248_in1;
	wire [0:0] andOp_248_out;
	andOp #(.WIDTH(1)) andOp_248(.in0(andOp_248_in0), .in1(andOp_248_in1), .out(andOp_248_out));

	reg [31:0] eq_249_in0;
	reg [31:0] eq_249_in1;
	wire [0:0] eq_249_out;
	eq #(.WIDTH(32)) eq_249(.in0(eq_249_in0), .in1(eq_249_in1), .out(eq_249_out));

	reg [0:0] andOp_250_in0;
	reg [0:0] andOp_250_in1;
	wire [0:0] andOp_250_out;
	andOp #(.WIDTH(1)) andOp_250(.in0(andOp_250_in0), .in1(andOp_250_in1), .out(andOp_250_out));

	reg [0:0] notOp_251_in0;
	wire [0:0] notOp_251_out;
	notOp #(.WIDTH(1)) notOp_251(.in(notOp_251_in0), .out(notOp_251_out));

	reg [0:0] andOp_252_in0;
	reg [0:0] andOp_252_in1;
	wire [0:0] andOp_252_out;
	andOp #(.WIDTH(1)) andOp_252(.in0(andOp_252_in0), .in1(andOp_252_in1), .out(andOp_252_out));

	reg [0:0] notOp_253_in0;
	wire [0:0] notOp_253_out;
	notOp #(.WIDTH(1)) notOp_253(.in(notOp_253_in0), .out(notOp_253_out));

	reg [0:0] andOp_254_in0;
	reg [0:0] andOp_254_in1;
	wire [0:0] andOp_254_out;
	andOp #(.WIDTH(1)) andOp_254(.in0(andOp_254_in0), .in1(andOp_254_in1), .out(andOp_254_out));

	reg [0:0] notOp_255_in0;
	wire [0:0] notOp_255_out;
	notOp #(.WIDTH(1)) notOp_255(.in(notOp_255_in0), .out(notOp_255_out));

	reg [0:0] andOp_256_in0;
	reg [0:0] andOp_256_in1;
	wire [0:0] andOp_256_out;
	andOp #(.WIDTH(1)) andOp_256(.in0(andOp_256_in0), .in1(andOp_256_in1), .out(andOp_256_out));

	reg [31:0] eq_257_in0;
	reg [31:0] eq_257_in1;
	wire [0:0] eq_257_out;
	eq #(.WIDTH(32)) eq_257(.in0(eq_257_in0), .in1(eq_257_in1), .out(eq_257_out));

	reg [0:0] andOp_258_in0;
	reg [0:0] andOp_258_in1;
	wire [0:0] andOp_258_out;
	andOp #(.WIDTH(1)) andOp_258(.in0(andOp_258_in0), .in1(andOp_258_in1), .out(andOp_258_out));

	reg [31:0] eq_259_in0;
	reg [31:0] eq_259_in1;
	wire [0:0] eq_259_out;
	eq #(.WIDTH(32)) eq_259(.in0(eq_259_in0), .in1(eq_259_in1), .out(eq_259_out));

	reg [0:0] andOp_260_in0;
	reg [0:0] andOp_260_in1;
	wire [0:0] andOp_260_out;
	andOp #(.WIDTH(1)) andOp_260(.in0(andOp_260_in0), .in1(andOp_260_in1), .out(andOp_260_out));

	reg [31:0] eq_261_in0;
	reg [31:0] eq_261_in1;
	wire [0:0] eq_261_out;
	eq #(.WIDTH(32)) eq_261(.in0(eq_261_in0), .in1(eq_261_in1), .out(eq_261_out));

	reg [0:0] andOp_262_in0;
	reg [0:0] andOp_262_in1;
	wire [0:0] andOp_262_out;
	andOp #(.WIDTH(1)) andOp_262(.in0(andOp_262_in0), .in1(andOp_262_in1), .out(andOp_262_out));

	reg [0:0] andOp_263_in0;
	reg [0:0] andOp_263_in1;
	wire [0:0] andOp_263_out;
	andOp #(.WIDTH(1)) andOp_263(.in0(andOp_263_in0), .in1(andOp_263_in1), .out(andOp_263_out));

	reg [31:0] eq_264_in0;
	reg [31:0] eq_264_in1;
	wire [0:0] eq_264_out;
	eq #(.WIDTH(32)) eq_264(.in0(eq_264_in0), .in1(eq_264_in1), .out(eq_264_out));

	reg [0:0] andOp_265_in0;
	reg [0:0] andOp_265_in1;
	wire [0:0] andOp_265_out;
	andOp #(.WIDTH(1)) andOp_265(.in0(andOp_265_in0), .in1(andOp_265_in1), .out(andOp_265_out));

	reg [0:0] notOp_266_in0;
	wire [0:0] notOp_266_out;
	notOp #(.WIDTH(1)) notOp_266(.in(notOp_266_in0), .out(notOp_266_out));

	reg [0:0] andOp_267_in0;
	reg [0:0] andOp_267_in1;
	wire [0:0] andOp_267_out;
	andOp #(.WIDTH(1)) andOp_267(.in0(andOp_267_in0), .in1(andOp_267_in1), .out(andOp_267_out));

	reg [0:0] notOp_268_in0;
	wire [0:0] notOp_268_out;
	notOp #(.WIDTH(1)) notOp_268(.in(notOp_268_in0), .out(notOp_268_out));

	reg [0:0] andOp_269_in0;
	reg [0:0] andOp_269_in1;
	wire [0:0] andOp_269_out;
	andOp #(.WIDTH(1)) andOp_269(.in0(andOp_269_in0), .in1(andOp_269_in1), .out(andOp_269_out));

	reg [0:0] notOp_270_in0;
	wire [0:0] notOp_270_out;
	notOp #(.WIDTH(1)) notOp_270(.in(notOp_270_in0), .out(notOp_270_out));

	reg [0:0] andOp_271_in0;
	reg [0:0] andOp_271_in1;
	wire [0:0] andOp_271_out;
	andOp #(.WIDTH(1)) andOp_271(.in0(andOp_271_in0), .in1(andOp_271_in1), .out(andOp_271_out));

	reg [0:0] andOp_272_in0;
	reg [0:0] andOp_272_in1;
	wire [0:0] andOp_272_out;
	andOp #(.WIDTH(1)) andOp_272(.in0(andOp_272_in0), .in1(andOp_272_in1), .out(andOp_272_out));

	reg [31:0] eq_273_in0;
	reg [31:0] eq_273_in1;
	wire [0:0] eq_273_out;
	eq #(.WIDTH(32)) eq_273(.in0(eq_273_in0), .in1(eq_273_in1), .out(eq_273_out));

	reg [0:0] andOp_274_in0;
	reg [0:0] andOp_274_in1;
	wire [0:0] andOp_274_out;
	andOp #(.WIDTH(1)) andOp_274(.in0(andOp_274_in0), .in1(andOp_274_in1), .out(andOp_274_out));

	reg [0:0] notOp_275_in0;
	wire [0:0] notOp_275_out;
	notOp #(.WIDTH(1)) notOp_275(.in(notOp_275_in0), .out(notOp_275_out));

	reg [0:0] andOp_276_in0;
	reg [0:0] andOp_276_in1;
	wire [0:0] andOp_276_out;
	andOp #(.WIDTH(1)) andOp_276(.in0(andOp_276_in0), .in1(andOp_276_in1), .out(andOp_276_out));

	reg [0:0] notOp_277_in0;
	wire [0:0] notOp_277_out;
	notOp #(.WIDTH(1)) notOp_277(.in(notOp_277_in0), .out(notOp_277_out));

	reg [0:0] andOp_278_in0;
	reg [0:0] andOp_278_in1;
	wire [0:0] andOp_278_out;
	andOp #(.WIDTH(1)) andOp_278(.in0(andOp_278_in0), .in1(andOp_278_in1), .out(andOp_278_out));

	reg [0:0] notOp_279_in0;
	wire [0:0] notOp_279_out;
	notOp #(.WIDTH(1)) notOp_279(.in(notOp_279_in0), .out(notOp_279_out));

	reg [0:0] andOp_280_in0;
	reg [0:0] andOp_280_in1;
	wire [0:0] andOp_280_out;
	andOp #(.WIDTH(1)) andOp_280(.in0(andOp_280_in0), .in1(andOp_280_in1), .out(andOp_280_out));

	reg [0:0] andOp_281_in0;
	reg [0:0] andOp_281_in1;
	wire [0:0] andOp_281_out;
	andOp #(.WIDTH(1)) andOp_281(.in0(andOp_281_in0), .in1(andOp_281_in1), .out(andOp_281_out));

	reg [31:0] eq_282_in0;
	reg [31:0] eq_282_in1;
	wire [0:0] eq_282_out;
	eq #(.WIDTH(32)) eq_282(.in0(eq_282_in0), .in1(eq_282_in1), .out(eq_282_out));

	reg [0:0] andOp_283_in0;
	reg [0:0] andOp_283_in1;
	wire [0:0] andOp_283_out;
	andOp #(.WIDTH(1)) andOp_283(.in0(andOp_283_in0), .in1(andOp_283_in1), .out(andOp_283_out));

	reg [0:0] notOp_284_in0;
	wire [0:0] notOp_284_out;
	notOp #(.WIDTH(1)) notOp_284(.in(notOp_284_in0), .out(notOp_284_out));

	reg [0:0] andOp_285_in0;
	reg [0:0] andOp_285_in1;
	wire [0:0] andOp_285_out;
	andOp #(.WIDTH(1)) andOp_285(.in0(andOp_285_in0), .in1(andOp_285_in1), .out(andOp_285_out));

	reg [0:0] notOp_286_in0;
	wire [0:0] notOp_286_out;
	notOp #(.WIDTH(1)) notOp_286(.in(notOp_286_in0), .out(notOp_286_out));

	reg [0:0] andOp_287_in0;
	reg [0:0] andOp_287_in1;
	wire [0:0] andOp_287_out;
	andOp #(.WIDTH(1)) andOp_287(.in0(andOp_287_in0), .in1(andOp_287_in1), .out(andOp_287_out));

	reg [0:0] notOp_288_in0;
	wire [0:0] notOp_288_out;
	notOp #(.WIDTH(1)) notOp_288(.in(notOp_288_in0), .out(notOp_288_out));

	reg [0:0] andOp_289_in0;
	reg [0:0] andOp_289_in1;
	wire [0:0] andOp_289_out;
	andOp #(.WIDTH(1)) andOp_289(.in0(andOp_289_in0), .in1(andOp_289_in1), .out(andOp_289_out));

	reg [0:0] andOp_290_in0;
	reg [0:0] andOp_290_in1;
	wire [0:0] andOp_290_out;
	andOp #(.WIDTH(1)) andOp_290(.in0(andOp_290_in0), .in1(andOp_290_in1), .out(andOp_290_out));

	reg [31:0] eq_291_in0;
	reg [31:0] eq_291_in1;
	wire [0:0] eq_291_out;
	eq #(.WIDTH(32)) eq_291(.in0(eq_291_in0), .in1(eq_291_in1), .out(eq_291_out));

	reg [0:0] andOp_292_in0;
	reg [0:0] andOp_292_in1;
	wire [0:0] andOp_292_out;
	andOp #(.WIDTH(1)) andOp_292(.in0(andOp_292_in0), .in1(andOp_292_in1), .out(andOp_292_out));

	reg [0:0] notOp_293_in0;
	wire [0:0] notOp_293_out;
	notOp #(.WIDTH(1)) notOp_293(.in(notOp_293_in0), .out(notOp_293_out));

	reg [0:0] andOp_294_in0;
	reg [0:0] andOp_294_in1;
	wire [0:0] andOp_294_out;
	andOp #(.WIDTH(1)) andOp_294(.in0(andOp_294_in0), .in1(andOp_294_in1), .out(andOp_294_out));

	reg [0:0] notOp_295_in0;
	wire [0:0] notOp_295_out;
	notOp #(.WIDTH(1)) notOp_295(.in(notOp_295_in0), .out(notOp_295_out));

	reg [0:0] andOp_296_in0;
	reg [0:0] andOp_296_in1;
	wire [0:0] andOp_296_out;
	andOp #(.WIDTH(1)) andOp_296(.in0(andOp_296_in0), .in1(andOp_296_in1), .out(andOp_296_out));

	reg [0:0] notOp_297_in0;
	wire [0:0] notOp_297_out;
	notOp #(.WIDTH(1)) notOp_297(.in(notOp_297_in0), .out(notOp_297_out));

	reg [0:0] andOp_298_in0;
	reg [0:0] andOp_298_in1;
	wire [0:0] andOp_298_out;
	andOp #(.WIDTH(1)) andOp_298(.in0(andOp_298_in0), .in1(andOp_298_in1), .out(andOp_298_out));

	reg [0:0] andOp_299_in0;
	reg [0:0] andOp_299_in1;
	wire [0:0] andOp_299_out;
	andOp #(.WIDTH(1)) andOp_299(.in0(andOp_299_in0), .in1(andOp_299_in1), .out(andOp_299_out));

	reg [31:0] eq_300_in0;
	reg [31:0] eq_300_in1;
	wire [0:0] eq_300_out;
	eq #(.WIDTH(32)) eq_300(.in0(eq_300_in0), .in1(eq_300_in1), .out(eq_300_out));

	reg [0:0] andOp_301_in0;
	reg [0:0] andOp_301_in1;
	wire [0:0] andOp_301_out;
	andOp #(.WIDTH(1)) andOp_301(.in0(andOp_301_in0), .in1(andOp_301_in1), .out(andOp_301_out));

	reg [0:0] notOp_302_in0;
	wire [0:0] notOp_302_out;
	notOp #(.WIDTH(1)) notOp_302(.in(notOp_302_in0), .out(notOp_302_out));

	reg [0:0] andOp_303_in0;
	reg [0:0] andOp_303_in1;
	wire [0:0] andOp_303_out;
	andOp #(.WIDTH(1)) andOp_303(.in0(andOp_303_in0), .in1(andOp_303_in1), .out(andOp_303_out));

	reg [0:0] notOp_304_in0;
	wire [0:0] notOp_304_out;
	notOp #(.WIDTH(1)) notOp_304(.in(notOp_304_in0), .out(notOp_304_out));

	reg [0:0] andOp_305_in0;
	reg [0:0] andOp_305_in1;
	wire [0:0] andOp_305_out;
	andOp #(.WIDTH(1)) andOp_305(.in0(andOp_305_in0), .in1(andOp_305_in1), .out(andOp_305_out));

	reg [0:0] notOp_306_in0;
	wire [0:0] notOp_306_out;
	notOp #(.WIDTH(1)) notOp_306(.in(notOp_306_in0), .out(notOp_306_out));

	reg [0:0] andOp_307_in0;
	reg [0:0] andOp_307_in1;
	wire [0:0] andOp_307_out;
	andOp #(.WIDTH(1)) andOp_307(.in0(andOp_307_in0), .in1(andOp_307_in1), .out(andOp_307_out));

	reg [0:0] andOp_308_in0;
	reg [0:0] andOp_308_in1;
	wire [0:0] andOp_308_out;
	andOp #(.WIDTH(1)) andOp_308(.in0(andOp_308_in0), .in1(andOp_308_in1), .out(andOp_308_out));

	reg [31:0] eq_309_in0;
	reg [31:0] eq_309_in1;
	wire [0:0] eq_309_out;
	eq #(.WIDTH(32)) eq_309(.in0(eq_309_in0), .in1(eq_309_in1), .out(eq_309_out));

	reg [0:0] andOp_310_in0;
	reg [0:0] andOp_310_in1;
	wire [0:0] andOp_310_out;
	andOp #(.WIDTH(1)) andOp_310(.in0(andOp_310_in0), .in1(andOp_310_in1), .out(andOp_310_out));

	reg [0:0] notOp_311_in0;
	wire [0:0] notOp_311_out;
	notOp #(.WIDTH(1)) notOp_311(.in(notOp_311_in0), .out(notOp_311_out));

	reg [0:0] andOp_312_in0;
	reg [0:0] andOp_312_in1;
	wire [0:0] andOp_312_out;
	andOp #(.WIDTH(1)) andOp_312(.in0(andOp_312_in0), .in1(andOp_312_in1), .out(andOp_312_out));

	reg [0:0] notOp_313_in0;
	wire [0:0] notOp_313_out;
	notOp #(.WIDTH(1)) notOp_313(.in(notOp_313_in0), .out(notOp_313_out));

	reg [0:0] andOp_314_in0;
	reg [0:0] andOp_314_in1;
	wire [0:0] andOp_314_out;
	andOp #(.WIDTH(1)) andOp_314(.in0(andOp_314_in0), .in1(andOp_314_in1), .out(andOp_314_out));

	reg [0:0] notOp_315_in0;
	wire [0:0] notOp_315_out;
	notOp #(.WIDTH(1)) notOp_315(.in(notOp_315_in0), .out(notOp_315_out));

	reg [0:0] andOp_316_in0;
	reg [0:0] andOp_316_in1;
	wire [0:0] andOp_316_out;
	andOp #(.WIDTH(1)) andOp_316(.in0(andOp_316_in0), .in1(andOp_316_in1), .out(andOp_316_out));

	reg [0:0] andOp_317_in0;
	reg [0:0] andOp_317_in1;
	wire [0:0] andOp_317_out;
	andOp #(.WIDTH(1)) andOp_317(.in0(andOp_317_in0), .in1(andOp_317_in1), .out(andOp_317_out));

	reg [31:0] eq_318_in0;
	reg [31:0] eq_318_in1;
	wire [0:0] eq_318_out;
	eq #(.WIDTH(32)) eq_318(.in0(eq_318_in0), .in1(eq_318_in1), .out(eq_318_out));

	reg [0:0] andOp_319_in0;
	reg [0:0] andOp_319_in1;
	wire [0:0] andOp_319_out;
	andOp #(.WIDTH(1)) andOp_319(.in0(andOp_319_in0), .in1(andOp_319_in1), .out(andOp_319_out));

	reg [0:0] notOp_320_in0;
	wire [0:0] notOp_320_out;
	notOp #(.WIDTH(1)) notOp_320(.in(notOp_320_in0), .out(notOp_320_out));

	reg [0:0] andOp_321_in0;
	reg [0:0] andOp_321_in1;
	wire [0:0] andOp_321_out;
	andOp #(.WIDTH(1)) andOp_321(.in0(andOp_321_in0), .in1(andOp_321_in1), .out(andOp_321_out));

	reg [0:0] notOp_322_in0;
	wire [0:0] notOp_322_out;
	notOp #(.WIDTH(1)) notOp_322(.in(notOp_322_in0), .out(notOp_322_out));

	reg [0:0] andOp_323_in0;
	reg [0:0] andOp_323_in1;
	wire [0:0] andOp_323_out;
	andOp #(.WIDTH(1)) andOp_323(.in0(andOp_323_in0), .in1(andOp_323_in1), .out(andOp_323_out));

	reg [0:0] notOp_324_in0;
	wire [0:0] notOp_324_out;
	notOp #(.WIDTH(1)) notOp_324(.in(notOp_324_in0), .out(notOp_324_out));

	reg [0:0] andOp_325_in0;
	reg [0:0] andOp_325_in1;
	wire [0:0] andOp_325_out;
	andOp #(.WIDTH(1)) andOp_325(.in0(andOp_325_in0), .in1(andOp_325_in1), .out(andOp_325_out));

	// End Functional Units

	reg [31:0] add_tmp_2;
	reg [31:0] data_store_0_0;
	reg [31:0] data_store_0_10;
	reg [0:0] data_store_0_12;
	reg [31:0] data_store_0_2;
	reg [31:0] data_store_0_4;
	reg [31:0] data_store_0_6;
	reg [31:0] data_store_0_8;
	reg [31:0] data_store_1_14;
	reg [31:0] data_store_1_16;
	reg [31:0] data_store_1_18;
	reg [31:0] data_store_1_20;
	reg [31:0] data_store_1_22;
	reg [31:0] data_store_1_24;
	reg [0:0] data_store_1_26;
	reg [31:0] data_store_2_28;
	reg [31:0] data_store_2_30;
	reg [31:0] data_store_2_32;
	reg [31:0] data_store_2_34;
	reg [31:0] data_store_2_36;
	reg [31:0] data_store_2_38;
	reg [0:0] data_store_2_40;
	reg [31:0] global_state;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;

	// controller for add_add_9.add_in0_add_9
	// controller for add_add_9.add_in1_add_9
	// Insensitive connections
	always @(*) begin
		add_in0_add_9 = valid ? phi_out_phi_8 : phi_out_phi_8;
		add_in1_add_9 = valid ? 32'd1 : 32'd1;
	end
	// controller for andOp_101.andOp_101_in0
	// controller for andOp_101.andOp_101_in1
	// Insensitive connections
	always @(*) begin
		andOp_101_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_101_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_102.andOp_102_in0
	// controller for andOp_102.andOp_102_in1
	// Insensitive connections
	always @(*) begin
		andOp_102_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_102_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_103.andOp_103_in0
	// controller for andOp_103.andOp_103_in1
	// Insensitive connections
	always @(*) begin
		andOp_103_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_103_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_104.andOp_104_in0
	// controller for andOp_104.andOp_104_in1
	// Insensitive connections
	always @(*) begin
		andOp_104_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_104_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_105.andOp_105_in0
	// controller for andOp_105.andOp_105_in1
	// Insensitive connections
	always @(*) begin
		andOp_105_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_105_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_106.andOp_106_in0
	// controller for andOp_106.andOp_106_in1
	// Insensitive connections
	always @(*) begin
		andOp_106_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_106_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_107.andOp_107_in0
	// controller for andOp_107.andOp_107_in1
	// Insensitive connections
	always @(*) begin
		andOp_107_in0 = valid ? bb_2_active_in_state_0_out_data : bb_2_active_in_state_0_out_data;
		andOp_107_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_108.andOp_108_in0
	// controller for andOp_108.andOp_108_in1
	// Insensitive connections
	always @(*) begin
		andOp_108_in0 = valid ? bb_2_active_in_state_1_out_data : bb_2_active_in_state_1_out_data;
		andOp_108_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_109.andOp_109_in0
	// controller for andOp_109.andOp_109_in1
	// Insensitive connections
	always @(*) begin
		andOp_109_in0 = valid ? bb_1_active_in_state_2_out_data : bb_1_active_in_state_2_out_data;
		andOp_109_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_111.andOp_111_in0
	// controller for andOp_111.andOp_111_in1
	// Insensitive connections
	always @(*) begin
		andOp_111_in0 = valid ? notOp_110_out : notOp_110_out;
		andOp_111_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_113.andOp_113_in0
	// controller for andOp_113.andOp_113_in1
	// Insensitive connections
	always @(*) begin
		andOp_113_in0 = valid ? notOp_112_out : notOp_112_out;
		andOp_113_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_115.andOp_115_in0
	// controller for andOp_115.andOp_115_in1
	// Insensitive connections
	always @(*) begin
		andOp_115_in0 = valid ? notOp_114_out : notOp_114_out;
		andOp_115_in1 = valid ? andOp_113_out : andOp_113_out;
	end
	// controller for andOp_117.andOp_117_in0
	// controller for andOp_117.andOp_117_in1
	// Insensitive connections
	always @(*) begin
		andOp_117_in0 = valid ? notOp_116_out : notOp_116_out;
		andOp_117_in1 = valid ? andOp_115_out : andOp_115_out;
	end
	// controller for andOp_118.andOp_118_in0
	// controller for andOp_118.andOp_118_in1
	// Insensitive connections
	always @(*) begin
		andOp_118_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_118_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_120.andOp_120_in0
	// controller for andOp_120.andOp_120_in1
	// Insensitive connections
	always @(*) begin
		andOp_120_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_120_in1 = valid ? eq_119_out : eq_119_out;
	end
	// controller for andOp_122.andOp_122_in0
	// controller for andOp_122.andOp_122_in1
	// Insensitive connections
	always @(*) begin
		andOp_122_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_122_in1 = valid ? eq_121_out : eq_121_out;
	end
	// controller for andOp_124.andOp_124_in0
	// controller for andOp_124.andOp_124_in1
	// Insensitive connections
	always @(*) begin
		andOp_124_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_124_in1 = valid ? eq_123_out : eq_123_out;
	end
	// controller for andOp_125.andOp_125_in0
	// controller for andOp_125.andOp_125_in1
	// Insensitive connections
	always @(*) begin
		andOp_125_in0 = valid ? 1'd0 : 1'd0;
		andOp_125_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_127.andOp_127_in0
	// controller for andOp_127.andOp_127_in1
	// Insensitive connections
	always @(*) begin
		andOp_127_in0 = valid ? andOp_125_out : andOp_125_out;
		andOp_127_in1 = valid ? eq_126_out : eq_126_out;
	end
	// controller for andOp_129.andOp_129_in0
	// controller for andOp_129.andOp_129_in1
	// Insensitive connections
	always @(*) begin
		andOp_129_in0 = valid ? andOp_125_out : andOp_125_out;
		andOp_129_in1 = valid ? notOp_128_out : notOp_128_out;
	end
	// controller for andOp_131.andOp_131_in0
	// controller for andOp_131.andOp_131_in1
	// Insensitive connections
	always @(*) begin
		andOp_131_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_131_in1 = valid ? notOp_130_out : notOp_130_out;
	end
	// controller for andOp_133.andOp_133_in0
	// controller for andOp_133.andOp_133_in1
	// Insensitive connections
	always @(*) begin
		andOp_133_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_133_in1 = valid ? notOp_132_out : notOp_132_out;
	end
	// controller for andOp_134.andOp_134_in0
	// controller for andOp_134.andOp_134_in1
	// Insensitive connections
	always @(*) begin
		andOp_134_in0 = valid ? 1'd0 : 1'd0;
		andOp_134_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_136.andOp_136_in0
	// controller for andOp_136.andOp_136_in1
	// Insensitive connections
	always @(*) begin
		andOp_136_in0 = valid ? andOp_134_out : andOp_134_out;
		andOp_136_in1 = valid ? eq_135_out : eq_135_out;
	end
	// controller for andOp_138.andOp_138_in0
	// controller for andOp_138.andOp_138_in1
	// Insensitive connections
	always @(*) begin
		andOp_138_in0 = valid ? andOp_134_out : andOp_134_out;
		andOp_138_in1 = valid ? notOp_137_out : notOp_137_out;
	end
	// controller for andOp_140.andOp_140_in0
	// controller for andOp_140.andOp_140_in1
	// Insensitive connections
	always @(*) begin
		andOp_140_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_140_in1 = valid ? notOp_139_out : notOp_139_out;
	end
	// controller for andOp_142.andOp_142_in0
	// controller for andOp_142.andOp_142_in1
	// Insensitive connections
	always @(*) begin
		andOp_142_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_142_in1 = valid ? notOp_141_out : notOp_141_out;
	end
	// controller for andOp_143.andOp_143_in0
	// controller for andOp_143.andOp_143_in1
	// Insensitive connections
	always @(*) begin
		andOp_143_in0 = valid ? 1'd0 : 1'd0;
		andOp_143_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_145.andOp_145_in0
	// controller for andOp_145.andOp_145_in1
	// Insensitive connections
	always @(*) begin
		andOp_145_in0 = valid ? andOp_143_out : andOp_143_out;
		andOp_145_in1 = valid ? eq_144_out : eq_144_out;
	end
	// controller for andOp_147.andOp_147_in0
	// controller for andOp_147.andOp_147_in1
	// Insensitive connections
	always @(*) begin
		andOp_147_in0 = valid ? andOp_143_out : andOp_143_out;
		andOp_147_in1 = valid ? notOp_146_out : notOp_146_out;
	end
	// controller for andOp_149.andOp_149_in0
	// controller for andOp_149.andOp_149_in1
	// Insensitive connections
	always @(*) begin
		andOp_149_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_149_in1 = valid ? notOp_148_out : notOp_148_out;
	end
	// controller for andOp_151.andOp_151_in0
	// controller for andOp_151.andOp_151_in1
	// Insensitive connections
	always @(*) begin
		andOp_151_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_151_in1 = valid ? notOp_150_out : notOp_150_out;
	end
	// controller for andOp_152.andOp_152_in0
	// controller for andOp_152.andOp_152_in1
	// Insensitive connections
	always @(*) begin
		andOp_152_in0 = valid ? 1'd0 : 1'd0;
		andOp_152_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_154.andOp_154_in0
	// controller for andOp_154.andOp_154_in1
	// Insensitive connections
	always @(*) begin
		andOp_154_in0 = valid ? andOp_152_out : andOp_152_out;
		andOp_154_in1 = valid ? eq_153_out : eq_153_out;
	end
	// controller for andOp_156.andOp_156_in0
	// controller for andOp_156.andOp_156_in1
	// Insensitive connections
	always @(*) begin
		andOp_156_in0 = valid ? andOp_152_out : andOp_152_out;
		andOp_156_in1 = valid ? notOp_155_out : notOp_155_out;
	end
	// controller for andOp_158.andOp_158_in0
	// controller for andOp_158.andOp_158_in1
	// Insensitive connections
	always @(*) begin
		andOp_158_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_158_in1 = valid ? notOp_157_out : notOp_157_out;
	end
	// controller for andOp_160.andOp_160_in0
	// controller for andOp_160.andOp_160_in1
	// Insensitive connections
	always @(*) begin
		andOp_160_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_160_in1 = valid ? notOp_159_out : notOp_159_out;
	end
	// controller for andOp_161.andOp_161_in0
	// controller for andOp_161.andOp_161_in1
	// Insensitive connections
	always @(*) begin
		andOp_161_in0 = valid ? 1'd0 : 1'd0;
		andOp_161_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_163.andOp_163_in0
	// controller for andOp_163.andOp_163_in1
	// Insensitive connections
	always @(*) begin
		andOp_163_in0 = valid ? andOp_161_out : andOp_161_out;
		andOp_163_in1 = valid ? eq_162_out : eq_162_out;
	end
	// controller for andOp_165.andOp_165_in0
	// controller for andOp_165.andOp_165_in1
	// Insensitive connections
	always @(*) begin
		andOp_165_in0 = valid ? andOp_161_out : andOp_161_out;
		andOp_165_in1 = valid ? notOp_164_out : notOp_164_out;
	end
	// controller for andOp_167.andOp_167_in0
	// controller for andOp_167.andOp_167_in1
	// Insensitive connections
	always @(*) begin
		andOp_167_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_167_in1 = valid ? notOp_166_out : notOp_166_out;
	end
	// controller for andOp_169.andOp_169_in0
	// controller for andOp_169.andOp_169_in1
	// Insensitive connections
	always @(*) begin
		andOp_169_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_169_in1 = valid ? notOp_168_out : notOp_168_out;
	end
	// controller for andOp_170.andOp_170_in0
	// controller for andOp_170.andOp_170_in1
	// Insensitive connections
	always @(*) begin
		andOp_170_in0 = valid ? 1'd0 : 1'd0;
		andOp_170_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_172.andOp_172_in0
	// controller for andOp_172.andOp_172_in1
	// Insensitive connections
	always @(*) begin
		andOp_172_in0 = valid ? andOp_170_out : andOp_170_out;
		andOp_172_in1 = valid ? eq_171_out : eq_171_out;
	end
	// controller for andOp_174.andOp_174_in0
	// controller for andOp_174.andOp_174_in1
	// Insensitive connections
	always @(*) begin
		andOp_174_in0 = valid ? andOp_170_out : andOp_170_out;
		andOp_174_in1 = valid ? notOp_173_out : notOp_173_out;
	end
	// controller for andOp_176.andOp_176_in0
	// controller for andOp_176.andOp_176_in1
	// Insensitive connections
	always @(*) begin
		andOp_176_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_176_in1 = valid ? notOp_175_out : notOp_175_out;
	end
	// controller for andOp_178.andOp_178_in0
	// controller for andOp_178.andOp_178_in1
	// Insensitive connections
	always @(*) begin
		andOp_178_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_178_in1 = valid ? notOp_177_out : notOp_177_out;
	end
	// controller for andOp_179.andOp_179_in0
	// controller for andOp_179.andOp_179_in1
	// Insensitive connections
	always @(*) begin
		andOp_179_in0 = valid ? 1'd0 : 1'd0;
		andOp_179_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_181.andOp_181_in0
	// controller for andOp_181.andOp_181_in1
	// Insensitive connections
	always @(*) begin
		andOp_181_in0 = valid ? andOp_179_out : andOp_179_out;
		andOp_181_in1 = valid ? eq_180_out : eq_180_out;
	end
	// controller for andOp_183.andOp_183_in0
	// controller for andOp_183.andOp_183_in1
	// Insensitive connections
	always @(*) begin
		andOp_183_in0 = valid ? andOp_179_out : andOp_179_out;
		andOp_183_in1 = valid ? notOp_182_out : notOp_182_out;
	end
	// controller for andOp_185.andOp_185_in0
	// controller for andOp_185.andOp_185_in1
	// Insensitive connections
	always @(*) begin
		andOp_185_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_185_in1 = valid ? notOp_184_out : notOp_184_out;
	end
	// controller for andOp_187.andOp_187_in0
	// controller for andOp_187.andOp_187_in1
	// Insensitive connections
	always @(*) begin
		andOp_187_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_187_in1 = valid ? notOp_186_out : notOp_186_out;
	end
	// controller for andOp_189.andOp_189_in0
	// controller for andOp_189.andOp_189_in1
	// Insensitive connections
	always @(*) begin
		andOp_189_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_189_in1 = valid ? eq_188_out : eq_188_out;
	end
	// controller for andOp_191.andOp_191_in0
	// controller for andOp_191.andOp_191_in1
	// Insensitive connections
	always @(*) begin
		andOp_191_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_191_in1 = valid ? eq_190_out : eq_190_out;
	end
	// controller for andOp_193.andOp_193_in0
	// controller for andOp_193.andOp_193_in1
	// Insensitive connections
	always @(*) begin
		andOp_193_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_193_in1 = valid ? eq_192_out : eq_192_out;
	end
	// controller for andOp_194.andOp_194_in0
	// controller for andOp_194.andOp_194_in1
	// Insensitive connections
	always @(*) begin
		andOp_194_in0 = valid ? 1'd0 : 1'd0;
		andOp_194_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_196.andOp_196_in0
	// controller for andOp_196.andOp_196_in1
	// Insensitive connections
	always @(*) begin
		andOp_196_in0 = valid ? andOp_194_out : andOp_194_out;
		andOp_196_in1 = valid ? eq_195_out : eq_195_out;
	end
	// controller for andOp_198.andOp_198_in0
	// controller for andOp_198.andOp_198_in1
	// Insensitive connections
	always @(*) begin
		andOp_198_in0 = valid ? andOp_194_out : andOp_194_out;
		andOp_198_in1 = valid ? notOp_197_out : notOp_197_out;
	end
	// controller for andOp_200.andOp_200_in0
	// controller for andOp_200.andOp_200_in1
	// Insensitive connections
	always @(*) begin
		andOp_200_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_200_in1 = valid ? notOp_199_out : notOp_199_out;
	end
	// controller for andOp_202.andOp_202_in0
	// controller for andOp_202.andOp_202_in1
	// Insensitive connections
	always @(*) begin
		andOp_202_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_202_in1 = valid ? notOp_201_out : notOp_201_out;
	end
	// controller for andOp_203.andOp_203_in0
	// controller for andOp_203.andOp_203_in1
	// Insensitive connections
	always @(*) begin
		andOp_203_in0 = valid ? 1'd0 : 1'd0;
		andOp_203_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_205.andOp_205_in0
	// controller for andOp_205.andOp_205_in1
	// Insensitive connections
	always @(*) begin
		andOp_205_in0 = valid ? andOp_203_out : andOp_203_out;
		andOp_205_in1 = valid ? eq_204_out : eq_204_out;
	end
	// controller for andOp_207.andOp_207_in0
	// controller for andOp_207.andOp_207_in1
	// Insensitive connections
	always @(*) begin
		andOp_207_in0 = valid ? andOp_203_out : andOp_203_out;
		andOp_207_in1 = valid ? notOp_206_out : notOp_206_out;
	end
	// controller for andOp_209.andOp_209_in0
	// controller for andOp_209.andOp_209_in1
	// Insensitive connections
	always @(*) begin
		andOp_209_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_209_in1 = valid ? notOp_208_out : notOp_208_out;
	end
	// controller for andOp_211.andOp_211_in0
	// controller for andOp_211.andOp_211_in1
	// Insensitive connections
	always @(*) begin
		andOp_211_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_211_in1 = valid ? notOp_210_out : notOp_210_out;
	end
	// controller for andOp_212.andOp_212_in0
	// controller for andOp_212.andOp_212_in1
	// Insensitive connections
	always @(*) begin
		andOp_212_in0 = valid ? 1'd0 : 1'd0;
		andOp_212_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_214.andOp_214_in0
	// controller for andOp_214.andOp_214_in1
	// Insensitive connections
	always @(*) begin
		andOp_214_in0 = valid ? andOp_212_out : andOp_212_out;
		andOp_214_in1 = valid ? eq_213_out : eq_213_out;
	end
	// controller for andOp_216.andOp_216_in0
	// controller for andOp_216.andOp_216_in1
	// Insensitive connections
	always @(*) begin
		andOp_216_in0 = valid ? andOp_212_out : andOp_212_out;
		andOp_216_in1 = valid ? notOp_215_out : notOp_215_out;
	end
	// controller for andOp_218.andOp_218_in0
	// controller for andOp_218.andOp_218_in1
	// Insensitive connections
	always @(*) begin
		andOp_218_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_218_in1 = valid ? notOp_217_out : notOp_217_out;
	end
	// controller for andOp_220.andOp_220_in0
	// controller for andOp_220.andOp_220_in1
	// Insensitive connections
	always @(*) begin
		andOp_220_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_220_in1 = valid ? notOp_219_out : notOp_219_out;
	end
	// controller for andOp_221.andOp_221_in0
	// controller for andOp_221.andOp_221_in1
	// Insensitive connections
	always @(*) begin
		andOp_221_in0 = valid ? 1'd0 : 1'd0;
		andOp_221_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_223.andOp_223_in0
	// controller for andOp_223.andOp_223_in1
	// Insensitive connections
	always @(*) begin
		andOp_223_in0 = valid ? andOp_221_out : andOp_221_out;
		andOp_223_in1 = valid ? eq_222_out : eq_222_out;
	end
	// controller for andOp_225.andOp_225_in0
	// controller for andOp_225.andOp_225_in1
	// Insensitive connections
	always @(*) begin
		andOp_225_in0 = valid ? andOp_221_out : andOp_221_out;
		andOp_225_in1 = valid ? notOp_224_out : notOp_224_out;
	end
	// controller for andOp_227.andOp_227_in0
	// controller for andOp_227.andOp_227_in1
	// Insensitive connections
	always @(*) begin
		andOp_227_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_227_in1 = valid ? notOp_226_out : notOp_226_out;
	end
	// controller for andOp_229.andOp_229_in0
	// controller for andOp_229.andOp_229_in1
	// Insensitive connections
	always @(*) begin
		andOp_229_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_229_in1 = valid ? notOp_228_out : notOp_228_out;
	end
	// controller for andOp_230.andOp_230_in0
	// controller for andOp_230.andOp_230_in1
	// Insensitive connections
	always @(*) begin
		andOp_230_in0 = valid ? 1'd0 : 1'd0;
		andOp_230_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_232.andOp_232_in0
	// controller for andOp_232.andOp_232_in1
	// Insensitive connections
	always @(*) begin
		andOp_232_in0 = valid ? andOp_230_out : andOp_230_out;
		andOp_232_in1 = valid ? eq_231_out : eq_231_out;
	end
	// controller for andOp_234.andOp_234_in0
	// controller for andOp_234.andOp_234_in1
	// Insensitive connections
	always @(*) begin
		andOp_234_in0 = valid ? andOp_230_out : andOp_230_out;
		andOp_234_in1 = valid ? notOp_233_out : notOp_233_out;
	end
	// controller for andOp_236.andOp_236_in0
	// controller for andOp_236.andOp_236_in1
	// Insensitive connections
	always @(*) begin
		andOp_236_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_236_in1 = valid ? notOp_235_out : notOp_235_out;
	end
	// controller for andOp_238.andOp_238_in0
	// controller for andOp_238.andOp_238_in1
	// Insensitive connections
	always @(*) begin
		andOp_238_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_238_in1 = valid ? notOp_237_out : notOp_237_out;
	end
	// controller for andOp_239.andOp_239_in0
	// controller for andOp_239.andOp_239_in1
	// Insensitive connections
	always @(*) begin
		andOp_239_in0 = valid ? 1'd0 : 1'd0;
		andOp_239_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_241.andOp_241_in0
	// controller for andOp_241.andOp_241_in1
	// Insensitive connections
	always @(*) begin
		andOp_241_in0 = valid ? andOp_239_out : andOp_239_out;
		andOp_241_in1 = valid ? eq_240_out : eq_240_out;
	end
	// controller for andOp_243.andOp_243_in0
	// controller for andOp_243.andOp_243_in1
	// Insensitive connections
	always @(*) begin
		andOp_243_in0 = valid ? andOp_239_out : andOp_239_out;
		andOp_243_in1 = valid ? notOp_242_out : notOp_242_out;
	end
	// controller for andOp_245.andOp_245_in0
	// controller for andOp_245.andOp_245_in1
	// Insensitive connections
	always @(*) begin
		andOp_245_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_245_in1 = valid ? notOp_244_out : notOp_244_out;
	end
	// controller for andOp_247.andOp_247_in0
	// controller for andOp_247.andOp_247_in1
	// Insensitive connections
	always @(*) begin
		andOp_247_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_247_in1 = valid ? notOp_246_out : notOp_246_out;
	end
	// controller for andOp_248.andOp_248_in0
	// controller for andOp_248.andOp_248_in1
	// Insensitive connections
	always @(*) begin
		andOp_248_in0 = valid ? 1'd0 : 1'd0;
		andOp_248_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_250.andOp_250_in0
	// controller for andOp_250.andOp_250_in1
	// Insensitive connections
	always @(*) begin
		andOp_250_in0 = valid ? andOp_248_out : andOp_248_out;
		andOp_250_in1 = valid ? eq_249_out : eq_249_out;
	end
	// controller for andOp_252.andOp_252_in0
	// controller for andOp_252.andOp_252_in1
	// Insensitive connections
	always @(*) begin
		andOp_252_in0 = valid ? andOp_248_out : andOp_248_out;
		andOp_252_in1 = valid ? notOp_251_out : notOp_251_out;
	end
	// controller for andOp_254.andOp_254_in0
	// controller for andOp_254.andOp_254_in1
	// Insensitive connections
	always @(*) begin
		andOp_254_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_254_in1 = valid ? notOp_253_out : notOp_253_out;
	end
	// controller for andOp_256.andOp_256_in0
	// controller for andOp_256.andOp_256_in1
	// Insensitive connections
	always @(*) begin
		andOp_256_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_256_in1 = valid ? notOp_255_out : notOp_255_out;
	end
	// controller for andOp_258.andOp_258_in0
	// controller for andOp_258.andOp_258_in1
	// Insensitive connections
	always @(*) begin
		andOp_258_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_258_in1 = valid ? eq_257_out : eq_257_out;
	end
	// controller for andOp_260.andOp_260_in0
	// controller for andOp_260.andOp_260_in1
	// Insensitive connections
	always @(*) begin
		andOp_260_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_260_in1 = valid ? eq_259_out : eq_259_out;
	end
	// controller for andOp_262.andOp_262_in0
	// controller for andOp_262.andOp_262_in1
	// Insensitive connections
	always @(*) begin
		andOp_262_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_262_in1 = valid ? eq_261_out : eq_261_out;
	end
	// controller for andOp_263.andOp_263_in0
	// controller for andOp_263.andOp_263_in1
	// Insensitive connections
	always @(*) begin
		andOp_263_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_263_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_265.andOp_265_in0
	// controller for andOp_265.andOp_265_in1
	// Insensitive connections
	always @(*) begin
		andOp_265_in0 = valid ? andOp_263_out : andOp_263_out;
		andOp_265_in1 = valid ? eq_264_out : eq_264_out;
	end
	// controller for andOp_267.andOp_267_in0
	// controller for andOp_267.andOp_267_in1
	// Insensitive connections
	always @(*) begin
		andOp_267_in0 = valid ? andOp_263_out : andOp_263_out;
		andOp_267_in1 = valid ? notOp_266_out : notOp_266_out;
	end
	// controller for andOp_269.andOp_269_in0
	// controller for andOp_269.andOp_269_in1
	// Insensitive connections
	always @(*) begin
		andOp_269_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_269_in1 = valid ? notOp_268_out : notOp_268_out;
	end
	// controller for andOp_271.andOp_271_in0
	// controller for andOp_271.andOp_271_in1
	// Insensitive connections
	always @(*) begin
		andOp_271_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_271_in1 = valid ? notOp_270_out : notOp_270_out;
	end
	// controller for andOp_272.andOp_272_in0
	// controller for andOp_272.andOp_272_in1
	// Insensitive connections
	always @(*) begin
		andOp_272_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_272_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_274.andOp_274_in0
	// controller for andOp_274.andOp_274_in1
	// Insensitive connections
	always @(*) begin
		andOp_274_in0 = valid ? andOp_272_out : andOp_272_out;
		andOp_274_in1 = valid ? eq_273_out : eq_273_out;
	end
	// controller for andOp_276.andOp_276_in0
	// controller for andOp_276.andOp_276_in1
	// Insensitive connections
	always @(*) begin
		andOp_276_in0 = valid ? andOp_272_out : andOp_272_out;
		andOp_276_in1 = valid ? notOp_275_out : notOp_275_out;
	end
	// controller for andOp_278.andOp_278_in0
	// controller for andOp_278.andOp_278_in1
	// Insensitive connections
	always @(*) begin
		andOp_278_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_278_in1 = valid ? notOp_277_out : notOp_277_out;
	end
	// controller for andOp_280.andOp_280_in0
	// controller for andOp_280.andOp_280_in1
	// Insensitive connections
	always @(*) begin
		andOp_280_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_280_in1 = valid ? notOp_279_out : notOp_279_out;
	end
	// controller for andOp_281.andOp_281_in0
	// controller for andOp_281.andOp_281_in1
	// Insensitive connections
	always @(*) begin
		andOp_281_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_281_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_283.andOp_283_in0
	// controller for andOp_283.andOp_283_in1
	// Insensitive connections
	always @(*) begin
		andOp_283_in0 = valid ? andOp_281_out : andOp_281_out;
		andOp_283_in1 = valid ? eq_282_out : eq_282_out;
	end
	// controller for andOp_285.andOp_285_in0
	// controller for andOp_285.andOp_285_in1
	// Insensitive connections
	always @(*) begin
		andOp_285_in0 = valid ? andOp_281_out : andOp_281_out;
		andOp_285_in1 = valid ? notOp_284_out : notOp_284_out;
	end
	// controller for andOp_287.andOp_287_in0
	// controller for andOp_287.andOp_287_in1
	// Insensitive connections
	always @(*) begin
		andOp_287_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_287_in1 = valid ? notOp_286_out : notOp_286_out;
	end
	// controller for andOp_289.andOp_289_in0
	// controller for andOp_289.andOp_289_in1
	// Insensitive connections
	always @(*) begin
		andOp_289_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_289_in1 = valid ? notOp_288_out : notOp_288_out;
	end
	// controller for andOp_290.andOp_290_in0
	// controller for andOp_290.andOp_290_in1
	// Insensitive connections
	always @(*) begin
		andOp_290_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_290_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_292.andOp_292_in0
	// controller for andOp_292.andOp_292_in1
	// Insensitive connections
	always @(*) begin
		andOp_292_in0 = valid ? andOp_290_out : andOp_290_out;
		andOp_292_in1 = valid ? eq_291_out : eq_291_out;
	end
	// controller for andOp_294.andOp_294_in0
	// controller for andOp_294.andOp_294_in1
	// Insensitive connections
	always @(*) begin
		andOp_294_in0 = valid ? andOp_290_out : andOp_290_out;
		andOp_294_in1 = valid ? notOp_293_out : notOp_293_out;
	end
	// controller for andOp_296.andOp_296_in0
	// controller for andOp_296.andOp_296_in1
	// Insensitive connections
	always @(*) begin
		andOp_296_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_296_in1 = valid ? notOp_295_out : notOp_295_out;
	end
	// controller for andOp_298.andOp_298_in0
	// controller for andOp_298.andOp_298_in1
	// Insensitive connections
	always @(*) begin
		andOp_298_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_298_in1 = valid ? notOp_297_out : notOp_297_out;
	end
	// controller for andOp_299.andOp_299_in0
	// controller for andOp_299.andOp_299_in1
	// Insensitive connections
	always @(*) begin
		andOp_299_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_299_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_301.andOp_301_in0
	// controller for andOp_301.andOp_301_in1
	// Insensitive connections
	always @(*) begin
		andOp_301_in0 = valid ? andOp_299_out : andOp_299_out;
		andOp_301_in1 = valid ? eq_300_out : eq_300_out;
	end
	// controller for andOp_303.andOp_303_in0
	// controller for andOp_303.andOp_303_in1
	// Insensitive connections
	always @(*) begin
		andOp_303_in0 = valid ? andOp_299_out : andOp_299_out;
		andOp_303_in1 = valid ? notOp_302_out : notOp_302_out;
	end
	// controller for andOp_305.andOp_305_in0
	// controller for andOp_305.andOp_305_in1
	// Insensitive connections
	always @(*) begin
		andOp_305_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_305_in1 = valid ? notOp_304_out : notOp_304_out;
	end
	// controller for andOp_307.andOp_307_in0
	// controller for andOp_307.andOp_307_in1
	// Insensitive connections
	always @(*) begin
		andOp_307_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_307_in1 = valid ? notOp_306_out : notOp_306_out;
	end
	// controller for andOp_308.andOp_308_in0
	// controller for andOp_308.andOp_308_in1
	// Insensitive connections
	always @(*) begin
		andOp_308_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_308_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_310.andOp_310_in0
	// controller for andOp_310.andOp_310_in1
	// Insensitive connections
	always @(*) begin
		andOp_310_in0 = valid ? andOp_308_out : andOp_308_out;
		andOp_310_in1 = valid ? eq_309_out : eq_309_out;
	end
	// controller for andOp_312.andOp_312_in0
	// controller for andOp_312.andOp_312_in1
	// Insensitive connections
	always @(*) begin
		andOp_312_in0 = valid ? andOp_308_out : andOp_308_out;
		andOp_312_in1 = valid ? notOp_311_out : notOp_311_out;
	end
	// controller for andOp_314.andOp_314_in0
	// controller for andOp_314.andOp_314_in1
	// Insensitive connections
	always @(*) begin
		andOp_314_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_314_in1 = valid ? notOp_313_out : notOp_313_out;
	end
	// controller for andOp_316.andOp_316_in0
	// controller for andOp_316.andOp_316_in1
	// Insensitive connections
	always @(*) begin
		andOp_316_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_316_in1 = valid ? notOp_315_out : notOp_315_out;
	end
	// controller for andOp_317.andOp_317_in0
	// controller for andOp_317.andOp_317_in1
	// Insensitive connections
	always @(*) begin
		andOp_317_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_317_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_319.andOp_319_in0
	// controller for andOp_319.andOp_319_in1
	// Insensitive connections
	always @(*) begin
		andOp_319_in0 = valid ? andOp_317_out : andOp_317_out;
		andOp_319_in1 = valid ? eq_318_out : eq_318_out;
	end
	// controller for andOp_321.andOp_321_in0
	// controller for andOp_321.andOp_321_in1
	// Insensitive connections
	always @(*) begin
		andOp_321_in0 = valid ? andOp_317_out : andOp_317_out;
		andOp_321_in1 = valid ? notOp_320_out : notOp_320_out;
	end
	// controller for andOp_323.andOp_323_in0
	// controller for andOp_323.andOp_323_in1
	// Insensitive connections
	always @(*) begin
		andOp_323_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_323_in1 = valid ? notOp_322_out : notOp_322_out;
	end
	// controller for andOp_325.andOp_325_in0
	// controller for andOp_325.andOp_325_in1
	// Insensitive connections
	always @(*) begin
		andOp_325_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_325_in1 = valid ? notOp_324_out : notOp_324_out;
	end
	// controller for andOp_42.andOp_42_in0
	// controller for andOp_42.andOp_42_in1
	// Insensitive connections
	always @(*) begin
		andOp_42_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_42_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_43.andOp_43_in0
	// controller for andOp_43.andOp_43_in1
	// Insensitive connections
	always @(*) begin
		andOp_43_in0 = valid ? andOp_42_out : andOp_42_out;
		andOp_43_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_45.andOp_45_in0
	// controller for andOp_45.andOp_45_in1
	// Insensitive connections
	always @(*) begin
		andOp_45_in0 = valid ? bb_2_active_in_state_2_out_data : bb_2_active_in_state_2_out_data;
		andOp_45_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_46.andOp_46_in0
	// controller for andOp_46.andOp_46_in1
	// Insensitive connections
	always @(*) begin
		andOp_46_in0 = valid ? andOp_45_out : andOp_45_out;
		andOp_46_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_48.andOp_48_in0
	// controller for andOp_48.andOp_48_in1
	// Insensitive connections
	always @(*) begin
		andOp_48_in0 = valid ? bb_2_active_in_state_2_out_data : bb_2_active_in_state_2_out_data;
		andOp_48_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_49.andOp_49_in0
	// controller for andOp_49.andOp_49_in1
	// Insensitive connections
	always @(*) begin
		andOp_49_in0 = valid ? andOp_48_out : andOp_48_out;
		andOp_49_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_51.andOp_51_in0
	// controller for andOp_51.andOp_51_in1
	// Insensitive connections
	always @(*) begin
		andOp_51_in0 = valid ? bb_2_active_in_state_2_out_data : bb_2_active_in_state_2_out_data;
		andOp_51_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_52.andOp_52_in0
	// controller for andOp_52.andOp_52_in1
	// Insensitive connections
	always @(*) begin
		andOp_52_in0 = valid ? andOp_51_out : andOp_51_out;
		andOp_52_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_54.andOp_54_in0
	// controller for andOp_54.andOp_54_in1
	// Insensitive connections
	always @(*) begin
		andOp_54_in0 = valid ? bb_3_active_in_state_2_out_data : bb_3_active_in_state_2_out_data;
		andOp_54_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_55.andOp_55_in0
	// controller for andOp_55.andOp_55_in1
	// Insensitive connections
	always @(*) begin
		andOp_55_in0 = valid ? andOp_54_out : andOp_54_out;
		andOp_55_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_57.andOp_57_in0
	// controller for andOp_57.andOp_57_in1
	// Insensitive connections
	always @(*) begin
		andOp_57_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_57_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_58.andOp_58_in0
	// controller for andOp_58.andOp_58_in1
	// Insensitive connections
	always @(*) begin
		andOp_58_in0 = valid ? andOp_57_out : andOp_57_out;
		andOp_58_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_60.andOp_60_in0
	// controller for andOp_60.andOp_60_in1
	// Insensitive connections
	always @(*) begin
		andOp_60_in0 = valid ? andOp_58_out : andOp_58_out;
		andOp_60_in1 = valid ? cmp_out_icmp_18 : cmp_out_icmp_18;
	end
	// controller for andOp_62.andOp_62_in0
	// controller for andOp_62.andOp_62_in1
	// Insensitive connections
	always @(*) begin
		andOp_62_in0 = valid ? andOp_58_out : andOp_58_out;
		andOp_62_in1 = valid ? notOp_61_out : notOp_61_out;
	end
	// controller for andOp_77.andOp_77_in0
	// controller for andOp_77.andOp_77_in1
	// Insensitive connections
	always @(*) begin
		andOp_77_in0 = valid ? notOp_76_out : notOp_76_out;
		andOp_77_in1 = valid ? andOp_43_out : andOp_43_out;
	end
	// controller for andOp_81.andOp_81_in0
	// controller for andOp_81.andOp_81_in1
	// Insensitive connections
	always @(*) begin
		andOp_81_in0 = valid ? notOp_80_out : notOp_80_out;
		andOp_81_in1 = valid ? andOp_55_out : andOp_55_out;
	end
	// controller for andOp_85.andOp_85_in0
	// controller for andOp_85.andOp_85_in1
	// Insensitive connections
	always @(*) begin
		andOp_85_in0 = valid ? notOp_84_out : notOp_84_out;
		andOp_85_in1 = valid ? andOp_62_out : andOp_62_out;
	end
	// controller for andOp_88.andOp_88_in0
	// controller for andOp_88.andOp_88_in1
	// Insensitive connections
	always @(*) begin
		andOp_88_in0 = valid ? notOp_87_out : notOp_87_out;
		andOp_88_in1 = valid ? andOp_46_out : andOp_46_out;
	end
	// controller for andOp_89.andOp_89_in0
	// controller for andOp_89.andOp_89_in1
	// Insensitive connections
	always @(*) begin
		andOp_89_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_89_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_90.andOp_90_in0
	// controller for andOp_90.andOp_90_in1
	// Insensitive connections
	always @(*) begin
		andOp_90_in0 = valid ? bb_2_active_in_state_0_out_data : bb_2_active_in_state_0_out_data;
		andOp_90_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_91.andOp_91_in0
	// controller for andOp_91.andOp_91_in1
	// Insensitive connections
	always @(*) begin
		andOp_91_in0 = valid ? bb_2_active_in_state_1_out_data : bb_2_active_in_state_1_out_data;
		andOp_91_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_92.andOp_92_in0
	// controller for andOp_92.andOp_92_in1
	// Insensitive connections
	always @(*) begin
		andOp_92_in0 = valid ? bb_2_active_in_state_2_out_data : bb_2_active_in_state_2_out_data;
		andOp_92_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_93.andOp_93_in0
	// controller for andOp_93.andOp_93_in1
	// Insensitive connections
	always @(*) begin
		andOp_93_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_93_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_94.andOp_94_in0
	// controller for andOp_94.andOp_94_in1
	// Insensitive connections
	always @(*) begin
		andOp_94_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_94_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_95.andOp_95_in0
	// controller for andOp_95.andOp_95_in1
	// Insensitive connections
	always @(*) begin
		andOp_95_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_95_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_96.andOp_96_in0
	// controller for andOp_96.andOp_96_in1
	// Insensitive connections
	always @(*) begin
		andOp_96_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_96_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_97.andOp_97_in0
	// controller for andOp_97.andOp_97_in1
	// Insensitive connections
	always @(*) begin
		andOp_97_in0 = valid ? bb_1_active_in_state_2_out_data : bb_1_active_in_state_2_out_data;
		andOp_97_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_98.andOp_98_in0
	// controller for andOp_98.andOp_98_in1
	// Insensitive connections
	always @(*) begin
		andOp_98_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
		andOp_98_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_63_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_74_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_2.bb_1_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_2_in_data = orOp_68_out;
		end else begin
			bb_1_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_2.bb_1_predecessor_in_state_2_in_data
	always @(*) begin
		if (andOp_81_out) begin 
			bb_1_predecessor_in_state_2_in_data = 32'd3;
		end else if (eq_79_out) begin 
			bb_1_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_0.bb_2_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_0_in_data = orOp_65_out;
		end else begin
			bb_2_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_1.bb_2_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_1_in_data = eq_66_out;
		end else begin
			bb_2_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_2.bb_2_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_2_in_data = eq_69_out;
		end else begin
			bb_2_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_0.bb_2_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_77_out) begin 
			bb_2_predecessor_in_state_0_in_data = 32'd0;
		end else if (eq_75_out) begin 
			bb_2_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_1.bb_2_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_78_out) begin 
			bb_2_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_2.bb_2_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_82_out) begin 
			bb_2_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_2.bb_3_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_2_in_data = orOp_71_out;
		end else begin
			bb_3_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_2.bb_3_predecessor_in_state_2_in_data
	always @(*) begin
		if (andOp_85_out) begin 
			bb_3_predecessor_in_state_2_in_data = 32'd4;
		end else if (eq_83_out) begin 
			bb_3_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_2.bb_4_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_2_in_data = orOp_73_out;
		end else begin
			bb_4_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_2.bb_4_predecessor_in_state_2_in_data
	always @(*) begin
		if (andOp_88_out) begin 
			bb_4_predecessor_in_state_2_in_data = 32'd2;
		end else if (eq_86_out) begin 
			bb_4_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_43_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_44_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_2_happened_in_state_0.br_2_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_46_out) begin 
			br_2_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_47_out) begin 
			br_2_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_2_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_2_happened_in_state_1.br_2_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_49_out) begin 
			br_2_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_50_out) begin 
			br_2_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_2_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_2_happened_in_state_2.br_2_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_52_out) begin 
			br_2_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_53_out) begin 
			br_2_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_2_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_2.br_3_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_55_out) begin 
			br_3_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_56_out) begin 
			br_3_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_2.br_4_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_58_out) begin 
			br_4_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_59_out) begin 
			br_4_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_2_in_data = 0;
		end
	end
	// controller for concat_100.concat_100_in0
	// controller for concat_100.concat_100_in1
	// Insensitive connections
	always @(*) begin
		concat_100_in0 = valid ? 32'd4 : 32'd4;
		concat_100_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for concat_99.concat_99_in0
	// controller for concat_99.concat_99_in1
	// Insensitive connections
	always @(*) begin
		concat_99_in0 = valid ? data_in_2_31_out_data : data_in_2_31_out_data;
		concat_99_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for data_in_0_1.data_in_0_1_in_data
	always @(*) begin
		if (andOp_120_out) begin 
			data_in_0_1_in_data = data_store_0_0;
		end else if (andOp_122_out) begin 
			data_in_0_1_in_data = data_store_1_14;
		end else if (andOp_124_out) begin 
			data_in_0_1_in_data = data_store_2_28;
		end else begin
			data_in_0_1_in_data = 0;
		end
	end
	// controller for data_in_0_11.data_in_0_11_in_data
	always @(*) begin
		if (andOp_120_out) begin 
			data_in_0_11_in_data = data_store_0_10;
		end else if (andOp_122_out) begin 
			data_in_0_11_in_data = data_store_1_24;
		end else if (andOp_124_out) begin 
			data_in_0_11_in_data = data_store_2_38;
		end else begin
			data_in_0_11_in_data = 0;
		end
	end
	// controller for data_in_0_13.data_in_0_13_in_data
	always @(*) begin
		if (andOp_120_out) begin 
			data_in_0_13_in_data = data_store_0_12;
		end else if (andOp_122_out) begin 
			data_in_0_13_in_data = data_store_1_26;
		end else if (andOp_124_out) begin 
			data_in_0_13_in_data = data_store_2_40;
		end else begin
			data_in_0_13_in_data = 0;
		end
	end
	// controller for data_in_0_3.data_in_0_3_in_data
	always @(*) begin
		if (andOp_120_out) begin 
			data_in_0_3_in_data = data_store_0_2;
		end else if (andOp_122_out) begin 
			data_in_0_3_in_data = data_store_1_16;
		end else if (andOp_124_out) begin 
			data_in_0_3_in_data = data_store_2_30;
		end else begin
			data_in_0_3_in_data = 0;
		end
	end
	// controller for data_in_0_5.data_in_0_5_in_data
	always @(*) begin
		if (andOp_120_out) begin 
			data_in_0_5_in_data = data_store_0_4;
		end else if (andOp_122_out) begin 
			data_in_0_5_in_data = data_store_1_18;
		end else if (andOp_124_out) begin 
			data_in_0_5_in_data = data_store_2_32;
		end else begin
			data_in_0_5_in_data = 0;
		end
	end
	// controller for data_in_0_7.data_in_0_7_in_data
	always @(*) begin
		if (andOp_120_out) begin 
			data_in_0_7_in_data = data_store_0_6;
		end else if (andOp_122_out) begin 
			data_in_0_7_in_data = data_store_1_20;
		end else if (andOp_124_out) begin 
			data_in_0_7_in_data = data_store_2_34;
		end else begin
			data_in_0_7_in_data = 0;
		end
	end
	// controller for data_in_0_9.data_in_0_9_in_data
	always @(*) begin
		if (andOp_120_out) begin 
			data_in_0_9_in_data = data_store_0_8;
		end else if (andOp_122_out) begin 
			data_in_0_9_in_data = data_store_1_22;
		end else if (andOp_124_out) begin 
			data_in_0_9_in_data = data_store_2_36;
		end else begin
			data_in_0_9_in_data = 0;
		end
	end
	// controller for data_in_1_15.data_in_1_15_in_data
	always @(*) begin
		if (andOp_189_out) begin 
			data_in_1_15_in_data = data_store_0_0;
		end else if (andOp_191_out) begin 
			data_in_1_15_in_data = data_store_1_14;
		end else if (andOp_193_out) begin 
			data_in_1_15_in_data = data_store_2_28;
		end else begin
			data_in_1_15_in_data = 0;
		end
	end
	// controller for data_in_1_17.data_in_1_17_in_data
	always @(*) begin
		if (andOp_189_out) begin 
			data_in_1_17_in_data = data_store_0_2;
		end else if (andOp_191_out) begin 
			data_in_1_17_in_data = data_store_1_16;
		end else if (andOp_193_out) begin 
			data_in_1_17_in_data = data_store_2_30;
		end else begin
			data_in_1_17_in_data = 0;
		end
	end
	// controller for data_in_1_19.data_in_1_19_in_data
	always @(*) begin
		if (andOp_189_out) begin 
			data_in_1_19_in_data = data_store_0_4;
		end else if (andOp_191_out) begin 
			data_in_1_19_in_data = data_store_1_18;
		end else if (andOp_193_out) begin 
			data_in_1_19_in_data = data_store_2_32;
		end else begin
			data_in_1_19_in_data = 0;
		end
	end
	// controller for data_in_1_21.data_in_1_21_in_data
	always @(*) begin
		if (andOp_189_out) begin 
			data_in_1_21_in_data = data_store_0_6;
		end else if (andOp_191_out) begin 
			data_in_1_21_in_data = data_store_1_20;
		end else if (andOp_193_out) begin 
			data_in_1_21_in_data = data_store_2_34;
		end else begin
			data_in_1_21_in_data = 0;
		end
	end
	// controller for data_in_1_23.data_in_1_23_in_data
	always @(*) begin
		if (andOp_189_out) begin 
			data_in_1_23_in_data = data_store_0_8;
		end else if (andOp_191_out) begin 
			data_in_1_23_in_data = data_store_1_22;
		end else if (andOp_193_out) begin 
			data_in_1_23_in_data = data_store_2_36;
		end else begin
			data_in_1_23_in_data = 0;
		end
	end
	// controller for data_in_1_25.data_in_1_25_in_data
	always @(*) begin
		if (andOp_189_out) begin 
			data_in_1_25_in_data = data_store_0_10;
		end else if (andOp_191_out) begin 
			data_in_1_25_in_data = data_store_1_24;
		end else if (andOp_193_out) begin 
			data_in_1_25_in_data = data_store_2_38;
		end else begin
			data_in_1_25_in_data = 0;
		end
	end
	// controller for data_in_1_27.data_in_1_27_in_data
	always @(*) begin
		if (andOp_189_out) begin 
			data_in_1_27_in_data = data_store_0_12;
		end else if (andOp_191_out) begin 
			data_in_1_27_in_data = data_store_1_26;
		end else if (andOp_193_out) begin 
			data_in_1_27_in_data = data_store_2_40;
		end else begin
			data_in_1_27_in_data = 0;
		end
	end
	// controller for data_in_2_29.data_in_2_29_in_data
	always @(*) begin
		if (andOp_258_out) begin 
			data_in_2_29_in_data = data_store_0_0;
		end else if (andOp_260_out) begin 
			data_in_2_29_in_data = data_store_1_14;
		end else if (andOp_262_out) begin 
			data_in_2_29_in_data = data_store_2_28;
		end else begin
			data_in_2_29_in_data = 0;
		end
	end
	// controller for data_in_2_31.data_in_2_31_in_data
	always @(*) begin
		if (andOp_258_out) begin 
			data_in_2_31_in_data = data_store_0_2;
		end else if (andOp_260_out) begin 
			data_in_2_31_in_data = data_store_1_16;
		end else if (andOp_262_out) begin 
			data_in_2_31_in_data = data_store_2_30;
		end else begin
			data_in_2_31_in_data = 0;
		end
	end
	// controller for data_in_2_33.data_in_2_33_in_data
	always @(*) begin
		if (andOp_258_out) begin 
			data_in_2_33_in_data = data_store_0_4;
		end else if (andOp_260_out) begin 
			data_in_2_33_in_data = data_store_1_18;
		end else if (andOp_262_out) begin 
			data_in_2_33_in_data = data_store_2_32;
		end else begin
			data_in_2_33_in_data = 0;
		end
	end
	// controller for data_in_2_35.data_in_2_35_in_data
	always @(*) begin
		if (andOp_258_out) begin 
			data_in_2_35_in_data = data_store_0_6;
		end else if (andOp_260_out) begin 
			data_in_2_35_in_data = data_store_1_20;
		end else if (andOp_262_out) begin 
			data_in_2_35_in_data = data_store_2_34;
		end else begin
			data_in_2_35_in_data = 0;
		end
	end
	// controller for data_in_2_37.data_in_2_37_in_data
	always @(*) begin
		if (andOp_258_out) begin 
			data_in_2_37_in_data = data_store_0_8;
		end else if (andOp_260_out) begin 
			data_in_2_37_in_data = data_store_1_22;
		end else if (andOp_262_out) begin 
			data_in_2_37_in_data = data_store_2_36;
		end else begin
			data_in_2_37_in_data = 0;
		end
	end
	// controller for data_in_2_39.data_in_2_39_in_data
	always @(*) begin
		if (andOp_258_out) begin 
			data_in_2_39_in_data = data_store_0_10;
		end else if (andOp_260_out) begin 
			data_in_2_39_in_data = data_store_1_24;
		end else if (andOp_262_out) begin 
			data_in_2_39_in_data = data_store_2_38;
		end else begin
			data_in_2_39_in_data = 0;
		end
	end
	// controller for data_in_2_41.data_in_2_41_in_data
	always @(*) begin
		if (andOp_258_out) begin 
			data_in_2_41_in_data = data_store_0_12;
		end else if (andOp_260_out) begin 
			data_in_2_41_in_data = data_store_1_26;
		end else if (andOp_262_out) begin 
			data_in_2_41_in_data = data_store_2_40;
		end else begin
			data_in_2_41_in_data = 0;
		end
	end
	// controller for eq_119.eq_119_in0
	// controller for eq_119.eq_119_in1
	// Insensitive connections
	always @(*) begin
		eq_119_in0 = valid ? 32'd0 : 32'd0;
		eq_119_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_121.eq_121_in0
	// controller for eq_121.eq_121_in1
	// Insensitive connections
	always @(*) begin
		eq_121_in0 = valid ? 32'd1 : 32'd1;
		eq_121_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_123.eq_123_in0
	// controller for eq_123.eq_123_in1
	// Insensitive connections
	always @(*) begin
		eq_123_in0 = valid ? 32'd2 : 32'd2;
		eq_123_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_126.eq_126_in0
	// controller for eq_126.eq_126_in1
	// Insensitive connections
	always @(*) begin
		eq_126_in0 = valid ? 32'd2 : 32'd2;
		eq_126_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_135.eq_135_in0
	// controller for eq_135.eq_135_in1
	// Insensitive connections
	always @(*) begin
		eq_135_in0 = valid ? 32'd2 : 32'd2;
		eq_135_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_144.eq_144_in0
	// controller for eq_144.eq_144_in1
	// Insensitive connections
	always @(*) begin
		eq_144_in0 = valid ? 32'd2 : 32'd2;
		eq_144_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_153.eq_153_in0
	// controller for eq_153.eq_153_in1
	// Insensitive connections
	always @(*) begin
		eq_153_in0 = valid ? 32'd2 : 32'd2;
		eq_153_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_162.eq_162_in0
	// controller for eq_162.eq_162_in1
	// Insensitive connections
	always @(*) begin
		eq_162_in0 = valid ? 32'd2 : 32'd2;
		eq_162_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_171.eq_171_in0
	// controller for eq_171.eq_171_in1
	// Insensitive connections
	always @(*) begin
		eq_171_in0 = valid ? 32'd2 : 32'd2;
		eq_171_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_180.eq_180_in0
	// controller for eq_180.eq_180_in1
	// Insensitive connections
	always @(*) begin
		eq_180_in0 = valid ? 32'd2 : 32'd2;
		eq_180_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_188.eq_188_in0
	// controller for eq_188.eq_188_in1
	// Insensitive connections
	always @(*) begin
		eq_188_in0 = valid ? 32'd0 : 32'd0;
		eq_188_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_190.eq_190_in0
	// controller for eq_190.eq_190_in1
	// Insensitive connections
	always @(*) begin
		eq_190_in0 = valid ? 32'd1 : 32'd1;
		eq_190_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_192.eq_192_in0
	// controller for eq_192.eq_192_in1
	// Insensitive connections
	always @(*) begin
		eq_192_in0 = valid ? 32'd2 : 32'd2;
		eq_192_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_195.eq_195_in0
	// controller for eq_195.eq_195_in1
	// Insensitive connections
	always @(*) begin
		eq_195_in0 = valid ? 32'd2 : 32'd2;
		eq_195_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_204.eq_204_in0
	// controller for eq_204.eq_204_in1
	// Insensitive connections
	always @(*) begin
		eq_204_in0 = valid ? 32'd2 : 32'd2;
		eq_204_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_213.eq_213_in0
	// controller for eq_213.eq_213_in1
	// Insensitive connections
	always @(*) begin
		eq_213_in0 = valid ? 32'd2 : 32'd2;
		eq_213_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_222.eq_222_in0
	// controller for eq_222.eq_222_in1
	// Insensitive connections
	always @(*) begin
		eq_222_in0 = valid ? 32'd2 : 32'd2;
		eq_222_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_231.eq_231_in0
	// controller for eq_231.eq_231_in1
	// Insensitive connections
	always @(*) begin
		eq_231_in0 = valid ? 32'd2 : 32'd2;
		eq_231_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_240.eq_240_in0
	// controller for eq_240.eq_240_in1
	// Insensitive connections
	always @(*) begin
		eq_240_in0 = valid ? 32'd2 : 32'd2;
		eq_240_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_249.eq_249_in0
	// controller for eq_249.eq_249_in1
	// Insensitive connections
	always @(*) begin
		eq_249_in0 = valid ? 32'd2 : 32'd2;
		eq_249_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_257.eq_257_in0
	// controller for eq_257.eq_257_in1
	// Insensitive connections
	always @(*) begin
		eq_257_in0 = valid ? 32'd0 : 32'd0;
		eq_257_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_259.eq_259_in0
	// controller for eq_259.eq_259_in1
	// Insensitive connections
	always @(*) begin
		eq_259_in0 = valid ? 32'd1 : 32'd1;
		eq_259_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_261.eq_261_in0
	// controller for eq_261.eq_261_in1
	// Insensitive connections
	always @(*) begin
		eq_261_in0 = valid ? 32'd2 : 32'd2;
		eq_261_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_264.eq_264_in0
	// controller for eq_264.eq_264_in1
	// Insensitive connections
	always @(*) begin
		eq_264_in0 = valid ? 32'd2 : 32'd2;
		eq_264_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_273.eq_273_in0
	// controller for eq_273.eq_273_in1
	// Insensitive connections
	always @(*) begin
		eq_273_in0 = valid ? 32'd2 : 32'd2;
		eq_273_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_282.eq_282_in0
	// controller for eq_282.eq_282_in1
	// Insensitive connections
	always @(*) begin
		eq_282_in0 = valid ? 32'd2 : 32'd2;
		eq_282_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_291.eq_291_in0
	// controller for eq_291.eq_291_in1
	// Insensitive connections
	always @(*) begin
		eq_291_in0 = valid ? 32'd2 : 32'd2;
		eq_291_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_300.eq_300_in0
	// controller for eq_300.eq_300_in1
	// Insensitive connections
	always @(*) begin
		eq_300_in0 = valid ? 32'd2 : 32'd2;
		eq_300_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_309.eq_309_in0
	// controller for eq_309.eq_309_in1
	// Insensitive connections
	always @(*) begin
		eq_309_in0 = valid ? 32'd2 : 32'd2;
		eq_309_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_318.eq_318_in0
	// controller for eq_318.eq_318_in1
	// Insensitive connections
	always @(*) begin
		eq_318_in0 = valid ? 32'd2 : 32'd2;
		eq_318_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_63.eq_63_in0
	// controller for eq_63.eq_63_in1
	// Insensitive connections
	always @(*) begin
		eq_63_in0 = valid ? 32'd0 : 32'd0;
		eq_63_in1 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
	end
	// controller for eq_64.eq_64_in0
	// controller for eq_64.eq_64_in1
	// Insensitive connections
	always @(*) begin
		eq_64_in0 = valid ? 32'd2 : 32'd2;
		eq_64_in1 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
	end
	// controller for eq_66.eq_66_in0
	// controller for eq_66.eq_66_in1
	// Insensitive connections
	always @(*) begin
		eq_66_in0 = valid ? 32'd2 : 32'd2;
		eq_66_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_67.eq_67_in0
	// controller for eq_67.eq_67_in1
	// Insensitive connections
	always @(*) begin
		eq_67_in0 = valid ? 32'd1 : 32'd1;
		eq_67_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_69.eq_69_in0
	// controller for eq_69.eq_69_in1
	// Insensitive connections
	always @(*) begin
		eq_69_in0 = valid ? 32'd2 : 32'd2;
		eq_69_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_70.eq_70_in0
	// controller for eq_70.eq_70_in1
	// Insensitive connections
	always @(*) begin
		eq_70_in0 = valid ? 32'd3 : 32'd3;
		eq_70_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_72.eq_72_in0
	// controller for eq_72.eq_72_in1
	// Insensitive connections
	always @(*) begin
		eq_72_in0 = valid ? 32'd4 : 32'd4;
		eq_72_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_74.eq_74_in0
	// controller for eq_74.eq_74_in1
	// Insensitive connections
	always @(*) begin
		eq_74_in0 = valid ? 32'd0 : 32'd0;
		eq_74_in1 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
	end
	// controller for eq_75.eq_75_in0
	// controller for eq_75.eq_75_in1
	// Insensitive connections
	always @(*) begin
		eq_75_in0 = valid ? 32'd2 : 32'd2;
		eq_75_in1 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
	end
	// controller for eq_78.eq_78_in0
	// controller for eq_78.eq_78_in1
	// Insensitive connections
	always @(*) begin
		eq_78_in0 = valid ? 32'd2 : 32'd2;
		eq_78_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_79.eq_79_in0
	// controller for eq_79.eq_79_in1
	// Insensitive connections
	always @(*) begin
		eq_79_in0 = valid ? 32'd1 : 32'd1;
		eq_79_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_82.eq_82_in0
	// controller for eq_82.eq_82_in1
	// Insensitive connections
	always @(*) begin
		eq_82_in0 = valid ? 32'd2 : 32'd2;
		eq_82_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_83.eq_83_in0
	// controller for eq_83.eq_83_in1
	// Insensitive connections
	always @(*) begin
		eq_83_in0 = valid ? 32'd3 : 32'd3;
		eq_83_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_86.eq_86_in0
	// controller for eq_86.eq_86_in1
	// Insensitive connections
	always @(*) begin
		eq_86_in0 = valid ? 32'd4 : 32'd4;
		eq_86_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for icmp_18.cmp_in0_icmp_18
	// controller for icmp_18.cmp_in1_icmp_18
	// Insensitive connections
	always @(*) begin
		cmp_in0_icmp_18 = valid ? add_out_add_9 : add_out_add_9;
		cmp_in1_icmp_18 = valid ? 32'd8533 : 32'd8533;
	end
	// controller for m.m_rst_n
	always @(*) begin
		if (andOp_90_out) begin 
			m_rst_n = -(1'd1);
		end else if (andOp_91_out) begin 
			m_rst_n = 1'd0;
		end else if (andOp_92_out) begin 
			m_rst_n = -(1'd1);
		end else begin
			m_rst_n = 0;
		end
	end
	// controller for m.m_word0
	always @(*) begin
		if (andOp_93_out) begin 
			m_word0 = in0_out_data;
		end else begin
			m_word0 = 0;
		end
	end
	// controller for m.m_word1
	always @(*) begin
		if (andOp_94_out) begin 
			m_word1 = in1_out_data;
		end else begin
			m_word1 = 0;
		end
	end
	// controller for m.m_word2
	always @(*) begin
		if (andOp_95_out) begin 
			m_word2 = in2_out_data;
		end else begin
			m_word2 = 0;
		end
	end
	// controller for notOp_110.notOp_110_in0
	// Insensitive connections
	always @(*) begin
		notOp_110_in0 = valid ? andOp_107_out : andOp_107_out;
	end
	// controller for notOp_112.notOp_112_in0
	// Insensitive connections
	always @(*) begin
		notOp_112_in0 = valid ? andOp_108_out : andOp_108_out;
	end
	// controller for notOp_114.notOp_114_in0
	// Insensitive connections
	always @(*) begin
		notOp_114_in0 = valid ? andOp_109_out : andOp_109_out;
	end
	// controller for notOp_116.notOp_116_in0
	// Insensitive connections
	always @(*) begin
		notOp_116_in0 = valid ? andOp_60_out : andOp_60_out;
	end
	// controller for notOp_128.notOp_128_in0
	// Insensitive connections
	always @(*) begin
		notOp_128_in0 = valid ? eq_126_out : eq_126_out;
	end
	// controller for notOp_130.notOp_130_in0
	// Insensitive connections
	always @(*) begin
		notOp_130_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_132.notOp_132_in0
	// Insensitive connections
	always @(*) begin
		notOp_132_in0 = valid ? andOp_127_out : andOp_127_out;
	end
	// controller for notOp_137.notOp_137_in0
	// Insensitive connections
	always @(*) begin
		notOp_137_in0 = valid ? eq_135_out : eq_135_out;
	end
	// controller for notOp_139.notOp_139_in0
	// Insensitive connections
	always @(*) begin
		notOp_139_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_141.notOp_141_in0
	// Insensitive connections
	always @(*) begin
		notOp_141_in0 = valid ? andOp_136_out : andOp_136_out;
	end
	// controller for notOp_146.notOp_146_in0
	// Insensitive connections
	always @(*) begin
		notOp_146_in0 = valid ? eq_144_out : eq_144_out;
	end
	// controller for notOp_148.notOp_148_in0
	// Insensitive connections
	always @(*) begin
		notOp_148_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_150.notOp_150_in0
	// Insensitive connections
	always @(*) begin
		notOp_150_in0 = valid ? andOp_145_out : andOp_145_out;
	end
	// controller for notOp_155.notOp_155_in0
	// Insensitive connections
	always @(*) begin
		notOp_155_in0 = valid ? eq_153_out : eq_153_out;
	end
	// controller for notOp_157.notOp_157_in0
	// Insensitive connections
	always @(*) begin
		notOp_157_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_159.notOp_159_in0
	// Insensitive connections
	always @(*) begin
		notOp_159_in0 = valid ? andOp_154_out : andOp_154_out;
	end
	// controller for notOp_164.notOp_164_in0
	// Insensitive connections
	always @(*) begin
		notOp_164_in0 = valid ? eq_162_out : eq_162_out;
	end
	// controller for notOp_166.notOp_166_in0
	// Insensitive connections
	always @(*) begin
		notOp_166_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_168.notOp_168_in0
	// Insensitive connections
	always @(*) begin
		notOp_168_in0 = valid ? andOp_163_out : andOp_163_out;
	end
	// controller for notOp_173.notOp_173_in0
	// Insensitive connections
	always @(*) begin
		notOp_173_in0 = valid ? eq_171_out : eq_171_out;
	end
	// controller for notOp_175.notOp_175_in0
	// Insensitive connections
	always @(*) begin
		notOp_175_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_177.notOp_177_in0
	// Insensitive connections
	always @(*) begin
		notOp_177_in0 = valid ? andOp_172_out : andOp_172_out;
	end
	// controller for notOp_182.notOp_182_in0
	// Insensitive connections
	always @(*) begin
		notOp_182_in0 = valid ? eq_180_out : eq_180_out;
	end
	// controller for notOp_184.notOp_184_in0
	// Insensitive connections
	always @(*) begin
		notOp_184_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_186.notOp_186_in0
	// Insensitive connections
	always @(*) begin
		notOp_186_in0 = valid ? andOp_181_out : andOp_181_out;
	end
	// controller for notOp_197.notOp_197_in0
	// Insensitive connections
	always @(*) begin
		notOp_197_in0 = valid ? eq_195_out : eq_195_out;
	end
	// controller for notOp_199.notOp_199_in0
	// Insensitive connections
	always @(*) begin
		notOp_199_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_201.notOp_201_in0
	// Insensitive connections
	always @(*) begin
		notOp_201_in0 = valid ? andOp_196_out : andOp_196_out;
	end
	// controller for notOp_206.notOp_206_in0
	// Insensitive connections
	always @(*) begin
		notOp_206_in0 = valid ? eq_204_out : eq_204_out;
	end
	// controller for notOp_208.notOp_208_in0
	// Insensitive connections
	always @(*) begin
		notOp_208_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_210.notOp_210_in0
	// Insensitive connections
	always @(*) begin
		notOp_210_in0 = valid ? andOp_205_out : andOp_205_out;
	end
	// controller for notOp_215.notOp_215_in0
	// Insensitive connections
	always @(*) begin
		notOp_215_in0 = valid ? eq_213_out : eq_213_out;
	end
	// controller for notOp_217.notOp_217_in0
	// Insensitive connections
	always @(*) begin
		notOp_217_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_219.notOp_219_in0
	// Insensitive connections
	always @(*) begin
		notOp_219_in0 = valid ? andOp_214_out : andOp_214_out;
	end
	// controller for notOp_224.notOp_224_in0
	// Insensitive connections
	always @(*) begin
		notOp_224_in0 = valid ? eq_222_out : eq_222_out;
	end
	// controller for notOp_226.notOp_226_in0
	// Insensitive connections
	always @(*) begin
		notOp_226_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_228.notOp_228_in0
	// Insensitive connections
	always @(*) begin
		notOp_228_in0 = valid ? andOp_223_out : andOp_223_out;
	end
	// controller for notOp_233.notOp_233_in0
	// Insensitive connections
	always @(*) begin
		notOp_233_in0 = valid ? eq_231_out : eq_231_out;
	end
	// controller for notOp_235.notOp_235_in0
	// Insensitive connections
	always @(*) begin
		notOp_235_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_237.notOp_237_in0
	// Insensitive connections
	always @(*) begin
		notOp_237_in0 = valid ? andOp_232_out : andOp_232_out;
	end
	// controller for notOp_242.notOp_242_in0
	// Insensitive connections
	always @(*) begin
		notOp_242_in0 = valid ? eq_240_out : eq_240_out;
	end
	// controller for notOp_244.notOp_244_in0
	// Insensitive connections
	always @(*) begin
		notOp_244_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_246.notOp_246_in0
	// Insensitive connections
	always @(*) begin
		notOp_246_in0 = valid ? andOp_241_out : andOp_241_out;
	end
	// controller for notOp_251.notOp_251_in0
	// Insensitive connections
	always @(*) begin
		notOp_251_in0 = valid ? eq_249_out : eq_249_out;
	end
	// controller for notOp_253.notOp_253_in0
	// Insensitive connections
	always @(*) begin
		notOp_253_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_255.notOp_255_in0
	// Insensitive connections
	always @(*) begin
		notOp_255_in0 = valid ? andOp_250_out : andOp_250_out;
	end
	// controller for notOp_266.notOp_266_in0
	// Insensitive connections
	always @(*) begin
		notOp_266_in0 = valid ? eq_264_out : eq_264_out;
	end
	// controller for notOp_268.notOp_268_in0
	// Insensitive connections
	always @(*) begin
		notOp_268_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
	end
	// controller for notOp_270.notOp_270_in0
	// Insensitive connections
	always @(*) begin
		notOp_270_in0 = valid ? andOp_265_out : andOp_265_out;
	end
	// controller for notOp_275.notOp_275_in0
	// Insensitive connections
	always @(*) begin
		notOp_275_in0 = valid ? eq_273_out : eq_273_out;
	end
	// controller for notOp_277.notOp_277_in0
	// Insensitive connections
	always @(*) begin
		notOp_277_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
	end
	// controller for notOp_279.notOp_279_in0
	// Insensitive connections
	always @(*) begin
		notOp_279_in0 = valid ? andOp_274_out : andOp_274_out;
	end
	// controller for notOp_284.notOp_284_in0
	// Insensitive connections
	always @(*) begin
		notOp_284_in0 = valid ? eq_282_out : eq_282_out;
	end
	// controller for notOp_286.notOp_286_in0
	// Insensitive connections
	always @(*) begin
		notOp_286_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
	end
	// controller for notOp_288.notOp_288_in0
	// Insensitive connections
	always @(*) begin
		notOp_288_in0 = valid ? andOp_283_out : andOp_283_out;
	end
	// controller for notOp_293.notOp_293_in0
	// Insensitive connections
	always @(*) begin
		notOp_293_in0 = valid ? eq_291_out : eq_291_out;
	end
	// controller for notOp_295.notOp_295_in0
	// Insensitive connections
	always @(*) begin
		notOp_295_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
	end
	// controller for notOp_297.notOp_297_in0
	// Insensitive connections
	always @(*) begin
		notOp_297_in0 = valid ? andOp_292_out : andOp_292_out;
	end
	// controller for notOp_302.notOp_302_in0
	// Insensitive connections
	always @(*) begin
		notOp_302_in0 = valid ? eq_300_out : eq_300_out;
	end
	// controller for notOp_304.notOp_304_in0
	// Insensitive connections
	always @(*) begin
		notOp_304_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
	end
	// controller for notOp_306.notOp_306_in0
	// Insensitive connections
	always @(*) begin
		notOp_306_in0 = valid ? andOp_301_out : andOp_301_out;
	end
	// controller for notOp_311.notOp_311_in0
	// Insensitive connections
	always @(*) begin
		notOp_311_in0 = valid ? eq_309_out : eq_309_out;
	end
	// controller for notOp_313.notOp_313_in0
	// Insensitive connections
	always @(*) begin
		notOp_313_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
	end
	// controller for notOp_315.notOp_315_in0
	// Insensitive connections
	always @(*) begin
		notOp_315_in0 = valid ? andOp_310_out : andOp_310_out;
	end
	// controller for notOp_320.notOp_320_in0
	// Insensitive connections
	always @(*) begin
		notOp_320_in0 = valid ? eq_318_out : eq_318_out;
	end
	// controller for notOp_322.notOp_322_in0
	// Insensitive connections
	always @(*) begin
		notOp_322_in0 = valid ? bb_4_active_in_state_2_out_data : bb_4_active_in_state_2_out_data;
	end
	// controller for notOp_324.notOp_324_in0
	// Insensitive connections
	always @(*) begin
		notOp_324_in0 = valid ? andOp_319_out : andOp_319_out;
	end
	// controller for notOp_44.notOp_44_in0
	// Insensitive connections
	always @(*) begin
		notOp_44_in0 = valid ? andOp_43_out : andOp_43_out;
	end
	// controller for notOp_47.notOp_47_in0
	// Insensitive connections
	always @(*) begin
		notOp_47_in0 = valid ? andOp_46_out : andOp_46_out;
	end
	// controller for notOp_50.notOp_50_in0
	// Insensitive connections
	always @(*) begin
		notOp_50_in0 = valid ? andOp_49_out : andOp_49_out;
	end
	// controller for notOp_53.notOp_53_in0
	// Insensitive connections
	always @(*) begin
		notOp_53_in0 = valid ? andOp_52_out : andOp_52_out;
	end
	// controller for notOp_56.notOp_56_in0
	// Insensitive connections
	always @(*) begin
		notOp_56_in0 = valid ? andOp_55_out : andOp_55_out;
	end
	// controller for notOp_59.notOp_59_in0
	// Insensitive connections
	always @(*) begin
		notOp_59_in0 = valid ? andOp_58_out : andOp_58_out;
	end
	// controller for notOp_61.notOp_61_in0
	// Insensitive connections
	always @(*) begin
		notOp_61_in0 = valid ? cmp_out_icmp_18 : cmp_out_icmp_18;
	end
	// controller for notOp_76.notOp_76_in0
	// Insensitive connections
	always @(*) begin
		notOp_76_in0 = valid ? eq_75_out : eq_75_out;
	end
	// controller for notOp_80.notOp_80_in0
	// Insensitive connections
	always @(*) begin
		notOp_80_in0 = valid ? eq_79_out : eq_79_out;
	end
	// controller for notOp_84.notOp_84_in0
	// Insensitive connections
	always @(*) begin
		notOp_84_in0 = valid ? eq_83_out : eq_83_out;
	end
	// controller for notOp_87.notOp_87_in0
	// Insensitive connections
	always @(*) begin
		notOp_87_in0 = valid ? eq_86_out : eq_86_out;
	end
	// controller for orOp_65.orOp_65_in0
	// controller for orOp_65.orOp_65_in1
	// Insensitive connections
	always @(*) begin
		orOp_65_in0 = valid ? eq_64_out : eq_64_out;
		orOp_65_in1 = valid ? andOp_43_out : andOp_43_out;
	end
	// controller for orOp_68.orOp_68_in0
	// controller for orOp_68.orOp_68_in1
	// Insensitive connections
	always @(*) begin
		orOp_68_in0 = valid ? eq_67_out : eq_67_out;
		orOp_68_in1 = valid ? andOp_55_out : andOp_55_out;
	end
	// controller for orOp_71.orOp_71_in0
	// controller for orOp_71.orOp_71_in1
	// Insensitive connections
	always @(*) begin
		orOp_71_in0 = valid ? eq_70_out : eq_70_out;
		orOp_71_in1 = valid ? andOp_62_out : andOp_62_out;
	end
	// controller for orOp_73.orOp_73_in0
	// controller for orOp_73.orOp_73_in1
	// Insensitive connections
	always @(*) begin
		orOp_73_in0 = valid ? eq_72_out : eq_72_out;
		orOp_73_in1 = valid ? andOp_46_out : andOp_46_out;
	end
	// controller for out.out_in_data_reg
	always @(*) begin
		if (andOp_105_out) begin 
			out_in_data_reg = m_median_word;
		end else begin
			out_in_data_reg = 0;
		end
	end
	// controller for phi_8.phi_in_phi_8
	// controller for phi_8.phi_last_block_phi_8
	// controller for phi_8.phi_s_phi_8
	// Insensitive connections
	always @(*) begin
		phi_in_phi_8 = valid ? concat_99_out : concat_99_out;
		phi_last_block_phi_8 = valid ? bb_4_predecessor_in_state_2_out_data : bb_4_predecessor_in_state_2_out_data;
		phi_s_phi_8 = valid ? concat_100_out : concat_100_out;
	end
	// controller for ret_4.valid_reg
	always @(*) begin
		if (andOp_97_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			add_tmp_2 <= 0;
		end else begin
			if (andOp_118_out) begin
				add_tmp_2 <= add_out_add_9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_0 <= 0;
		end else begin
			if (andOp_127_out) begin
				data_store_0_0 <= phi_out_phi_8;
			end
			if (andOp_133_out) begin
				data_store_0_0 <= data_in_0_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_10 <= 0;
		end else begin
			if (andOp_172_out) begin
				data_store_0_10 <= m_median_word;
			end
			if (andOp_178_out) begin
				data_store_0_10 <= data_in_0_11_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_12 <= 0;
		end else begin
			if (andOp_181_out) begin
				data_store_0_12 <= cmp_out_icmp_18;
			end
			if (andOp_187_out) begin
				data_store_0_12 <= data_in_0_13_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_2 <= 0;
		end else begin
			if (andOp_136_out) begin
				data_store_0_2 <= add_out_add_9;
			end
			if (andOp_142_out) begin
				data_store_0_2 <= data_in_0_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_4 <= 0;
		end else begin
			if (andOp_145_out) begin
				data_store_0_4 <= in0_out_data;
			end
			if (andOp_151_out) begin
				data_store_0_4 <= data_in_0_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_6 <= 0;
		end else begin
			if (andOp_154_out) begin
				data_store_0_6 <= in1_out_data;
			end
			if (andOp_160_out) begin
				data_store_0_6 <= data_in_0_7_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_8 <= 0;
		end else begin
			if (andOp_163_out) begin
				data_store_0_8 <= in2_out_data;
			end
			if (andOp_169_out) begin
				data_store_0_8 <= data_in_0_9_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_14 <= 0;
		end else begin
			if (andOp_196_out) begin
				data_store_1_14 <= phi_out_phi_8;
			end
			if (andOp_202_out) begin
				data_store_1_14 <= data_in_1_15_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_16 <= 0;
		end else begin
			if (andOp_205_out) begin
				data_store_1_16 <= add_out_add_9;
			end
			if (andOp_211_out) begin
				data_store_1_16 <= data_in_1_17_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_18 <= 0;
		end else begin
			if (andOp_214_out) begin
				data_store_1_18 <= in0_out_data;
			end
			if (andOp_220_out) begin
				data_store_1_18 <= data_in_1_19_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_20 <= 0;
		end else begin
			if (andOp_223_out) begin
				data_store_1_20 <= in1_out_data;
			end
			if (andOp_229_out) begin
				data_store_1_20 <= data_in_1_21_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_22 <= 0;
		end else begin
			if (andOp_232_out) begin
				data_store_1_22 <= in2_out_data;
			end
			if (andOp_238_out) begin
				data_store_1_22 <= data_in_1_23_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_24 <= 0;
		end else begin
			if (andOp_241_out) begin
				data_store_1_24 <= m_median_word;
			end
			if (andOp_247_out) begin
				data_store_1_24 <= data_in_1_25_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_26 <= 0;
		end else begin
			if (andOp_250_out) begin
				data_store_1_26 <= cmp_out_icmp_18;
			end
			if (andOp_256_out) begin
				data_store_1_26 <= data_in_1_27_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_28 <= 0;
		end else begin
			if (andOp_265_out) begin
				data_store_2_28 <= phi_out_phi_8;
			end
			if (andOp_271_out) begin
				data_store_2_28 <= data_in_2_29_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_30 <= 0;
		end else begin
			if (andOp_274_out) begin
				data_store_2_30 <= add_out_add_9;
			end
			if (andOp_280_out) begin
				data_store_2_30 <= data_in_2_31_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_32 <= 0;
		end else begin
			if (andOp_283_out) begin
				data_store_2_32 <= in0_out_data;
			end
			if (andOp_289_out) begin
				data_store_2_32 <= data_in_2_33_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_34 <= 0;
		end else begin
			if (andOp_292_out) begin
				data_store_2_34 <= in1_out_data;
			end
			if (andOp_298_out) begin
				data_store_2_34 <= data_in_2_35_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_36 <= 0;
		end else begin
			if (andOp_301_out) begin
				data_store_2_36 <= in2_out_data;
			end
			if (andOp_307_out) begin
				data_store_2_36 <= data_in_2_37_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_38 <= 0;
		end else begin
			if (andOp_310_out) begin
				data_store_2_38 <= m_median_word;
			end
			if (andOp_316_out) begin
				data_store_2_38 <= data_in_2_39_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_40 <= 0;
		end else begin
			if (andOp_319_out) begin
				data_store_2_40 <= cmp_out_icmp_18;
			end
			if (andOp_325_out) begin
				data_store_2_40 <= data_in_2_41_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_107_out) begin
				global_state <= 32'd1;
			end
			if (andOp_108_out) begin
				global_state <= 32'd2;
			end
			if (andOp_109_out) begin
				global_state <= 32'd2;
			end
			if (andOp_60_out) begin
				global_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (1'd1) begin
				state_0_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
			if (andOp_43_out) begin
				state_0_last_BB_reg <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_107_out) begin
				state_1_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_107_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_111_out) begin
				state_1_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_107_out) begin
				state_1_last_state <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_108_out) begin
				state_2_entry_BB_reg <= 32'd2;
			end
			if (andOp_109_out) begin
				state_2_entry_BB_reg <= 32'd1;
			end
			if (andOp_60_out) begin
				state_2_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_108_out) begin
				state_2_is_active <= 1'd1;
			end
			if (andOp_109_out) begin
				state_2_is_active <= 1'd1;
			end
			if (andOp_117_out) begin
				state_2_is_active <= 1'd0;
			end
			if (andOp_60_out) begin
				state_2_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_55_out) begin
				state_2_last_BB_reg <= 32'd3;
			end
			if (andOp_60_out) begin
				state_2_last_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_108_out) begin
				state_2_last_state <= 32'd1;
			end
			if (andOp_109_out) begin
				state_2_last_state <= 32'd2;
			end
			if (andOp_60_out) begin
				state_2_last_state <= 32'd2;
			end
		end
	end

endmodule

