module matrix_add(input [0:0] clk, input [0:0] rst, output [0:0] valid, output [8:0] a_debug_addr, input [31:0] a_debug_data, output [8:0] a_debug_write_addr, output [31:0] a_debug_write_data, output [0:0] a_debug_write_en, output [8:0] a_raddr_0, input [31:0] a_rdata_0, output [0:0] a_rst, output [8:0] a_waddr_0, output [31:0] a_wdata_0, output [0:0] a_wen_0, output [8:0] b_debug_addr, input [31:0] b_debug_data, output [8:0] b_debug_write_addr, output [31:0] b_debug_write_data, output [0:0] b_debug_write_en, output [8:0] b_raddr_0, input [31:0] b_rdata_0, output [0:0] b_rst, output [8:0] b_waddr_0, output [31:0] b_wdata_0, output [0:0] b_wen_0, output [8:0] c_debug_addr, input [31:0] c_debug_data, output [8:0] c_debug_write_addr, output [31:0] c_debug_write_data, output [0:0] c_debug_write_en, output [8:0] c_raddr_0, input [31:0] c_rdata_0, output [0:0] c_rst, output [8:0] c_waddr_0, output [31:0] c_wdata_0, output [0:0] c_wen_0);

	reg [0:0] valid_reg;
	reg [8:0] a_debug_addr_reg;
	reg [8:0] a_debug_write_addr_reg;
	reg [31:0] a_debug_write_data_reg;
	reg [0:0] a_debug_write_en_reg;
	reg [8:0] a_raddr_0_reg;
	reg [0:0] a_rst_reg;
	reg [8:0] a_waddr_0_reg;
	reg [31:0] a_wdata_0_reg;
	reg [0:0] a_wen_0_reg;
	reg [8:0] b_debug_addr_reg;
	reg [8:0] b_debug_write_addr_reg;
	reg [31:0] b_debug_write_data_reg;
	reg [0:0] b_debug_write_en_reg;
	reg [8:0] b_raddr_0_reg;
	reg [0:0] b_rst_reg;
	reg [8:0] b_waddr_0_reg;
	reg [31:0] b_wdata_0_reg;
	reg [0:0] b_wen_0_reg;
	reg [8:0] c_debug_addr_reg;
	reg [8:0] c_debug_write_addr_reg;
	reg [31:0] c_debug_write_data_reg;
	reg [0:0] c_debug_write_en_reg;
	reg [8:0] c_raddr_0_reg;
	reg [0:0] c_rst_reg;
	reg [8:0] c_waddr_0_reg;
	reg [31:0] c_wdata_0_reg;
	reg [0:0] c_wen_0_reg;

	assign valid = valid_reg;
	assign a_debug_addr = a_debug_addr_reg;
	assign a_debug_write_addr = a_debug_write_addr_reg;
	assign a_debug_write_data = a_debug_write_data_reg;
	assign a_debug_write_en = a_debug_write_en_reg;
	assign a_raddr_0 = a_raddr_0_reg;
	assign a_rst = a_rst_reg;
	assign a_waddr_0 = a_waddr_0_reg;
	assign a_wdata_0 = a_wdata_0_reg;
	assign a_wen_0 = a_wen_0_reg;
	assign b_debug_addr = b_debug_addr_reg;
	assign b_debug_write_addr = b_debug_write_addr_reg;
	assign b_debug_write_data = b_debug_write_data_reg;
	assign b_debug_write_en = b_debug_write_en_reg;
	assign b_raddr_0 = b_raddr_0_reg;
	assign b_rst = b_rst_reg;
	assign b_waddr_0 = b_waddr_0_reg;
	assign b_wdata_0 = b_wdata_0_reg;
	assign b_wen_0 = b_wen_0_reg;
	assign c_debug_addr = c_debug_addr_reg;
	assign c_debug_write_addr = c_debug_write_addr_reg;
	assign c_debug_write_data = c_debug_write_data_reg;
	assign c_debug_write_en = c_debug_write_en_reg;
	assign c_raddr_0 = c_raddr_0_reg;
	assign c_rst = c_rst_reg;
	assign c_waddr_0 = c_waddr_0_reg;
	assign c_wdata_0 = c_wdata_0_reg;
	assign c_wen_0 = c_wen_0_reg;

	// Start debug wires and ports

	initial begin
	end






	// End debug wires and ports

	// Start Functional Units
	wire [31:0] add_add12_in0;
	wire [31:0] add_add12_in1;
	wire [31:0] add_add12_out;
	add #(.WIDTH(32)) add_add12(.in0(add_add12_in0), .in1(add_add12_in1), .out(add_add12_out));

	br_dummy br_unit();

	wire [31:0] add_add17_in0;
	wire [31:0] add_add17_in1;
	wire [31:0] add_add17_out;
	add #(.WIDTH(32)) add_add17(.in0(add_add17_in0), .in1(add_add17_in1), .out(add_add17_out));

	wire [31:0] shl_shl2_in0;
	wire [31:0] shl_shl2_in1;
	wire [31:0] shl_shl2_out;
	shlOp #(.WIDTH(32)) shl_shl2(.in0(shl_shl2_in0), .in1(shl_shl2_in1), .out(shl_shl2_out));

	wire [63:0] phi_phi3_in;
	wire [31:0] phi_phi3_last_block;
	wire [63:0] phi_phi3_s;
	wire [31:0] phi_phi3_out;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_phi3(.in(phi_phi3_in), .last_block(phi_phi3_last_block), .out(phi_phi3_out), .s(phi_phi3_s));

	wire [31:0] icmp_icmp18_in0;
	wire [31:0] icmp_icmp18_in1;
	wire [0:0] icmp_icmp18_out;
	eq #(.WIDTH(32)) icmp_icmp18(.in0(icmp_icmp18_in0), .in1(icmp_icmp18_in1), .out(icmp_icmp18_out));

	wire [63:0] phi_phi4_in;
	wire [31:0] phi_phi4_last_block;
	wire [63:0] phi_phi4_s;
	wire [31:0] phi_phi4_out;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_phi4(.in(phi_phi4_in), .last_block(phi_phi4_last_block), .out(phi_phi4_out), .s(phi_phi4_s));

	wire [31:0] add_add8_in0;
	wire [31:0] add_add8_in1;
	wire [31:0] add_add8_out;
	add #(.WIDTH(32)) add_add8(.in0(add_add8_in0), .in1(add_add8_in1), .out(add_add8_out));

	wire [31:0] add_add6_in0;
	wire [31:0] add_add6_in1;
	wire [31:0] add_add6_out;
	add #(.WIDTH(32)) add_add6(.in0(add_add6_in0), .in1(add_add6_in1), .out(add_add6_out));

	wire [31:0] icmp_icmp7_in0;
	wire [31:0] icmp_icmp7_in1;
	wire [0:0] icmp_icmp7_out;
	eq #(.WIDTH(32)) icmp_icmp7(.in0(icmp_icmp7_in0), .in1(icmp_icmp7_in1), .out(icmp_icmp7_out));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] bb_1_active_in_state_1_in_data;
	wire [0:0] bb_1_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_1(.in_data(bb_1_active_in_state_1_in_data), .out_data(bb_1_active_in_state_1_out_data));

	reg [31:0] bb_1_predecessor_in_state_1_in_data;
	wire [31:0] bb_1_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_1(.in_data(bb_1_predecessor_in_state_1_in_data), .out_data(bb_1_predecessor_in_state_1_out_data));

	reg [0:0] br_1_happened_in_state_1_in_data;
	wire [0:0] br_1_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened_in_state_1(.in_data(br_1_happened_in_state_1_in_data), .out_data(br_1_happened_in_state_1_out_data));

	reg [0:0] bb_4_active_in_state_1_in_data;
	wire [0:0] bb_4_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_1(.in_data(bb_4_active_in_state_1_in_data), .out_data(bb_4_active_in_state_1_out_data));

	reg [31:0] bb_4_predecessor_in_state_1_in_data;
	wire [31:0] bb_4_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_1(.in_data(bb_4_predecessor_in_state_1_in_data), .out_data(bb_4_predecessor_in_state_1_out_data));

	reg [0:0] br_4_happened_in_state_1_in_data;
	wire [0:0] br_4_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_1(.in_data(br_4_happened_in_state_1_in_data), .out_data(br_4_happened_in_state_1_out_data));

	reg [0:0] bb_4_active_in_state_2_in_data;
	wire [0:0] bb_4_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_2(.in_data(bb_4_active_in_state_2_in_data), .out_data(bb_4_active_in_state_2_out_data));

	reg [31:0] bb_4_predecessor_in_state_2_in_data;
	wire [31:0] bb_4_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_2(.in_data(bb_4_predecessor_in_state_2_in_data), .out_data(bb_4_predecessor_in_state_2_out_data));

	reg [0:0] br_4_happened_in_state_2_in_data;
	wire [0:0] br_4_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_2(.in_data(br_4_happened_in_state_2_in_data), .out_data(br_4_happened_in_state_2_out_data));

	reg [0:0] bb_4_active_in_state_3_in_data;
	wire [0:0] bb_4_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_3(.in_data(bb_4_active_in_state_3_in_data), .out_data(bb_4_active_in_state_3_out_data));

	reg [31:0] bb_4_predecessor_in_state_3_in_data;
	wire [31:0] bb_4_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_3(.in_data(bb_4_predecessor_in_state_3_in_data), .out_data(bb_4_predecessor_in_state_3_out_data));

	reg [0:0] br_4_happened_in_state_3_in_data;
	wire [0:0] br_4_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_3(.in_data(br_4_happened_in_state_3_in_data), .out_data(br_4_happened_in_state_3_out_data));

	reg [0:0] bb_4_active_in_state_4_in_data;
	wire [0:0] bb_4_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_4(.in_data(bb_4_active_in_state_4_in_data), .out_data(bb_4_active_in_state_4_out_data));

	reg [31:0] bb_4_predecessor_in_state_4_in_data;
	wire [31:0] bb_4_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_4(.in_data(bb_4_predecessor_in_state_4_in_data), .out_data(bb_4_predecessor_in_state_4_out_data));

	reg [0:0] br_4_happened_in_state_4_in_data;
	wire [0:0] br_4_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_4(.in_data(br_4_happened_in_state_4_in_data), .out_data(br_4_happened_in_state_4_out_data));

	reg [0:0] bb_4_active_in_state_5_in_data;
	wire [0:0] bb_4_active_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_5(.in_data(bb_4_active_in_state_5_in_data), .out_data(bb_4_active_in_state_5_out_data));

	reg [31:0] bb_4_predecessor_in_state_5_in_data;
	wire [31:0] bb_4_predecessor_in_state_5_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_5(.in_data(bb_4_predecessor_in_state_5_in_data), .out_data(bb_4_predecessor_in_state_5_out_data));

	reg [0:0] br_4_happened_in_state_5_in_data;
	wire [0:0] br_4_happened_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_5(.in_data(br_4_happened_in_state_5_in_data), .out_data(br_4_happened_in_state_5_out_data));

	reg [0:0] bb_4_active_in_state_6_in_data;
	wire [0:0] bb_4_active_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_6(.in_data(bb_4_active_in_state_6_in_data), .out_data(bb_4_active_in_state_6_out_data));

	reg [31:0] bb_4_predecessor_in_state_6_in_data;
	wire [31:0] bb_4_predecessor_in_state_6_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_6(.in_data(bb_4_predecessor_in_state_6_in_data), .out_data(bb_4_predecessor_in_state_6_out_data));

	reg [0:0] br_4_happened_in_state_6_in_data;
	wire [0:0] br_4_happened_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_6(.in_data(br_4_happened_in_state_6_in_data), .out_data(br_4_happened_in_state_6_out_data));

	reg [0:0] bb_3_active_in_state_7_in_data;
	wire [0:0] bb_3_active_in_state_7_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_7(.in_data(bb_3_active_in_state_7_in_data), .out_data(bb_3_active_in_state_7_out_data));

	reg [31:0] bb_3_predecessor_in_state_7_in_data;
	wire [31:0] bb_3_predecessor_in_state_7_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_7(.in_data(bb_3_predecessor_in_state_7_in_data), .out_data(bb_3_predecessor_in_state_7_out_data));

	reg [0:0] br_3_happened_in_state_7_in_data;
	wire [0:0] br_3_happened_in_state_7_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_7(.in_data(br_3_happened_in_state_7_in_data), .out_data(br_3_happened_in_state_7_out_data));

	reg [0:0] bb_4_active_in_state_7_in_data;
	wire [0:0] bb_4_active_in_state_7_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_7(.in_data(bb_4_active_in_state_7_in_data), .out_data(bb_4_active_in_state_7_out_data));

	reg [31:0] bb_4_predecessor_in_state_7_in_data;
	wire [31:0] bb_4_predecessor_in_state_7_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_7(.in_data(bb_4_predecessor_in_state_7_in_data), .out_data(bb_4_predecessor_in_state_7_out_data));

	reg [0:0] br_4_happened_in_state_7_in_data;
	wire [0:0] br_4_happened_in_state_7_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_7(.in_data(br_4_happened_in_state_7_in_data), .out_data(br_4_happened_in_state_7_out_data));

	reg [0:0] bb_2_active_in_state_8_in_data;
	wire [0:0] bb_2_active_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_8(.in_data(bb_2_active_in_state_8_in_data), .out_data(bb_2_active_in_state_8_out_data));

	reg [31:0] bb_2_predecessor_in_state_8_in_data;
	wire [31:0] bb_2_predecessor_in_state_8_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_8(.in_data(bb_2_predecessor_in_state_8_in_data), .out_data(bb_2_predecessor_in_state_8_out_data));

	reg [31:0] data_in_0_1_in_data;
	wire [31:0] data_in_0_1_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_1(.in_data(data_in_0_1_in_data), .out_data(data_in_0_1_out_data));

	reg [31:0] data_in_0_3_in_data;
	wire [31:0] data_in_0_3_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_3(.in_data(data_in_0_3_in_data), .out_data(data_in_0_3_out_data));

	reg [31:0] data_in_0_5_in_data;
	wire [31:0] data_in_0_5_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_5(.in_data(data_in_0_5_in_data), .out_data(data_in_0_5_out_data));

	reg [31:0] data_in_0_7_in_data;
	wire [31:0] data_in_0_7_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_7(.in_data(data_in_0_7_in_data), .out_data(data_in_0_7_out_data));

	reg [31:0] data_in_1_9_in_data;
	wire [31:0] data_in_1_9_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_9(.in_data(data_in_1_9_in_data), .out_data(data_in_1_9_out_data));

	reg [31:0] data_in_1_11_in_data;
	wire [31:0] data_in_1_11_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_11(.in_data(data_in_1_11_in_data), .out_data(data_in_1_11_out_data));

	reg [31:0] data_in_1_13_in_data;
	wire [31:0] data_in_1_13_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_13(.in_data(data_in_1_13_in_data), .out_data(data_in_1_13_out_data));

	reg [31:0] data_in_1_16_in_data;
	wire [31:0] data_in_1_16_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_16(.in_data(data_in_1_16_in_data), .out_data(data_in_1_16_out_data));

	reg [31:0] data_in_2_18_in_data;
	wire [31:0] data_in_2_18_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_18(.in_data(data_in_2_18_in_data), .out_data(data_in_2_18_out_data));

	reg [31:0] data_in_2_20_in_data;
	wire [31:0] data_in_2_20_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_20(.in_data(data_in_2_20_in_data), .out_data(data_in_2_20_out_data));

	reg [31:0] data_in_2_22_in_data;
	wire [31:0] data_in_2_22_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_22(.in_data(data_in_2_22_in_data), .out_data(data_in_2_22_out_data));

	reg [31:0] data_in_2_23_in_data;
	wire [31:0] data_in_2_23_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_23(.in_data(data_in_2_23_in_data), .out_data(data_in_2_23_out_data));

	reg [31:0] data_in_2_26_in_data;
	wire [31:0] data_in_2_26_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_26(.in_data(data_in_2_26_in_data), .out_data(data_in_2_26_out_data));

	reg [31:0] data_in_3_28_in_data;
	wire [31:0] data_in_3_28_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_28(.in_data(data_in_3_28_in_data), .out_data(data_in_3_28_out_data));

	reg [31:0] data_in_3_30_in_data;
	wire [31:0] data_in_3_30_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_30(.in_data(data_in_3_30_in_data), .out_data(data_in_3_30_out_data));

	reg [31:0] data_in_3_32_in_data;
	wire [31:0] data_in_3_32_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_32(.in_data(data_in_3_32_in_data), .out_data(data_in_3_32_out_data));

	reg [31:0] data_in_3_34_in_data;
	wire [31:0] data_in_3_34_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_34(.in_data(data_in_3_34_in_data), .out_data(data_in_3_34_out_data));

	reg [31:0] data_in_3_36_in_data;
	wire [31:0] data_in_3_36_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_36(.in_data(data_in_3_36_in_data), .out_data(data_in_3_36_out_data));

	reg [31:0] data_in_4_39_in_data;
	wire [31:0] data_in_4_39_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_39(.in_data(data_in_4_39_in_data), .out_data(data_in_4_39_out_data));

	reg [31:0] data_in_4_41_in_data;
	wire [31:0] data_in_4_41_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_41(.in_data(data_in_4_41_in_data), .out_data(data_in_4_41_out_data));

	reg [31:0] data_in_4_43_in_data;
	wire [31:0] data_in_4_43_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_43(.in_data(data_in_4_43_in_data), .out_data(data_in_4_43_out_data));

	reg [31:0] data_in_4_44_in_data;
	wire [31:0] data_in_4_44_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_44(.in_data(data_in_4_44_in_data), .out_data(data_in_4_44_out_data));

	reg [31:0] data_in_4_46_in_data;
	wire [31:0] data_in_4_46_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_46(.in_data(data_in_4_46_in_data), .out_data(data_in_4_46_out_data));

	reg [31:0] data_in_4_47_in_data;
	wire [31:0] data_in_4_47_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_47(.in_data(data_in_4_47_in_data), .out_data(data_in_4_47_out_data));

	reg [31:0] data_in_5_49_in_data;
	wire [31:0] data_in_5_49_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_49(.in_data(data_in_5_49_in_data), .out_data(data_in_5_49_out_data));

	reg [31:0] data_in_5_51_in_data;
	wire [31:0] data_in_5_51_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_51(.in_data(data_in_5_51_in_data), .out_data(data_in_5_51_out_data));

	reg [31:0] data_in_5_53_in_data;
	wire [31:0] data_in_5_53_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_53(.in_data(data_in_5_53_in_data), .out_data(data_in_5_53_out_data));

	reg [31:0] data_in_5_55_in_data;
	wire [31:0] data_in_5_55_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_55(.in_data(data_in_5_55_in_data), .out_data(data_in_5_55_out_data));

	reg [31:0] data_in_6_57_in_data;
	wire [31:0] data_in_6_57_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_57(.in_data(data_in_6_57_in_data), .out_data(data_in_6_57_out_data));

	reg [31:0] data_in_6_59_in_data;
	wire [31:0] data_in_6_59_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_59(.in_data(data_in_6_59_in_data), .out_data(data_in_6_59_out_data));

	reg [31:0] data_in_6_61_in_data;
	wire [31:0] data_in_6_61_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_61(.in_data(data_in_6_61_in_data), .out_data(data_in_6_61_out_data));

	reg [31:0] data_in_6_63_in_data;
	wire [31:0] data_in_6_63_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_63(.in_data(data_in_6_63_in_data), .out_data(data_in_6_63_out_data));

	reg [31:0] data_in_7_65_in_data;
	wire [31:0] data_in_7_65_out_data;
	hls_wire #(.WIDTH(32)) data_in_7_65(.in_data(data_in_7_65_in_data), .out_data(data_in_7_65_out_data));

	reg [31:0] data_in_7_67_in_data;
	wire [31:0] data_in_7_67_out_data;
	hls_wire #(.WIDTH(32)) data_in_7_67(.in_data(data_in_7_67_in_data), .out_data(data_in_7_67_out_data));

	reg [31:0] data_in_7_69_in_data;
	wire [31:0] data_in_7_69_out_data;
	hls_wire #(.WIDTH(32)) data_in_7_69(.in_data(data_in_7_69_in_data), .out_data(data_in_7_69_out_data));

	reg [31:0] data_in_7_71_in_data;
	wire [31:0] data_in_7_71_out_data;
	hls_wire #(.WIDTH(32)) data_in_7_71(.in_data(data_in_7_71_in_data), .out_data(data_in_7_71_out_data));

	wire [0:0] andOp_72_in0;
	wire [0:0] andOp_72_in1;
	wire [0:0] andOp_72_out;
	andOp #(.WIDTH(1)) andOp_72(.in0(andOp_72_in0), .in1(andOp_72_in1), .out(andOp_72_out));

	wire [0:0] notOp_73_in0;
	wire [0:0] notOp_73_out;
	notOp #(.WIDTH(1)) notOp_73(.in(notOp_73_in0), .out(notOp_73_out));

	wire [0:0] andOp_74_in0;
	wire [0:0] andOp_74_in1;
	wire [0:0] andOp_74_out;
	andOp #(.WIDTH(1)) andOp_74(.in0(andOp_74_in0), .in1(andOp_74_in1), .out(andOp_74_out));

	wire [0:0] notOp_75_in0;
	wire [0:0] notOp_75_out;
	notOp #(.WIDTH(1)) notOp_75(.in(notOp_75_in0), .out(notOp_75_out));

	wire [0:0] andOp_76_in0;
	wire [0:0] andOp_76_in1;
	wire [0:0] andOp_76_out;
	andOp #(.WIDTH(1)) andOp_76(.in0(andOp_76_in0), .in1(andOp_76_in1), .out(andOp_76_out));

	wire [0:0] notOp_77_in0;
	wire [0:0] notOp_77_out;
	notOp #(.WIDTH(1)) notOp_77(.in(notOp_77_in0), .out(notOp_77_out));

	wire [0:0] andOp_78_in0;
	wire [0:0] andOp_78_in1;
	wire [0:0] andOp_78_out;
	andOp #(.WIDTH(1)) andOp_78(.in0(andOp_78_in0), .in1(andOp_78_in1), .out(andOp_78_out));

	wire [0:0] notOp_79_in0;
	wire [0:0] notOp_79_out;
	notOp #(.WIDTH(1)) notOp_79(.in(notOp_79_in0), .out(notOp_79_out));

	wire [0:0] andOp_80_in0;
	wire [0:0] andOp_80_in1;
	wire [0:0] andOp_80_out;
	andOp #(.WIDTH(1)) andOp_80(.in0(andOp_80_in0), .in1(andOp_80_in1), .out(andOp_80_out));

	wire [0:0] andOp_81_in0;
	wire [0:0] andOp_81_in1;
	wire [0:0] andOp_81_out;
	andOp #(.WIDTH(1)) andOp_81(.in0(andOp_81_in0), .in1(andOp_81_in1), .out(andOp_81_out));

	wire [0:0] notOp_82_in0;
	wire [0:0] notOp_82_out;
	notOp #(.WIDTH(1)) notOp_82(.in(notOp_82_in0), .out(notOp_82_out));

	wire [0:0] andOp_83_in0;
	wire [0:0] andOp_83_in1;
	wire [0:0] andOp_83_out;
	andOp #(.WIDTH(1)) andOp_83(.in0(andOp_83_in0), .in1(andOp_83_in1), .out(andOp_83_out));

	wire [0:0] notOp_84_in0;
	wire [0:0] notOp_84_out;
	notOp #(.WIDTH(1)) notOp_84(.in(notOp_84_in0), .out(notOp_84_out));

	wire [0:0] andOp_85_in0;
	wire [0:0] andOp_85_in1;
	wire [0:0] andOp_85_out;
	andOp #(.WIDTH(1)) andOp_85(.in0(andOp_85_in0), .in1(andOp_85_in1), .out(andOp_85_out));

	wire [0:0] andOp_86_in0;
	wire [0:0] andOp_86_in1;
	wire [0:0] andOp_86_out;
	andOp #(.WIDTH(1)) andOp_86(.in0(andOp_86_in0), .in1(andOp_86_in1), .out(andOp_86_out));

	wire [0:0] notOp_87_in0;
	wire [0:0] notOp_87_out;
	notOp #(.WIDTH(1)) notOp_87(.in(notOp_87_in0), .out(notOp_87_out));

	wire [0:0] andOp_88_in0;
	wire [0:0] andOp_88_in1;
	wire [0:0] andOp_88_out;
	andOp #(.WIDTH(1)) andOp_88(.in0(andOp_88_in0), .in1(andOp_88_in1), .out(andOp_88_out));

	wire [0:0] notOp_89_in0;
	wire [0:0] notOp_89_out;
	notOp #(.WIDTH(1)) notOp_89(.in(notOp_89_in0), .out(notOp_89_out));

	wire [0:0] andOp_90_in0;
	wire [0:0] andOp_90_in1;
	wire [0:0] andOp_90_out;
	andOp #(.WIDTH(1)) andOp_90(.in0(andOp_90_in0), .in1(andOp_90_in1), .out(andOp_90_out));

	wire [0:0] andOp_91_in0;
	wire [0:0] andOp_91_in1;
	wire [0:0] andOp_91_out;
	andOp #(.WIDTH(1)) andOp_91(.in0(andOp_91_in0), .in1(andOp_91_in1), .out(andOp_91_out));

	wire [0:0] notOp_92_in0;
	wire [0:0] notOp_92_out;
	notOp #(.WIDTH(1)) notOp_92(.in(notOp_92_in0), .out(notOp_92_out));

	wire [0:0] andOp_93_in0;
	wire [0:0] andOp_93_in1;
	wire [0:0] andOp_93_out;
	andOp #(.WIDTH(1)) andOp_93(.in0(andOp_93_in0), .in1(andOp_93_in1), .out(andOp_93_out));

	wire [0:0] notOp_94_in0;
	wire [0:0] notOp_94_out;
	notOp #(.WIDTH(1)) notOp_94(.in(notOp_94_in0), .out(notOp_94_out));

	wire [0:0] andOp_95_in0;
	wire [0:0] andOp_95_in1;
	wire [0:0] andOp_95_out;
	andOp #(.WIDTH(1)) andOp_95(.in0(andOp_95_in0), .in1(andOp_95_in1), .out(andOp_95_out));

	wire [0:0] andOp_96_in0;
	wire [0:0] andOp_96_in1;
	wire [0:0] andOp_96_out;
	andOp #(.WIDTH(1)) andOp_96(.in0(andOp_96_in0), .in1(andOp_96_in1), .out(andOp_96_out));

	wire [0:0] notOp_97_in0;
	wire [0:0] notOp_97_out;
	notOp #(.WIDTH(1)) notOp_97(.in(notOp_97_in0), .out(notOp_97_out));

	wire [0:0] andOp_98_in0;
	wire [0:0] andOp_98_in1;
	wire [0:0] andOp_98_out;
	andOp #(.WIDTH(1)) andOp_98(.in0(andOp_98_in0), .in1(andOp_98_in1), .out(andOp_98_out));

	wire [0:0] notOp_99_in0;
	wire [0:0] notOp_99_out;
	notOp #(.WIDTH(1)) notOp_99(.in(notOp_99_in0), .out(notOp_99_out));

	wire [0:0] andOp_100_in0;
	wire [0:0] andOp_100_in1;
	wire [0:0] andOp_100_out;
	andOp #(.WIDTH(1)) andOp_100(.in0(andOp_100_in0), .in1(andOp_100_in1), .out(andOp_100_out));

	wire [0:0] andOp_101_in0;
	wire [0:0] andOp_101_in1;
	wire [0:0] andOp_101_out;
	andOp #(.WIDTH(1)) andOp_101(.in0(andOp_101_in0), .in1(andOp_101_in1), .out(andOp_101_out));

	wire [0:0] notOp_102_in0;
	wire [0:0] notOp_102_out;
	notOp #(.WIDTH(1)) notOp_102(.in(notOp_102_in0), .out(notOp_102_out));

	wire [0:0] andOp_103_in0;
	wire [0:0] andOp_103_in1;
	wire [0:0] andOp_103_out;
	andOp #(.WIDTH(1)) andOp_103(.in0(andOp_103_in0), .in1(andOp_103_in1), .out(andOp_103_out));

	wire [0:0] notOp_104_in0;
	wire [0:0] notOp_104_out;
	notOp #(.WIDTH(1)) notOp_104(.in(notOp_104_in0), .out(notOp_104_out));

	wire [0:0] andOp_105_in0;
	wire [0:0] andOp_105_in1;
	wire [0:0] andOp_105_out;
	andOp #(.WIDTH(1)) andOp_105(.in0(andOp_105_in0), .in1(andOp_105_in1), .out(andOp_105_out));

	wire [0:0] andOp_106_in0;
	wire [0:0] andOp_106_in1;
	wire [0:0] andOp_106_out;
	andOp #(.WIDTH(1)) andOp_106(.in0(andOp_106_in0), .in1(andOp_106_in1), .out(andOp_106_out));

	wire [0:0] notOp_107_in0;
	wire [0:0] notOp_107_out;
	notOp #(.WIDTH(1)) notOp_107(.in(notOp_107_in0), .out(notOp_107_out));

	wire [0:0] andOp_108_in0;
	wire [0:0] andOp_108_in1;
	wire [0:0] andOp_108_out;
	andOp #(.WIDTH(1)) andOp_108(.in0(andOp_108_in0), .in1(andOp_108_in1), .out(andOp_108_out));

	wire [0:0] notOp_109_in0;
	wire [0:0] notOp_109_out;
	notOp #(.WIDTH(1)) notOp_109(.in(notOp_109_in0), .out(notOp_109_out));

	wire [0:0] andOp_110_in0;
	wire [0:0] andOp_110_in1;
	wire [0:0] andOp_110_out;
	andOp #(.WIDTH(1)) andOp_110(.in0(andOp_110_in0), .in1(andOp_110_in1), .out(andOp_110_out));

	wire [0:0] andOp_111_in0;
	wire [0:0] andOp_111_in1;
	wire [0:0] andOp_111_out;
	andOp #(.WIDTH(1)) andOp_111(.in0(andOp_111_in0), .in1(andOp_111_in1), .out(andOp_111_out));

	wire [0:0] notOp_112_in0;
	wire [0:0] notOp_112_out;
	notOp #(.WIDTH(1)) notOp_112(.in(notOp_112_in0), .out(notOp_112_out));

	wire [0:0] andOp_113_in0;
	wire [0:0] andOp_113_in1;
	wire [0:0] andOp_113_out;
	andOp #(.WIDTH(1)) andOp_113(.in0(andOp_113_in0), .in1(andOp_113_in1), .out(andOp_113_out));

	wire [0:0] notOp_114_in0;
	wire [0:0] notOp_114_out;
	notOp #(.WIDTH(1)) notOp_114(.in(notOp_114_in0), .out(notOp_114_out));

	wire [0:0] andOp_115_in0;
	wire [0:0] andOp_115_in1;
	wire [0:0] andOp_115_out;
	andOp #(.WIDTH(1)) andOp_115(.in0(andOp_115_in0), .in1(andOp_115_in1), .out(andOp_115_out));

	wire [31:0] eq_116_in0;
	wire [31:0] eq_116_in1;
	wire [0:0] eq_116_out;
	eq #(.WIDTH(32)) eq_116(.in0(eq_116_in0), .in1(eq_116_in1), .out(eq_116_out));

	wire [31:0] eq_117_in0;
	wire [31:0] eq_117_in1;
	wire [0:0] eq_117_out;
	eq #(.WIDTH(32)) eq_117(.in0(eq_117_in0), .in1(eq_117_in1), .out(eq_117_out));

	wire [31:0] eq_118_in0;
	wire [31:0] eq_118_in1;
	wire [0:0] eq_118_out;
	eq #(.WIDTH(32)) eq_118(.in0(eq_118_in0), .in1(eq_118_in1), .out(eq_118_out));

	wire [0:0] orOp_119_in0;
	wire [0:0] orOp_119_in1;
	wire [0:0] orOp_119_out;
	orOp #(.WIDTH(1)) orOp_119(.in0(orOp_119_in0), .in1(orOp_119_in1), .out(orOp_119_out));

	wire [31:0] eq_120_in0;
	wire [31:0] eq_120_in1;
	wire [0:0] eq_120_out;
	eq #(.WIDTH(32)) eq_120(.in0(eq_120_in0), .in1(eq_120_in1), .out(eq_120_out));

	wire [31:0] eq_121_in0;
	wire [31:0] eq_121_in1;
	wire [0:0] eq_121_out;
	eq #(.WIDTH(32)) eq_121(.in0(eq_121_in0), .in1(eq_121_in1), .out(eq_121_out));

	wire [31:0] eq_122_in0;
	wire [31:0] eq_122_in1;
	wire [0:0] eq_122_out;
	eq #(.WIDTH(32)) eq_122(.in0(eq_122_in0), .in1(eq_122_in1), .out(eq_122_out));

	wire [31:0] eq_123_in0;
	wire [31:0] eq_123_in1;
	wire [0:0] eq_123_out;
	eq #(.WIDTH(32)) eq_123(.in0(eq_123_in0), .in1(eq_123_in1), .out(eq_123_out));

	wire [31:0] eq_124_in0;
	wire [31:0] eq_124_in1;
	wire [0:0] eq_124_out;
	eq #(.WIDTH(32)) eq_124(.in0(eq_124_in0), .in1(eq_124_in1), .out(eq_124_out));

	wire [31:0] eq_125_in0;
	wire [31:0] eq_125_in1;
	wire [0:0] eq_125_out;
	eq #(.WIDTH(32)) eq_125(.in0(eq_125_in0), .in1(eq_125_in1), .out(eq_125_out));

	wire [0:0] orOp_126_in0;
	wire [0:0] orOp_126_in1;
	wire [0:0] orOp_126_out;
	orOp #(.WIDTH(1)) orOp_126(.in0(orOp_126_in0), .in1(orOp_126_in1), .out(orOp_126_out));

	wire [31:0] eq_127_in0;
	wire [31:0] eq_127_in1;
	wire [0:0] eq_127_out;
	eq #(.WIDTH(32)) eq_127(.in0(eq_127_in0), .in1(eq_127_in1), .out(eq_127_out));

	wire [31:0] eq_128_in0;
	wire [31:0] eq_128_in1;
	wire [0:0] eq_128_out;
	eq #(.WIDTH(32)) eq_128(.in0(eq_128_in0), .in1(eq_128_in1), .out(eq_128_out));

	wire [31:0] eq_129_in0;
	wire [31:0] eq_129_in1;
	wire [0:0] eq_129_out;
	eq #(.WIDTH(32)) eq_129(.in0(eq_129_in0), .in1(eq_129_in1), .out(eq_129_out));

	wire [31:0] eq_130_in0;
	wire [31:0] eq_130_in1;
	wire [0:0] eq_130_out;
	eq #(.WIDTH(32)) eq_130(.in0(eq_130_in0), .in1(eq_130_in1), .out(eq_130_out));

	wire [31:0] eq_131_in0;
	wire [31:0] eq_131_in1;
	wire [0:0] eq_131_out;
	eq #(.WIDTH(32)) eq_131(.in0(eq_131_in0), .in1(eq_131_in1), .out(eq_131_out));

	wire [0:0] notOp_132_in0;
	wire [0:0] notOp_132_out;
	notOp #(.WIDTH(1)) notOp_132(.in(notOp_132_in0), .out(notOp_132_out));

	wire [0:0] andOp_133_in0;
	wire [0:0] andOp_133_in1;
	wire [0:0] andOp_133_out;
	andOp #(.WIDTH(1)) andOp_133(.in0(andOp_133_in0), .in1(andOp_133_in1), .out(andOp_133_out));

	wire [31:0] eq_134_in0;
	wire [31:0] eq_134_in1;
	wire [0:0] eq_134_out;
	eq #(.WIDTH(32)) eq_134(.in0(eq_134_in0), .in1(eq_134_in1), .out(eq_134_out));

	wire [31:0] eq_135_in0;
	wire [31:0] eq_135_in1;
	wire [0:0] eq_135_out;
	eq #(.WIDTH(32)) eq_135(.in0(eq_135_in0), .in1(eq_135_in1), .out(eq_135_out));

	wire [31:0] eq_136_in0;
	wire [31:0] eq_136_in1;
	wire [0:0] eq_136_out;
	eq #(.WIDTH(32)) eq_136(.in0(eq_136_in0), .in1(eq_136_in1), .out(eq_136_out));

	wire [31:0] eq_137_in0;
	wire [31:0] eq_137_in1;
	wire [0:0] eq_137_out;
	eq #(.WIDTH(32)) eq_137(.in0(eq_137_in0), .in1(eq_137_in1), .out(eq_137_out));

	wire [31:0] eq_138_in0;
	wire [31:0] eq_138_in1;
	wire [0:0] eq_138_out;
	eq #(.WIDTH(32)) eq_138(.in0(eq_138_in0), .in1(eq_138_in1), .out(eq_138_out));

	wire [31:0] eq_139_in0;
	wire [31:0] eq_139_in1;
	wire [0:0] eq_139_out;
	eq #(.WIDTH(32)) eq_139(.in0(eq_139_in0), .in1(eq_139_in1), .out(eq_139_out));

	wire [0:0] notOp_140_in0;
	wire [0:0] notOp_140_out;
	notOp #(.WIDTH(1)) notOp_140(.in(notOp_140_in0), .out(notOp_140_out));

	wire [0:0] andOp_141_in0;
	wire [0:0] andOp_141_in1;
	wire [0:0] andOp_141_out;
	andOp #(.WIDTH(1)) andOp_141(.in0(andOp_141_in0), .in1(andOp_141_in1), .out(andOp_141_out));

	wire [31:0] eq_142_in0;
	wire [31:0] eq_142_in1;
	wire [0:0] eq_142_out;
	eq #(.WIDTH(32)) eq_142(.in0(eq_142_in0), .in1(eq_142_in1), .out(eq_142_out));

	wire [31:0] eq_143_in0;
	wire [31:0] eq_143_in1;
	wire [0:0] eq_143_out;
	eq #(.WIDTH(32)) eq_143(.in0(eq_143_in0), .in1(eq_143_in1), .out(eq_143_out));

	wire [0:0] andOp_144_in0;
	wire [0:0] andOp_144_in1;
	wire [0:0] andOp_144_out;
	andOp #(.WIDTH(1)) andOp_144(.in0(andOp_144_in0), .in1(andOp_144_in1), .out(andOp_144_out));

	wire [0:0] andOp_145_in0;
	wire [0:0] andOp_145_in1;
	wire [0:0] andOp_145_out;
	andOp #(.WIDTH(1)) andOp_145(.in0(andOp_145_in0), .in1(andOp_145_in1), .out(andOp_145_out));

	wire [31:0] concat_146_in0;
	wire [31:0] concat_146_in1;
	wire [63:0] concat_146_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_146(.in0(concat_146_in0), .in1(concat_146_in1), .out(concat_146_out));

	wire [31:0] concat_147_in0;
	wire [31:0] concat_147_in1;
	wire [63:0] concat_147_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_147(.in0(concat_147_in0), .in1(concat_147_in1), .out(concat_147_out));

	wire [0:0] andOp_148_in0;
	wire [0:0] andOp_148_in1;
	wire [0:0] andOp_148_out;
	andOp #(.WIDTH(1)) andOp_148(.in0(andOp_148_in0), .in1(andOp_148_in1), .out(andOp_148_out));

	wire [31:0] concat_149_in0;
	wire [31:0] concat_149_in1;
	wire [63:0] concat_149_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_149(.in0(concat_149_in0), .in1(concat_149_in1), .out(concat_149_out));

	wire [31:0] concat_150_in0;
	wire [31:0] concat_150_in1;
	wire [63:0] concat_150_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_150(.in0(concat_150_in0), .in1(concat_150_in1), .out(concat_150_out));

	wire [0:0] andOp_151_in0;
	wire [0:0] andOp_151_in1;
	wire [0:0] andOp_151_out;
	andOp #(.WIDTH(1)) andOp_151(.in0(andOp_151_in0), .in1(andOp_151_in1), .out(andOp_151_out));

	wire [0:0] andOp_152_in0;
	wire [0:0] andOp_152_in1;
	wire [0:0] andOp_152_out;
	andOp #(.WIDTH(1)) andOp_152(.in0(andOp_152_in0), .in1(andOp_152_in1), .out(andOp_152_out));

	wire [0:0] andOp_153_in0;
	wire [0:0] andOp_153_in1;
	wire [0:0] andOp_153_out;
	andOp #(.WIDTH(1)) andOp_153(.in0(andOp_153_in0), .in1(andOp_153_in1), .out(andOp_153_out));

	wire [0:0] andOp_154_in0;
	wire [0:0] andOp_154_in1;
	wire [0:0] andOp_154_out;
	andOp #(.WIDTH(1)) andOp_154(.in0(andOp_154_in0), .in1(andOp_154_in1), .out(andOp_154_out));

	wire [0:0] andOp_155_in0;
	wire [0:0] andOp_155_in1;
	wire [0:0] andOp_155_out;
	andOp #(.WIDTH(1)) andOp_155(.in0(andOp_155_in0), .in1(andOp_155_in1), .out(andOp_155_out));

	wire [0:0] andOp_156_in0;
	wire [0:0] andOp_156_in1;
	wire [0:0] andOp_156_out;
	andOp #(.WIDTH(1)) andOp_156(.in0(andOp_156_in0), .in1(andOp_156_in1), .out(andOp_156_out));

	wire [0:0] andOp_157_in0;
	wire [0:0] andOp_157_in1;
	wire [0:0] andOp_157_out;
	andOp #(.WIDTH(1)) andOp_157(.in0(andOp_157_in0), .in1(andOp_157_in1), .out(andOp_157_out));

	wire [0:0] andOp_158_in0;
	wire [0:0] andOp_158_in1;
	wire [0:0] andOp_158_out;
	andOp #(.WIDTH(1)) andOp_158(.in0(andOp_158_in0), .in1(andOp_158_in1), .out(andOp_158_out));

	wire [0:0] andOp_159_in0;
	wire [0:0] andOp_159_in1;
	wire [0:0] andOp_159_out;
	andOp #(.WIDTH(1)) andOp_159(.in0(andOp_159_in0), .in1(andOp_159_in1), .out(andOp_159_out));

	wire [0:0] andOp_160_in0;
	wire [0:0] andOp_160_in1;
	wire [0:0] andOp_160_out;
	andOp #(.WIDTH(1)) andOp_160(.in0(andOp_160_in0), .in1(andOp_160_in1), .out(andOp_160_out));

	wire [0:0] andOp_161_in0;
	wire [0:0] andOp_161_in1;
	wire [0:0] andOp_161_out;
	andOp #(.WIDTH(1)) andOp_161(.in0(andOp_161_in0), .in1(andOp_161_in1), .out(andOp_161_out));

	wire [0:0] andOp_162_in0;
	wire [0:0] andOp_162_in1;
	wire [0:0] andOp_162_out;
	andOp #(.WIDTH(1)) andOp_162(.in0(andOp_162_in0), .in1(andOp_162_in1), .out(andOp_162_out));

	wire [0:0] andOp_163_in0;
	wire [0:0] andOp_163_in1;
	wire [0:0] andOp_163_out;
	andOp #(.WIDTH(1)) andOp_163(.in0(andOp_163_in0), .in1(andOp_163_in1), .out(andOp_163_out));

	wire [0:0] andOp_164_in0;
	wire [0:0] andOp_164_in1;
	wire [0:0] andOp_164_out;
	andOp #(.WIDTH(1)) andOp_164(.in0(andOp_164_in0), .in1(andOp_164_in1), .out(andOp_164_out));

	wire [0:0] andOp_165_in0;
	wire [0:0] andOp_165_in1;
	wire [0:0] andOp_165_out;
	andOp #(.WIDTH(1)) andOp_165(.in0(andOp_165_in0), .in1(andOp_165_in1), .out(andOp_165_out));

	wire [0:0] andOp_166_in0;
	wire [0:0] andOp_166_in1;
	wire [0:0] andOp_166_out;
	andOp #(.WIDTH(1)) andOp_166(.in0(andOp_166_in0), .in1(andOp_166_in1), .out(andOp_166_out));

	wire [0:0] andOp_167_in0;
	wire [0:0] andOp_167_in1;
	wire [0:0] andOp_167_out;
	andOp #(.WIDTH(1)) andOp_167(.in0(andOp_167_in0), .in1(andOp_167_in1), .out(andOp_167_out));

	wire [0:0] andOp_168_in0;
	wire [0:0] andOp_168_in1;
	wire [0:0] andOp_168_out;
	andOp #(.WIDTH(1)) andOp_168(.in0(andOp_168_in0), .in1(andOp_168_in1), .out(andOp_168_out));

	wire [0:0] andOp_169_in0;
	wire [0:0] andOp_169_in1;
	wire [0:0] andOp_169_out;
	andOp #(.WIDTH(1)) andOp_169(.in0(andOp_169_in0), .in1(andOp_169_in1), .out(andOp_169_out));

	wire [0:0] andOp_170_in0;
	wire [0:0] andOp_170_in1;
	wire [0:0] andOp_170_out;
	andOp #(.WIDTH(1)) andOp_170(.in0(andOp_170_in0), .in1(andOp_170_in1), .out(andOp_170_out));

	wire [0:0] notOp_171_in0;
	wire [0:0] notOp_171_out;
	notOp #(.WIDTH(1)) notOp_171(.in(notOp_171_in0), .out(notOp_171_out));

	wire [0:0] andOp_172_in0;
	wire [0:0] andOp_172_in1;
	wire [0:0] andOp_172_out;
	andOp #(.WIDTH(1)) andOp_172(.in0(andOp_172_in0), .in1(andOp_172_in1), .out(andOp_172_out));

	wire [0:0] notOp_173_in0;
	wire [0:0] notOp_173_out;
	notOp #(.WIDTH(1)) notOp_173(.in(notOp_173_in0), .out(notOp_173_out));

	wire [0:0] andOp_174_in0;
	wire [0:0] andOp_174_in1;
	wire [0:0] andOp_174_out;
	andOp #(.WIDTH(1)) andOp_174(.in0(andOp_174_in0), .in1(andOp_174_in1), .out(andOp_174_out));

	wire [0:0] notOp_175_in0;
	wire [0:0] notOp_175_out;
	notOp #(.WIDTH(1)) notOp_175(.in(notOp_175_in0), .out(notOp_175_out));

	wire [0:0] andOp_176_in0;
	wire [0:0] andOp_176_in1;
	wire [0:0] andOp_176_out;
	andOp #(.WIDTH(1)) andOp_176(.in0(andOp_176_in0), .in1(andOp_176_in1), .out(andOp_176_out));

	wire [0:0] notOp_177_in0;
	wire [0:0] notOp_177_out;
	notOp #(.WIDTH(1)) notOp_177(.in(notOp_177_in0), .out(notOp_177_out));

	wire [0:0] andOp_178_in0;
	wire [0:0] andOp_178_in1;
	wire [0:0] andOp_178_out;
	andOp #(.WIDTH(1)) andOp_178(.in0(andOp_178_in0), .in1(andOp_178_in1), .out(andOp_178_out));

	wire [0:0] notOp_179_in0;
	wire [0:0] notOp_179_out;
	notOp #(.WIDTH(1)) notOp_179(.in(notOp_179_in0), .out(notOp_179_out));

	wire [0:0] andOp_180_in0;
	wire [0:0] andOp_180_in1;
	wire [0:0] andOp_180_out;
	andOp #(.WIDTH(1)) andOp_180(.in0(andOp_180_in0), .in1(andOp_180_in1), .out(andOp_180_out));

	wire [0:0] notOp_181_in0;
	wire [0:0] notOp_181_out;
	notOp #(.WIDTH(1)) notOp_181(.in(notOp_181_in0), .out(notOp_181_out));

	wire [0:0] andOp_182_in0;
	wire [0:0] andOp_182_in1;
	wire [0:0] andOp_182_out;
	andOp #(.WIDTH(1)) andOp_182(.in0(andOp_182_in0), .in1(andOp_182_in1), .out(andOp_182_out));

	wire [0:0] andOp_183_in0;
	wire [0:0] andOp_183_in1;
	wire [0:0] andOp_183_out;
	andOp #(.WIDTH(1)) andOp_183(.in0(andOp_183_in0), .in1(andOp_183_in1), .out(andOp_183_out));

	wire [0:0] andOp_184_in0;
	wire [0:0] andOp_184_in1;
	wire [0:0] andOp_184_out;
	andOp #(.WIDTH(1)) andOp_184(.in0(andOp_184_in0), .in1(andOp_184_in1), .out(andOp_184_out));

	wire [0:0] andOp_185_in0;
	wire [0:0] andOp_185_in1;
	wire [0:0] andOp_185_out;
	andOp #(.WIDTH(1)) andOp_185(.in0(andOp_185_in0), .in1(andOp_185_in1), .out(andOp_185_out));

	wire [0:0] notOp_186_in0;
	wire [0:0] notOp_186_out;
	notOp #(.WIDTH(1)) notOp_186(.in(notOp_186_in0), .out(notOp_186_out));

	wire [0:0] andOp_187_in0;
	wire [0:0] andOp_187_in1;
	wire [0:0] andOp_187_out;
	andOp #(.WIDTH(1)) andOp_187(.in0(andOp_187_in0), .in1(andOp_187_in1), .out(andOp_187_out));

	wire [0:0] notOp_188_in0;
	wire [0:0] notOp_188_out;
	notOp #(.WIDTH(1)) notOp_188(.in(notOp_188_in0), .out(notOp_188_out));

	wire [0:0] andOp_189_in0;
	wire [0:0] andOp_189_in1;
	wire [0:0] andOp_189_out;
	andOp #(.WIDTH(1)) andOp_189(.in0(andOp_189_in0), .in1(andOp_189_in1), .out(andOp_189_out));

	wire [0:0] notOp_190_in0;
	wire [0:0] notOp_190_out;
	notOp #(.WIDTH(1)) notOp_190(.in(notOp_190_in0), .out(notOp_190_out));

	wire [0:0] andOp_191_in0;
	wire [0:0] andOp_191_in1;
	wire [0:0] andOp_191_out;
	andOp #(.WIDTH(1)) andOp_191(.in0(andOp_191_in0), .in1(andOp_191_in1), .out(andOp_191_out));

	wire [0:0] notOp_192_in0;
	wire [0:0] notOp_192_out;
	notOp #(.WIDTH(1)) notOp_192(.in(notOp_192_in0), .out(notOp_192_out));

	wire [0:0] andOp_193_in0;
	wire [0:0] andOp_193_in1;
	wire [0:0] andOp_193_out;
	andOp #(.WIDTH(1)) andOp_193(.in0(andOp_193_in0), .in1(andOp_193_in1), .out(andOp_193_out));

	wire [0:0] notOp_194_in0;
	wire [0:0] notOp_194_out;
	notOp #(.WIDTH(1)) notOp_194(.in(notOp_194_in0), .out(notOp_194_out));

	wire [0:0] andOp_195_in0;
	wire [0:0] andOp_195_in1;
	wire [0:0] andOp_195_out;
	andOp #(.WIDTH(1)) andOp_195(.in0(andOp_195_in0), .in1(andOp_195_in1), .out(andOp_195_out));

	wire [0:0] notOp_196_in0;
	wire [0:0] notOp_196_out;
	notOp #(.WIDTH(1)) notOp_196(.in(notOp_196_in0), .out(notOp_196_out));

	wire [0:0] andOp_197_in0;
	wire [0:0] andOp_197_in1;
	wire [0:0] andOp_197_out;
	andOp #(.WIDTH(1)) andOp_197(.in0(andOp_197_in0), .in1(andOp_197_in1), .out(andOp_197_out));

	wire [0:0] andOp_198_in0;
	wire [0:0] andOp_198_in1;
	wire [0:0] andOp_198_out;
	andOp #(.WIDTH(1)) andOp_198(.in0(andOp_198_in0), .in1(andOp_198_in1), .out(andOp_198_out));

	wire [0:0] andOp_199_in0;
	wire [0:0] andOp_199_in1;
	wire [0:0] andOp_199_out;
	andOp #(.WIDTH(1)) andOp_199(.in0(andOp_199_in0), .in1(andOp_199_in1), .out(andOp_199_out));

	wire [0:0] andOp_200_in0;
	wire [0:0] andOp_200_in1;
	wire [0:0] andOp_200_out;
	andOp #(.WIDTH(1)) andOp_200(.in0(andOp_200_in0), .in1(andOp_200_in1), .out(andOp_200_out));

	wire [0:0] notOp_201_in0;
	wire [0:0] notOp_201_out;
	notOp #(.WIDTH(1)) notOp_201(.in(notOp_201_in0), .out(notOp_201_out));

	wire [0:0] andOp_202_in0;
	wire [0:0] andOp_202_in1;
	wire [0:0] andOp_202_out;
	andOp #(.WIDTH(1)) andOp_202(.in0(andOp_202_in0), .in1(andOp_202_in1), .out(andOp_202_out));

	wire [0:0] notOp_203_in0;
	wire [0:0] notOp_203_out;
	notOp #(.WIDTH(1)) notOp_203(.in(notOp_203_in0), .out(notOp_203_out));

	wire [0:0] andOp_204_in0;
	wire [0:0] andOp_204_in1;
	wire [0:0] andOp_204_out;
	andOp #(.WIDTH(1)) andOp_204(.in0(andOp_204_in0), .in1(andOp_204_in1), .out(andOp_204_out));

	wire [0:0] notOp_205_in0;
	wire [0:0] notOp_205_out;
	notOp #(.WIDTH(1)) notOp_205(.in(notOp_205_in0), .out(notOp_205_out));

	wire [0:0] andOp_206_in0;
	wire [0:0] andOp_206_in1;
	wire [0:0] andOp_206_out;
	andOp #(.WIDTH(1)) andOp_206(.in0(andOp_206_in0), .in1(andOp_206_in1), .out(andOp_206_out));

	wire [0:0] notOp_207_in0;
	wire [0:0] notOp_207_out;
	notOp #(.WIDTH(1)) notOp_207(.in(notOp_207_in0), .out(notOp_207_out));

	wire [0:0] andOp_208_in0;
	wire [0:0] andOp_208_in1;
	wire [0:0] andOp_208_out;
	andOp #(.WIDTH(1)) andOp_208(.in0(andOp_208_in0), .in1(andOp_208_in1), .out(andOp_208_out));

	wire [0:0] notOp_209_in0;
	wire [0:0] notOp_209_out;
	notOp #(.WIDTH(1)) notOp_209(.in(notOp_209_in0), .out(notOp_209_out));

	wire [0:0] andOp_210_in0;
	wire [0:0] andOp_210_in1;
	wire [0:0] andOp_210_out;
	andOp #(.WIDTH(1)) andOp_210(.in0(andOp_210_in0), .in1(andOp_210_in1), .out(andOp_210_out));

	wire [0:0] notOp_211_in0;
	wire [0:0] notOp_211_out;
	notOp #(.WIDTH(1)) notOp_211(.in(notOp_211_in0), .out(notOp_211_out));

	wire [0:0] andOp_212_in0;
	wire [0:0] andOp_212_in1;
	wire [0:0] andOp_212_out;
	andOp #(.WIDTH(1)) andOp_212(.in0(andOp_212_in0), .in1(andOp_212_in1), .out(andOp_212_out));

	wire [0:0] notOp_213_in0;
	wire [0:0] notOp_213_out;
	notOp #(.WIDTH(1)) notOp_213(.in(notOp_213_in0), .out(notOp_213_out));

	wire [0:0] andOp_214_in0;
	wire [0:0] andOp_214_in1;
	wire [0:0] andOp_214_out;
	andOp #(.WIDTH(1)) andOp_214(.in0(andOp_214_in0), .in1(andOp_214_in1), .out(andOp_214_out));

	wire [0:0] notOp_215_in0;
	wire [0:0] notOp_215_out;
	notOp #(.WIDTH(1)) notOp_215(.in(notOp_215_in0), .out(notOp_215_out));

	wire [0:0] andOp_216_in0;
	wire [0:0] andOp_216_in1;
	wire [0:0] andOp_216_out;
	andOp #(.WIDTH(1)) andOp_216(.in0(andOp_216_in0), .in1(andOp_216_in1), .out(andOp_216_out));

	wire [0:0] notOp_217_in0;
	wire [0:0] notOp_217_out;
	notOp #(.WIDTH(1)) notOp_217(.in(notOp_217_in0), .out(notOp_217_out));

	wire [0:0] andOp_218_in0;
	wire [0:0] andOp_218_in1;
	wire [0:0] andOp_218_out;
	andOp #(.WIDTH(1)) andOp_218(.in0(andOp_218_in0), .in1(andOp_218_in1), .out(andOp_218_out));

	wire [0:0] notOp_219_in0;
	wire [0:0] notOp_219_out;
	notOp #(.WIDTH(1)) notOp_219(.in(notOp_219_in0), .out(notOp_219_out));

	wire [0:0] andOp_220_in0;
	wire [0:0] andOp_220_in1;
	wire [0:0] andOp_220_out;
	andOp #(.WIDTH(1)) andOp_220(.in0(andOp_220_in0), .in1(andOp_220_in1), .out(andOp_220_out));

	wire [0:0] notOp_221_in0;
	wire [0:0] notOp_221_out;
	notOp #(.WIDTH(1)) notOp_221(.in(notOp_221_in0), .out(notOp_221_out));

	wire [0:0] andOp_222_in0;
	wire [0:0] andOp_222_in1;
	wire [0:0] andOp_222_out;
	andOp #(.WIDTH(1)) andOp_222(.in0(andOp_222_in0), .in1(andOp_222_in1), .out(andOp_222_out));

	wire [0:0] notOp_223_in0;
	wire [0:0] notOp_223_out;
	notOp #(.WIDTH(1)) notOp_223(.in(notOp_223_in0), .out(notOp_223_out));

	wire [0:0] andOp_224_in0;
	wire [0:0] andOp_224_in1;
	wire [0:0] andOp_224_out;
	andOp #(.WIDTH(1)) andOp_224(.in0(andOp_224_in0), .in1(andOp_224_in1), .out(andOp_224_out));

	reg [0:0] in_pipeline_0_in_data;
	wire [0:0] in_pipeline_0_out_data;
	hls_wire #(.WIDTH(1)) in_pipeline_0(.in_data(in_pipeline_0_in_data), .out_data(in_pipeline_0_out_data));

	wire [0:0] orOp_225_in0;
	wire [0:0] orOp_225_in1;
	wire [0:0] orOp_225_out;
	orOp #(.WIDTH(1)) orOp_225(.in0(orOp_225_in0), .in1(orOp_225_in1), .out(orOp_225_out));

	wire [0:0] orOp_226_in0;
	wire [0:0] orOp_226_in1;
	wire [0:0] orOp_226_out;
	orOp #(.WIDTH(1)) orOp_226(.in0(orOp_226_in0), .in1(orOp_226_in1), .out(orOp_226_out));

	wire [0:0] orOp_227_in0;
	wire [0:0] orOp_227_in1;
	wire [0:0] orOp_227_out;
	orOp #(.WIDTH(1)) orOp_227(.in0(orOp_227_in0), .in1(orOp_227_in1), .out(orOp_227_out));

	wire [0:0] orOp_228_in0;
	wire [0:0] orOp_228_in1;
	wire [0:0] orOp_228_out;
	orOp #(.WIDTH(1)) orOp_228(.in0(orOp_228_in0), .in1(orOp_228_in1), .out(orOp_228_out));

	wire [0:0] orOp_229_in0;
	wire [0:0] orOp_229_in1;
	wire [0:0] orOp_229_out;
	orOp #(.WIDTH(1)) orOp_229(.in0(orOp_229_in0), .in1(orOp_229_in1), .out(orOp_229_out));

	wire [0:0] orOp_230_in0;
	wire [0:0] orOp_230_in1;
	wire [0:0] orOp_230_out;
	orOp #(.WIDTH(1)) orOp_230(.in0(orOp_230_in0), .in1(orOp_230_in1), .out(orOp_230_out));

	wire [0:0] orOp_231_in0;
	wire [0:0] orOp_231_in1;
	wire [0:0] orOp_231_out;
	orOp #(.WIDTH(1)) orOp_231(.in0(orOp_231_in0), .in1(orOp_231_in1), .out(orOp_231_out));

	wire [31:0] eq_232_in0;
	wire [31:0] eq_232_in1;
	wire [0:0] eq_232_out;
	eq #(.WIDTH(32)) eq_232(.in0(eq_232_in0), .in1(eq_232_in1), .out(eq_232_out));

	wire [31:0] eq_233_in0;
	wire [31:0] eq_233_in1;
	wire [0:0] eq_233_out;
	eq #(.WIDTH(32)) eq_233(.in0(eq_233_in0), .in1(eq_233_in1), .out(eq_233_out));

	wire [31:0] eq_234_in0;
	wire [31:0] eq_234_in1;
	wire [0:0] eq_234_out;
	eq #(.WIDTH(32)) eq_234(.in0(eq_234_in0), .in1(eq_234_in1), .out(eq_234_out));

	wire [31:0] eq_235_in0;
	wire [31:0] eq_235_in1;
	wire [0:0] eq_235_out;
	eq #(.WIDTH(32)) eq_235(.in0(eq_235_in0), .in1(eq_235_in1), .out(eq_235_out));

	wire [0:0] andOp_236_in0;
	wire [0:0] andOp_236_in1;
	wire [0:0] andOp_236_out;
	andOp #(.WIDTH(1)) andOp_236(.in0(andOp_236_in0), .in1(andOp_236_in1), .out(andOp_236_out));

	wire [0:0] andOp_237_in0;
	wire [0:0] andOp_237_in1;
	wire [0:0] andOp_237_out;
	andOp #(.WIDTH(1)) andOp_237(.in0(andOp_237_in0), .in1(andOp_237_in1), .out(andOp_237_out));

	wire [0:0] andOp_238_in0;
	wire [0:0] andOp_238_in1;
	wire [0:0] andOp_238_out;
	andOp #(.WIDTH(1)) andOp_238(.in0(andOp_238_in0), .in1(andOp_238_in1), .out(andOp_238_out));

	wire [0:0] andOp_239_in0;
	wire [0:0] andOp_239_in1;
	wire [0:0] andOp_239_out;
	andOp #(.WIDTH(1)) andOp_239(.in0(andOp_239_in0), .in1(andOp_239_in1), .out(andOp_239_out));

	wire [31:0] eq_240_in0;
	wire [31:0] eq_240_in1;
	wire [0:0] eq_240_out;
	eq #(.WIDTH(32)) eq_240(.in0(eq_240_in0), .in1(eq_240_in1), .out(eq_240_out));

	wire [31:0] eq_241_in0;
	wire [31:0] eq_241_in1;
	wire [0:0] eq_241_out;
	eq #(.WIDTH(32)) eq_241(.in0(eq_241_in0), .in1(eq_241_in1), .out(eq_241_out));

	wire [0:0] andOp_242_in0;
	wire [0:0] andOp_242_in1;
	wire [0:0] andOp_242_out;
	andOp #(.WIDTH(1)) andOp_242(.in0(andOp_242_in0), .in1(andOp_242_in1), .out(andOp_242_out));

	wire [31:0] eq_243_in0;
	wire [31:0] eq_243_in1;
	wire [0:0] eq_243_out;
	eq #(.WIDTH(32)) eq_243(.in0(eq_243_in0), .in1(eq_243_in1), .out(eq_243_out));

	wire [31:0] eq_244_in0;
	wire [31:0] eq_244_in1;
	wire [0:0] eq_244_out;
	eq #(.WIDTH(32)) eq_244(.in0(eq_244_in0), .in1(eq_244_in1), .out(eq_244_out));

	wire [0:0] andOp_245_in0;
	wire [0:0] andOp_245_in1;
	wire [0:0] andOp_245_out;
	andOp #(.WIDTH(1)) andOp_245(.in0(andOp_245_in0), .in1(andOp_245_in1), .out(andOp_245_out));

	wire [31:0] eq_246_in0;
	wire [31:0] eq_246_in1;
	wire [0:0] eq_246_out;
	eq #(.WIDTH(32)) eq_246(.in0(eq_246_in0), .in1(eq_246_in1), .out(eq_246_out));

	wire [31:0] eq_247_in0;
	wire [31:0] eq_247_in1;
	wire [0:0] eq_247_out;
	eq #(.WIDTH(32)) eq_247(.in0(eq_247_in0), .in1(eq_247_in1), .out(eq_247_out));

	wire [31:0] eq_248_in0;
	wire [31:0] eq_248_in1;
	wire [0:0] eq_248_out;
	eq #(.WIDTH(32)) eq_248(.in0(eq_248_in0), .in1(eq_248_in1), .out(eq_248_out));

	wire [31:0] eq_249_in0;
	wire [31:0] eq_249_in1;
	wire [0:0] eq_249_out;
	eq #(.WIDTH(32)) eq_249(.in0(eq_249_in0), .in1(eq_249_in1), .out(eq_249_out));

	wire [31:0] eq_250_in0;
	wire [31:0] eq_250_in1;
	wire [0:0] eq_250_out;
	eq #(.WIDTH(32)) eq_250(.in0(eq_250_in0), .in1(eq_250_in1), .out(eq_250_out));

	wire [31:0] eq_251_in0;
	wire [31:0] eq_251_in1;
	wire [0:0] eq_251_out;
	eq #(.WIDTH(32)) eq_251(.in0(eq_251_in0), .in1(eq_251_in1), .out(eq_251_out));

	wire [31:0] eq_252_in0;
	wire [31:0] eq_252_in1;
	wire [0:0] eq_252_out;
	eq #(.WIDTH(32)) eq_252(.in0(eq_252_in0), .in1(eq_252_in1), .out(eq_252_out));

	wire [31:0] eq_253_in0;
	wire [31:0] eq_253_in1;
	wire [0:0] eq_253_out;
	eq #(.WIDTH(32)) eq_253(.in0(eq_253_in0), .in1(eq_253_in1), .out(eq_253_out));

	wire [31:0] eq_254_in0;
	wire [31:0] eq_254_in1;
	wire [0:0] eq_254_out;
	eq #(.WIDTH(32)) eq_254(.in0(eq_254_in0), .in1(eq_254_in1), .out(eq_254_out));

	wire [0:0] andOp_255_in0;
	wire [0:0] andOp_255_in1;
	wire [0:0] andOp_255_out;
	andOp #(.WIDTH(1)) andOp_255(.in0(andOp_255_in0), .in1(andOp_255_in1), .out(andOp_255_out));

	wire [31:0] eq_256_in0;
	wire [31:0] eq_256_in1;
	wire [0:0] eq_256_out;
	eq #(.WIDTH(32)) eq_256(.in0(eq_256_in0), .in1(eq_256_in1), .out(eq_256_out));

	wire [31:0] eq_257_in0;
	wire [31:0] eq_257_in1;
	wire [0:0] eq_257_out;
	eq #(.WIDTH(32)) eq_257(.in0(eq_257_in0), .in1(eq_257_in1), .out(eq_257_out));

	// End Functional Units

	reg [31:0] data_store_0_0;
	reg [31:0] data_store_0_2;
	reg [31:0] data_store_0_4;
	reg [31:0] data_store_0_6;
	reg [31:0] data_store_1_10;
	reg [31:0] data_store_1_12;
	reg [31:0] data_store_1_14;
	reg [31:0] data_store_1_15;
	reg [31:0] data_store_1_8;
	reg [31:0] data_store_2_17;
	reg [31:0] data_store_2_19;
	reg [31:0] data_store_2_21;
	reg [31:0] data_store_2_24;
	reg [31:0] data_store_2_25;
	reg [31:0] data_store_3_27;
	reg [31:0] data_store_3_29;
	reg [31:0] data_store_3_31;
	reg [31:0] data_store_3_33;
	reg [31:0] data_store_3_35;
	reg [31:0] data_store_3_37;
	reg [31:0] data_store_4_38;
	reg [31:0] data_store_4_40;
	reg [31:0] data_store_4_42;
	reg [31:0] data_store_4_45;
	reg [31:0] data_store_5_48;
	reg [31:0] data_store_5_50;
	reg [31:0] data_store_5_52;
	reg [31:0] data_store_5_54;
	reg [31:0] data_store_6_56;
	reg [31:0] data_store_6_58;
	reg [31:0] data_store_6_60;
	reg [31:0] data_store_6_62;
	reg [31:0] data_store_7_64;
	reg [31:0] data_store_7_66;
	reg [31:0] data_store_7_68;
	reg [31:0] data_store_7_70;
	reg [31:0] global_state;
	reg [0:0] out_of_pipe_7_8;
	reg [0:0] out_of_pipe_bb_7_8;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_3_last_state;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;
	reg [31:0] state_4_last_state;
	reg [31:0] state_5_entry_BB_reg;
	reg [0:0] state_5_is_active;
	reg [31:0] state_5_last_BB_reg;
	reg [31:0] state_5_last_state;
	reg [31:0] state_6_entry_BB_reg;
	reg [0:0] state_6_is_active;
	reg [31:0] state_6_last_BB_reg;
	reg [31:0] state_6_last_state;
	reg [31:0] state_7_entry_BB_reg;
	reg [0:0] state_7_is_active;
	reg [31:0] state_7_last_BB_reg;
	reg [31:0] state_7_last_state;
	reg [31:0] state_8_entry_BB_reg;
	reg [0:0] state_8_is_active;
	reg [31:0] state_8_last_BB_reg;
	reg [31:0] state_8_last_state;

	// controller for a.a_raddr_0_reg
	always @(*) begin
		if (andOp_154_out) begin 
			a_raddr_0_reg = add_add8_out;
		end else begin
			a_raddr_0_reg = 0;
		end
	end
	// controller for add_add12.add_add12_in0
	// controller for add_add12.add_add12_in1
	// Insensitive connections
	assign add_add12_in0 = b_rdata_0;
	assign add_add12_in1 = data_in_4_47_out_data;
	// controller for add_add17.add_add17_in0
	// controller for add_add17.add_add17_in1
	// Insensitive connections
	assign add_add17_in0 = data_in_7_69_out_data;
	assign add_add17_in1 = 32'd1;
	// controller for add_add6.add_add6_in0
	// controller for add_add6.add_add6_in1
	// Insensitive connections
	assign add_add6_in0 = phi_phi4_out;
	assign add_add6_in1 = 32'd1;
	// controller for add_add8.add_add8_in0
	// controller for add_add8.add_add8_in1
	// Insensitive connections
	assign add_add8_in0 = data_in_2_23_out_data;
	assign add_add8_in1 = data_in_2_20_out_data;
	// controller for andOp_100.andOp_100_in0
	// controller for andOp_100.andOp_100_in1
	// Insensitive connections
	assign andOp_100_in0 = andOp_96_out;
	assign andOp_100_in1 = notOp_99_out;
	// controller for andOp_101.andOp_101_in0
	// controller for andOp_101.andOp_101_in1
	// Insensitive connections
	assign andOp_101_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_101_in1 = state_1_is_active;
	// controller for andOp_103.andOp_103_in0
	// controller for andOp_103.andOp_103_in1
	// Insensitive connections
	assign andOp_103_in0 = andOp_101_out;
	assign andOp_103_in1 = icmp_icmp7_out;
	// controller for andOp_105.andOp_105_in0
	// controller for andOp_105.andOp_105_in1
	// Insensitive connections
	assign andOp_105_in0 = andOp_101_out;
	assign andOp_105_in1 = notOp_104_out;
	// controller for andOp_106.andOp_106_in0
	// controller for andOp_106.andOp_106_in1
	// Insensitive connections
	assign andOp_106_in0 = bb_3_active_in_state_7_out_data;
	assign andOp_106_in1 = state_7_is_active;
	// controller for andOp_108.andOp_108_in0
	// controller for andOp_108.andOp_108_in1
	// Insensitive connections
	assign andOp_108_in0 = andOp_106_out;
	assign andOp_108_in1 = icmp_icmp18_out;
	// controller for andOp_110.andOp_110_in0
	// controller for andOp_110.andOp_110_in1
	// Insensitive connections
	assign andOp_110_in0 = andOp_106_out;
	assign andOp_110_in1 = notOp_109_out;
	// controller for andOp_111.andOp_111_in0
	// controller for andOp_111.andOp_111_in1
	// Insensitive connections
	assign andOp_111_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_111_in1 = state_1_is_active;
	// controller for andOp_113.andOp_113_in0
	// controller for andOp_113.andOp_113_in1
	// Insensitive connections
	assign andOp_113_in0 = andOp_111_out;
	assign andOp_113_in1 = icmp_icmp7_out;
	// controller for andOp_115.andOp_115_in0
	// controller for andOp_115.andOp_115_in1
	// Insensitive connections
	assign andOp_115_in0 = andOp_111_out;
	assign andOp_115_in1 = notOp_114_out;
	// controller for andOp_133.andOp_133_in0
	// controller for andOp_133.andOp_133_in1
	// Insensitive connections
	assign andOp_133_in0 = notOp_132_out;
	assign andOp_133_in1 = andOp_74_out;
	// controller for andOp_141.andOp_141_in0
	// controller for andOp_141.andOp_141_in1
	// Insensitive connections
	assign andOp_141_in0 = notOp_140_out;
	assign andOp_141_in1 = andOp_78_out;
	// controller for andOp_144.andOp_144_in0
	// controller for andOp_144.andOp_144_in1
	// Insensitive connections
	assign andOp_144_in0 = bb_1_active_in_state_1_out_data;
	assign andOp_144_in1 = state_1_is_active;
	// controller for andOp_145.andOp_145_in0
	// controller for andOp_145.andOp_145_in1
	// Insensitive connections
	assign andOp_145_in0 = bb_1_active_in_state_1_out_data;
	assign andOp_145_in1 = state_1_is_active;
	// controller for andOp_148.andOp_148_in0
	// controller for andOp_148.andOp_148_in1
	// Insensitive connections
	assign andOp_148_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_148_in1 = state_1_is_active;
	// controller for andOp_151.andOp_151_in0
	// controller for andOp_151.andOp_151_in1
	// Insensitive connections
	assign andOp_151_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_151_in1 = state_1_is_active;
	// controller for andOp_152.andOp_152_in0
	// controller for andOp_152.andOp_152_in1
	// Insensitive connections
	assign andOp_152_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_152_in1 = state_1_is_active;
	// controller for andOp_153.andOp_153_in0
	// controller for andOp_153.andOp_153_in1
	// Insensitive connections
	assign andOp_153_in0 = bb_4_active_in_state_2_out_data;
	assign andOp_153_in1 = state_2_is_active;
	// controller for andOp_154.andOp_154_in0
	// controller for andOp_154.andOp_154_in1
	// Insensitive connections
	assign andOp_154_in0 = bb_4_active_in_state_2_out_data;
	assign andOp_154_in1 = state_2_is_active;
	// controller for andOp_155.andOp_155_in0
	// controller for andOp_155.andOp_155_in1
	// Insensitive connections
	assign andOp_155_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_155_in1 = state_3_is_active;
	// controller for andOp_156.andOp_156_in0
	// controller for andOp_156.andOp_156_in1
	// Insensitive connections
	assign andOp_156_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_156_in1 = state_3_is_active;
	// controller for andOp_157.andOp_157_in0
	// controller for andOp_157.andOp_157_in1
	// Insensitive connections
	assign andOp_157_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_157_in1 = state_4_is_active;
	// controller for andOp_158.andOp_158_in0
	// controller for andOp_158.andOp_158_in1
	// Insensitive connections
	assign andOp_158_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_158_in1 = state_4_is_active;
	// controller for andOp_159.andOp_159_in0
	// controller for andOp_159.andOp_159_in1
	// Insensitive connections
	assign andOp_159_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_159_in1 = state_4_is_active;
	// controller for andOp_160.andOp_160_in0
	// controller for andOp_160.andOp_160_in1
	// Insensitive connections
	assign andOp_160_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_160_in1 = state_4_is_active;
	// controller for andOp_161.andOp_161_in0
	// controller for andOp_161.andOp_161_in1
	// Insensitive connections
	assign andOp_161_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_161_in1 = state_4_is_active;
	// controller for andOp_162.andOp_162_in0
	// controller for andOp_162.andOp_162_in1
	// Insensitive connections
	assign andOp_162_in0 = bb_3_active_in_state_7_out_data;
	assign andOp_162_in1 = state_7_is_active;
	// controller for andOp_163.andOp_163_in0
	// controller for andOp_163.andOp_163_in1
	// Insensitive connections
	assign andOp_163_in0 = bb_3_active_in_state_7_out_data;
	assign andOp_163_in1 = state_7_is_active;
	// controller for andOp_164.andOp_164_in0
	// controller for andOp_164.andOp_164_in1
	// Insensitive connections
	assign andOp_164_in0 = bb_2_active_in_state_8_out_data;
	assign andOp_164_in1 = state_8_is_active;
	// controller for andOp_165.andOp_165_in0
	// controller for andOp_165.andOp_165_in1
	// Insensitive connections
	assign andOp_165_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_165_in1 = state_1_is_active;
	// controller for andOp_166.andOp_166_in0
	// controller for andOp_166.andOp_166_in1
	// Insensitive connections
	assign andOp_166_in0 = bb_4_active_in_state_2_out_data;
	assign andOp_166_in1 = state_2_is_active;
	// controller for andOp_167.andOp_167_in0
	// controller for andOp_167.andOp_167_in1
	// Insensitive connections
	assign andOp_167_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_167_in1 = state_3_is_active;
	// controller for andOp_168.andOp_168_in0
	// controller for andOp_168.andOp_168_in1
	// Insensitive connections
	assign andOp_168_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_168_in1 = state_4_is_active;
	// controller for andOp_169.andOp_169_in0
	// controller for andOp_169.andOp_169_in1
	// Insensitive connections
	assign andOp_169_in0 = bb_4_active_in_state_5_out_data;
	assign andOp_169_in1 = state_5_is_active;
	// controller for andOp_170.andOp_170_in0
	// controller for andOp_170.andOp_170_in1
	// Insensitive connections
	assign andOp_170_in0 = bb_4_active_in_state_6_out_data;
	assign andOp_170_in1 = state_6_is_active;
	// controller for andOp_172.andOp_172_in0
	// controller for andOp_172.andOp_172_in1
	// Insensitive connections
	assign andOp_172_in0 = 1'd1;
	assign andOp_172_in1 = notOp_171_out;
	// controller for andOp_174.andOp_174_in0
	// controller for andOp_174.andOp_174_in1
	// Insensitive connections
	assign andOp_174_in0 = andOp_172_out;
	assign andOp_174_in1 = notOp_173_out;
	// controller for andOp_176.andOp_176_in0
	// controller for andOp_176.andOp_176_in1
	// Insensitive connections
	assign andOp_176_in0 = andOp_174_out;
	assign andOp_176_in1 = notOp_175_out;
	// controller for andOp_178.andOp_178_in0
	// controller for andOp_178.andOp_178_in1
	// Insensitive connections
	assign andOp_178_in0 = andOp_176_out;
	assign andOp_178_in1 = notOp_177_out;
	// controller for andOp_180.andOp_180_in0
	// controller for andOp_180.andOp_180_in1
	// Insensitive connections
	assign andOp_180_in0 = andOp_178_out;
	assign andOp_180_in1 = notOp_179_out;
	// controller for andOp_182.andOp_182_in0
	// controller for andOp_182.andOp_182_in1
	// Insensitive connections
	assign andOp_182_in0 = andOp_180_out;
	assign andOp_182_in1 = notOp_181_out;
	// controller for andOp_183.andOp_183_in0
	// controller for andOp_183.andOp_183_in1
	// Insensitive connections
	assign andOp_183_in0 = in_pipeline_0_out_data;
	assign andOp_183_in1 = andOp_182_out;
	// controller for andOp_184.andOp_184_in0
	// controller for andOp_184.andOp_184_in1
	// Insensitive connections
	assign andOp_184_in0 = andOp_183_out;
	assign andOp_184_in1 = out_of_pipe_7_8;
	// controller for andOp_185.andOp_185_in0
	// controller for andOp_185.andOp_185_in1
	// Insensitive connections
	assign andOp_185_in0 = andOp_183_out;
	assign andOp_185_in1 = out_of_pipe_7_8;
	// controller for andOp_187.andOp_187_in0
	// controller for andOp_187.andOp_187_in1
	// Insensitive connections
	assign andOp_187_in0 = 1'd1;
	assign andOp_187_in1 = notOp_186_out;
	// controller for andOp_189.andOp_189_in0
	// controller for andOp_189.andOp_189_in1
	// Insensitive connections
	assign andOp_189_in0 = andOp_187_out;
	assign andOp_189_in1 = notOp_188_out;
	// controller for andOp_191.andOp_191_in0
	// controller for andOp_191.andOp_191_in1
	// Insensitive connections
	assign andOp_191_in0 = andOp_189_out;
	assign andOp_191_in1 = notOp_190_out;
	// controller for andOp_193.andOp_193_in0
	// controller for andOp_193.andOp_193_in1
	// Insensitive connections
	assign andOp_193_in0 = andOp_191_out;
	assign andOp_193_in1 = notOp_192_out;
	// controller for andOp_195.andOp_195_in0
	// controller for andOp_195.andOp_195_in1
	// Insensitive connections
	assign andOp_195_in0 = andOp_193_out;
	assign andOp_195_in1 = notOp_194_out;
	// controller for andOp_197.andOp_197_in0
	// controller for andOp_197.andOp_197_in1
	// Insensitive connections
	assign andOp_197_in0 = andOp_195_out;
	assign andOp_197_in1 = notOp_196_out;
	// controller for andOp_198.andOp_198_in0
	// controller for andOp_198.andOp_198_in1
	// Insensitive connections
	assign andOp_198_in0 = in_pipeline_0_out_data;
	assign andOp_198_in1 = andOp_197_out;
	// controller for andOp_199.andOp_199_in0
	// controller for andOp_199.andOp_199_in1
	// Insensitive connections
	assign andOp_199_in0 = andOp_198_out;
	assign andOp_199_in1 = out_of_pipe_bb_7_8;
	// controller for andOp_200.andOp_200_in0
	// controller for andOp_200.andOp_200_in1
	// Insensitive connections
	assign andOp_200_in0 = bb_2_active_in_state_8_out_data;
	assign andOp_200_in1 = state_8_is_active;
	// controller for andOp_202.andOp_202_in0
	// controller for andOp_202.andOp_202_in1
	// Insensitive connections
	assign andOp_202_in0 = notOp_201_out;
	assign andOp_202_in1 = 1'd1;
	// controller for andOp_204.andOp_204_in0
	// controller for andOp_204.andOp_204_in1
	// Insensitive connections
	assign andOp_204_in0 = notOp_203_out;
	assign andOp_204_in1 = andOp_202_out;
	// controller for andOp_206.andOp_206_in0
	// controller for andOp_206.andOp_206_in1
	// Insensitive connections
	assign andOp_206_in0 = notOp_205_out;
	assign andOp_206_in1 = andOp_204_out;
	// controller for andOp_208.andOp_208_in0
	// controller for andOp_208.andOp_208_in1
	// Insensitive connections
	assign andOp_208_in0 = notOp_207_out;
	assign andOp_208_in1 = 1'd1;
	// controller for andOp_210.andOp_210_in0
	// controller for andOp_210.andOp_210_in1
	// Insensitive connections
	assign andOp_210_in0 = notOp_209_out;
	assign andOp_210_in1 = 1'd1;
	// controller for andOp_212.andOp_212_in0
	// controller for andOp_212.andOp_212_in1
	// Insensitive connections
	assign andOp_212_in0 = notOp_211_out;
	assign andOp_212_in1 = 1'd1;
	// controller for andOp_214.andOp_214_in0
	// controller for andOp_214.andOp_214_in1
	// Insensitive connections
	assign andOp_214_in0 = notOp_213_out;
	assign andOp_214_in1 = 1'd1;
	// controller for andOp_216.andOp_216_in0
	// controller for andOp_216.andOp_216_in1
	// Insensitive connections
	assign andOp_216_in0 = notOp_215_out;
	assign andOp_216_in1 = 1'd1;
	// controller for andOp_218.andOp_218_in0
	// controller for andOp_218.andOp_218_in1
	// Insensitive connections
	assign andOp_218_in0 = notOp_217_out;
	assign andOp_218_in1 = 1'd1;
	// controller for andOp_220.andOp_220_in0
	// controller for andOp_220.andOp_220_in1
	// Insensitive connections
	assign andOp_220_in0 = notOp_219_out;
	assign andOp_220_in1 = andOp_218_out;
	// controller for andOp_222.andOp_222_in0
	// controller for andOp_222.andOp_222_in1
	// Insensitive connections
	assign andOp_222_in0 = notOp_221_out;
	assign andOp_222_in1 = 1'd1;
	// controller for andOp_224.andOp_224_in0
	// controller for andOp_224.andOp_224_in1
	// Insensitive connections
	assign andOp_224_in0 = notOp_223_out;
	assign andOp_224_in1 = andOp_222_out;
	// controller for andOp_236.andOp_236_in0
	// controller for andOp_236.andOp_236_in1
	// Insensitive connections
	assign andOp_236_in0 = bb_1_active_in_state_1_out_data;
	assign andOp_236_in1 = state_1_is_active;
	// controller for andOp_237.andOp_237_in0
	// controller for andOp_237.andOp_237_in1
	// Insensitive connections
	assign andOp_237_in0 = bb_1_active_in_state_1_out_data;
	assign andOp_237_in1 = state_1_is_active;
	// controller for andOp_238.andOp_238_in0
	// controller for andOp_238.andOp_238_in1
	// Insensitive connections
	assign andOp_238_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_238_in1 = state_1_is_active;
	// controller for andOp_239.andOp_239_in0
	// controller for andOp_239.andOp_239_in1
	// Insensitive connections
	assign andOp_239_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_239_in1 = state_1_is_active;
	// controller for andOp_242.andOp_242_in0
	// controller for andOp_242.andOp_242_in1
	// Insensitive connections
	assign andOp_242_in0 = bb_4_active_in_state_2_out_data;
	assign andOp_242_in1 = state_2_is_active;
	// controller for andOp_245.andOp_245_in0
	// controller for andOp_245.andOp_245_in1
	// Insensitive connections
	assign andOp_245_in0 = bb_4_active_in_state_3_out_data;
	assign andOp_245_in1 = state_3_is_active;
	// controller for andOp_255.andOp_255_in0
	// controller for andOp_255.andOp_255_in1
	// Insensitive connections
	assign andOp_255_in0 = bb_3_active_in_state_7_out_data;
	assign andOp_255_in1 = state_7_is_active;
	// controller for andOp_72.andOp_72_in0
	// controller for andOp_72.andOp_72_in1
	// Insensitive connections
	assign andOp_72_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_72_in1 = state_0_is_active;
	// controller for andOp_74.andOp_74_in0
	// controller for andOp_74.andOp_74_in1
	// Insensitive connections
	assign andOp_74_in0 = bb_1_active_in_state_1_out_data;
	assign andOp_74_in1 = state_1_is_active;
	// controller for andOp_76.andOp_76_in0
	// controller for andOp_76.andOp_76_in1
	// Insensitive connections
	assign andOp_76_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_76_in1 = state_1_is_active;
	// controller for andOp_78.andOp_78_in0
	// controller for andOp_78.andOp_78_in1
	// Insensitive connections
	assign andOp_78_in0 = andOp_76_out;
	assign andOp_78_in1 = icmp_icmp7_out;
	// controller for andOp_80.andOp_80_in0
	// controller for andOp_80.andOp_80_in1
	// Insensitive connections
	assign andOp_80_in0 = andOp_76_out;
	assign andOp_80_in1 = notOp_79_out;
	// controller for andOp_81.andOp_81_in0
	// controller for andOp_81.andOp_81_in1
	// Insensitive connections
	assign andOp_81_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_81_in1 = state_1_is_active;
	// controller for andOp_83.andOp_83_in0
	// controller for andOp_83.andOp_83_in1
	// Insensitive connections
	assign andOp_83_in0 = andOp_81_out;
	assign andOp_83_in1 = icmp_icmp7_out;
	// controller for andOp_85.andOp_85_in0
	// controller for andOp_85.andOp_85_in1
	// Insensitive connections
	assign andOp_85_in0 = andOp_81_out;
	assign andOp_85_in1 = notOp_84_out;
	// controller for andOp_86.andOp_86_in0
	// controller for andOp_86.andOp_86_in1
	// Insensitive connections
	assign andOp_86_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_86_in1 = state_1_is_active;
	// controller for andOp_88.andOp_88_in0
	// controller for andOp_88.andOp_88_in1
	// Insensitive connections
	assign andOp_88_in0 = andOp_86_out;
	assign andOp_88_in1 = icmp_icmp7_out;
	// controller for andOp_90.andOp_90_in0
	// controller for andOp_90.andOp_90_in1
	// Insensitive connections
	assign andOp_90_in0 = andOp_86_out;
	assign andOp_90_in1 = notOp_89_out;
	// controller for andOp_91.andOp_91_in0
	// controller for andOp_91.andOp_91_in1
	// Insensitive connections
	assign andOp_91_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_91_in1 = state_1_is_active;
	// controller for andOp_93.andOp_93_in0
	// controller for andOp_93.andOp_93_in1
	// Insensitive connections
	assign andOp_93_in0 = andOp_91_out;
	assign andOp_93_in1 = icmp_icmp7_out;
	// controller for andOp_95.andOp_95_in0
	// controller for andOp_95.andOp_95_in1
	// Insensitive connections
	assign andOp_95_in0 = andOp_91_out;
	assign andOp_95_in1 = notOp_94_out;
	// controller for andOp_96.andOp_96_in0
	// controller for andOp_96.andOp_96_in1
	// Insensitive connections
	assign andOp_96_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_96_in1 = state_1_is_active;
	// controller for andOp_98.andOp_98_in0
	// controller for andOp_98.andOp_98_in1
	// Insensitive connections
	assign andOp_98_in0 = andOp_96_out;
	assign andOp_98_in1 = icmp_icmp7_out;
	// controller for b.b_raddr_0_reg
	always @(*) begin
		if (andOp_156_out) begin 
			b_raddr_0_reg = data_in_3_34_out_data;
		end else begin
			b_raddr_0_reg = 0;
		end
	end
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_116_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_129_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_1.bb_1_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_1_in_data = eq_117_out;
		end else begin
			bb_1_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_1.bb_1_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_130_out) begin 
			bb_1_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_8.bb_2_active_in_state_8_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_8_in_data = eq_128_out;
		end else begin
			bb_2_active_in_state_8_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_8.bb_2_predecessor_in_state_8_in_data
	always @(*) begin
		if (eq_143_out) begin 
			bb_2_predecessor_in_state_8_in_data = state_8_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_8_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_7.bb_3_active_in_state_7_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_7_in_data = orOp_126_out;
		end else begin
			bb_3_active_in_state_7_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_7.bb_3_predecessor_in_state_7_in_data
	always @(*) begin
		if (andOp_141_out) begin 
			bb_3_predecessor_in_state_7_in_data = 32'd4;
		end else if (eq_139_out) begin 
			bb_3_predecessor_in_state_7_in_data = state_7_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_7_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_1.bb_4_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_1_in_data = orOp_119_out;
		end else begin
			bb_4_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_2.bb_4_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_2_in_data = eq_120_out;
		end else begin
			bb_4_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_3.bb_4_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_3_in_data = eq_121_out;
		end else begin
			bb_4_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_4.bb_4_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_4_in_data = eq_122_out;
		end else begin
			bb_4_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_5.bb_4_active_in_state_5_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_5_in_data = eq_123_out;
		end else begin
			bb_4_active_in_state_5_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_6.bb_4_active_in_state_6_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_6_in_data = eq_124_out;
		end else begin
			bb_4_active_in_state_6_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_7.bb_4_active_in_state_7_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_7_in_data = eq_127_out;
		end else begin
			bb_4_active_in_state_7_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_1.bb_4_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_133_out) begin 
			bb_4_predecessor_in_state_1_in_data = 32'd1;
		end else if (eq_131_out) begin 
			bb_4_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_2.bb_4_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_134_out) begin 
			bb_4_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_3.bb_4_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_135_out) begin 
			bb_4_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_4.bb_4_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_136_out) begin 
			bb_4_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_5.bb_4_predecessor_in_state_5_in_data
	always @(*) begin
		if (eq_137_out) begin 
			bb_4_predecessor_in_state_5_in_data = state_5_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_5_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_6.bb_4_predecessor_in_state_6_in_data
	always @(*) begin
		if (eq_138_out) begin 
			bb_4_predecessor_in_state_6_in_data = state_6_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_6_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_7.bb_4_predecessor_in_state_7_in_data
	always @(*) begin
		if (eq_142_out) begin 
			bb_4_predecessor_in_state_7_in_data = state_7_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_7_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_72_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_73_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_1_happened_in_state_1.br_1_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_74_out) begin 
			br_1_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_75_out) begin 
			br_1_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_1_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_7.br_3_happened_in_state_7_in_data
	always @(*) begin
		if (andOp_106_out) begin 
			br_3_happened_in_state_7_in_data = 1'd1;
		end else if (notOp_107_out) begin 
			br_3_happened_in_state_7_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_7_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_1.br_4_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_76_out) begin 
			br_4_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_77_out) begin 
			br_4_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_2.br_4_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_81_out) begin 
			br_4_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_82_out) begin 
			br_4_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_3.br_4_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_86_out) begin 
			br_4_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_87_out) begin 
			br_4_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_4.br_4_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_91_out) begin 
			br_4_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_92_out) begin 
			br_4_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_5.br_4_happened_in_state_5_in_data
	always @(*) begin
		if (andOp_96_out) begin 
			br_4_happened_in_state_5_in_data = 1'd1;
		end else if (notOp_97_out) begin 
			br_4_happened_in_state_5_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_5_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_6.br_4_happened_in_state_6_in_data
	always @(*) begin
		if (andOp_101_out) begin 
			br_4_happened_in_state_6_in_data = 1'd1;
		end else if (notOp_102_out) begin 
			br_4_happened_in_state_6_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_6_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_7.br_4_happened_in_state_7_in_data
	always @(*) begin
		if (andOp_111_out) begin 
			br_4_happened_in_state_7_in_data = 1'd1;
		end else if (notOp_112_out) begin 
			br_4_happened_in_state_7_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_7_in_data = 0;
		end
	end
	// controller for c.c_waddr_0_reg
	always @(*) begin
		if (andOp_160_out) begin 
			c_waddr_0_reg = data_in_4_44_out_data;
		end else begin
			c_waddr_0_reg = 0;
		end
	end
	// controller for c.c_wdata_0_reg
	always @(*) begin
		if (andOp_161_out) begin 
			c_wdata_0_reg = add_add12_out;
		end else begin
			c_wdata_0_reg = 0;
		end
	end
	// controller for c.c_wen_0_reg
	always @(*) begin
		if (andOp_159_out) begin 
			c_wen_0_reg = -(1'd1);
		end else begin
			c_wen_0_reg = 0;
		end
	end
	// controller for concat_146.concat_146_in0
	// controller for concat_146.concat_146_in1
	// Insensitive connections
	assign concat_146_in0 = data_in_1_9_out_data;
	assign concat_146_in1 = 32'd0;
	// controller for concat_147.concat_147_in0
	// controller for concat_147.concat_147_in1
	// Insensitive connections
	assign concat_147_in0 = 32'd3;
	assign concat_147_in1 = 32'd0;
	// controller for concat_149.concat_149_in0
	// controller for concat_149.concat_149_in1
	// Insensitive connections
	assign concat_149_in0 = data_in_1_16_out_data;
	assign concat_149_in1 = 32'd0;
	// controller for concat_150.concat_150_in0
	// controller for concat_150.concat_150_in1
	// Insensitive connections
	assign concat_150_in0 = 32'd4;
	assign concat_150_in1 = 32'd1;
	// controller for data_in_0_1.data_in_0_1_in_data
	always @(*) begin
		if (eq_232_out) begin 
			data_in_0_1_in_data = data_store_0_0;
		end else begin
			data_in_0_1_in_data = 0;
		end
	end
	// controller for data_in_0_3.data_in_0_3_in_data
	always @(*) begin
		if (eq_232_out) begin 
			data_in_0_3_in_data = data_store_0_2;
		end else begin
			data_in_0_3_in_data = 0;
		end
	end
	// controller for data_in_0_5.data_in_0_5_in_data
	always @(*) begin
		if (eq_232_out) begin 
			data_in_0_5_in_data = data_store_0_4;
		end else begin
			data_in_0_5_in_data = 0;
		end
	end
	// controller for data_in_0_7.data_in_0_7_in_data
	always @(*) begin
		if (eq_232_out) begin 
			data_in_0_7_in_data = data_store_0_6;
		end else begin
			data_in_0_7_in_data = 0;
		end
	end
	// controller for data_in_1_11.data_in_1_11_in_data
	always @(*) begin
		if (eq_233_out) begin 
			data_in_1_11_in_data = data_store_0_2;
		end else if (eq_234_out) begin 
			data_in_1_11_in_data = data_store_1_10;
		end else if (eq_235_out) begin 
			data_in_1_11_in_data = data_store_7_66;
		end else begin
			data_in_1_11_in_data = 0;
		end
	end
	// controller for data_in_1_13.data_in_1_13_in_data
	always @(*) begin
		if (eq_233_out) begin 
			data_in_1_13_in_data = data_store_0_4;
		end else if (eq_234_out) begin 
			data_in_1_13_in_data = data_store_1_12;
		end else if (eq_235_out) begin 
			data_in_1_13_in_data = data_store_7_68;
		end else begin
			data_in_1_13_in_data = 0;
		end
	end
	// controller for data_in_1_16.data_in_1_16_in_data
	always @(*) begin
		if (eq_233_out) begin 
			data_in_1_16_in_data = data_store_0_6;
		end else if (eq_234_out) begin 
			data_in_1_16_in_data = data_store_1_15;
		end else if (eq_235_out) begin 
			data_in_1_16_in_data = data_store_7_70;
		end else begin
			data_in_1_16_in_data = 0;
		end
	end
	// controller for data_in_1_9.data_in_1_9_in_data
	always @(*) begin
		if (eq_233_out) begin 
			data_in_1_9_in_data = data_store_0_0;
		end else if (eq_234_out) begin 
			data_in_1_9_in_data = data_store_1_8;
		end else if (eq_235_out) begin 
			data_in_1_9_in_data = data_store_7_64;
		end else begin
			data_in_1_9_in_data = 0;
		end
	end
	// controller for data_in_2_18.data_in_2_18_in_data
	always @(*) begin
		if (eq_240_out) begin 
			data_in_2_18_in_data = data_store_1_8;
		end else if (eq_241_out) begin 
			data_in_2_18_in_data = data_store_2_17;
		end else begin
			data_in_2_18_in_data = 0;
		end
	end
	// controller for data_in_2_20.data_in_2_20_in_data
	always @(*) begin
		if (eq_240_out) begin 
			data_in_2_20_in_data = data_store_1_10;
		end else if (eq_241_out) begin 
			data_in_2_20_in_data = data_store_2_19;
		end else begin
			data_in_2_20_in_data = 0;
		end
	end
	// controller for data_in_2_22.data_in_2_22_in_data
	always @(*) begin
		if (eq_240_out) begin 
			data_in_2_22_in_data = data_store_1_12;
		end else if (eq_241_out) begin 
			data_in_2_22_in_data = data_store_2_21;
		end else begin
			data_in_2_22_in_data = 0;
		end
	end
	// controller for data_in_2_23.data_in_2_23_in_data
	always @(*) begin
		if (eq_240_out) begin 
			data_in_2_23_in_data = data_store_1_14;
		end else if (eq_241_out) begin 
			data_in_2_23_in_data = 32'd0;
		end else begin
			data_in_2_23_in_data = 0;
		end
	end
	// controller for data_in_2_26.data_in_2_26_in_data
	always @(*) begin
		if (eq_240_out) begin 
			data_in_2_26_in_data = data_store_1_15;
		end else if (eq_241_out) begin 
			data_in_2_26_in_data = data_store_2_25;
		end else begin
			data_in_2_26_in_data = 0;
		end
	end
	// controller for data_in_3_28.data_in_3_28_in_data
	always @(*) begin
		if (eq_243_out) begin 
			data_in_3_28_in_data = data_store_2_17;
		end else if (eq_244_out) begin 
			data_in_3_28_in_data = data_store_3_27;
		end else begin
			data_in_3_28_in_data = 0;
		end
	end
	// controller for data_in_3_30.data_in_3_30_in_data
	always @(*) begin
		if (eq_243_out) begin 
			data_in_3_30_in_data = data_store_2_19;
		end else if (eq_244_out) begin 
			data_in_3_30_in_data = data_store_3_29;
		end else begin
			data_in_3_30_in_data = 0;
		end
	end
	// controller for data_in_3_32.data_in_3_32_in_data
	always @(*) begin
		if (eq_243_out) begin 
			data_in_3_32_in_data = data_store_2_21;
		end else if (eq_244_out) begin 
			data_in_3_32_in_data = data_store_3_31;
		end else begin
			data_in_3_32_in_data = 0;
		end
	end
	// controller for data_in_3_34.data_in_3_34_in_data
	always @(*) begin
		if (eq_243_out) begin 
			data_in_3_34_in_data = data_store_2_24;
		end else if (eq_244_out) begin 
			data_in_3_34_in_data = data_store_3_33;
		end else begin
			data_in_3_34_in_data = 0;
		end
	end
	// controller for data_in_3_36.data_in_3_36_in_data
	always @(*) begin
		if (eq_243_out) begin 
			data_in_3_36_in_data = data_store_2_25;
		end else if (eq_244_out) begin 
			data_in_3_36_in_data = data_store_3_35;
		end else begin
			data_in_3_36_in_data = 0;
		end
	end
	// controller for data_in_4_39.data_in_4_39_in_data
	always @(*) begin
		if (eq_246_out) begin 
			data_in_4_39_in_data = data_store_3_27;
		end else if (eq_247_out) begin 
			data_in_4_39_in_data = data_store_4_38;
		end else begin
			data_in_4_39_in_data = 0;
		end
	end
	// controller for data_in_4_41.data_in_4_41_in_data
	always @(*) begin
		if (eq_246_out) begin 
			data_in_4_41_in_data = data_store_3_29;
		end else if (eq_247_out) begin 
			data_in_4_41_in_data = data_store_4_40;
		end else begin
			data_in_4_41_in_data = 0;
		end
	end
	// controller for data_in_4_43.data_in_4_43_in_data
	always @(*) begin
		if (eq_246_out) begin 
			data_in_4_43_in_data = data_store_3_31;
		end else if (eq_247_out) begin 
			data_in_4_43_in_data = data_store_4_42;
		end else begin
			data_in_4_43_in_data = 0;
		end
	end
	// controller for data_in_4_44.data_in_4_44_in_data
	always @(*) begin
		if (eq_246_out) begin 
			data_in_4_44_in_data = data_store_3_33;
		end else if (eq_247_out) begin 
			data_in_4_44_in_data = 32'd0;
		end else begin
			data_in_4_44_in_data = 0;
		end
	end
	// controller for data_in_4_46.data_in_4_46_in_data
	always @(*) begin
		if (eq_246_out) begin 
			data_in_4_46_in_data = data_store_3_35;
		end else if (eq_247_out) begin 
			data_in_4_46_in_data = data_store_4_45;
		end else begin
			data_in_4_46_in_data = 0;
		end
	end
	// controller for data_in_4_47.data_in_4_47_in_data
	always @(*) begin
		if (eq_246_out) begin 
			data_in_4_47_in_data = data_store_3_37;
		end else if (eq_247_out) begin 
			data_in_4_47_in_data = 32'd0;
		end else begin
			data_in_4_47_in_data = 0;
		end
	end
	// controller for data_in_5_49.data_in_5_49_in_data
	always @(*) begin
		if (eq_248_out) begin 
			data_in_5_49_in_data = data_store_4_38;
		end else if (eq_249_out) begin 
			data_in_5_49_in_data = data_store_5_48;
		end else begin
			data_in_5_49_in_data = 0;
		end
	end
	// controller for data_in_5_51.data_in_5_51_in_data
	always @(*) begin
		if (eq_248_out) begin 
			data_in_5_51_in_data = data_store_4_40;
		end else if (eq_249_out) begin 
			data_in_5_51_in_data = data_store_5_50;
		end else begin
			data_in_5_51_in_data = 0;
		end
	end
	// controller for data_in_5_53.data_in_5_53_in_data
	always @(*) begin
		if (eq_248_out) begin 
			data_in_5_53_in_data = data_store_4_42;
		end else if (eq_249_out) begin 
			data_in_5_53_in_data = data_store_5_52;
		end else begin
			data_in_5_53_in_data = 0;
		end
	end
	// controller for data_in_5_55.data_in_5_55_in_data
	always @(*) begin
		if (eq_248_out) begin 
			data_in_5_55_in_data = data_store_4_45;
		end else if (eq_249_out) begin 
			data_in_5_55_in_data = data_store_5_54;
		end else begin
			data_in_5_55_in_data = 0;
		end
	end
	// controller for data_in_6_57.data_in_6_57_in_data
	always @(*) begin
		if (eq_250_out) begin 
			data_in_6_57_in_data = data_store_5_48;
		end else if (eq_251_out) begin 
			data_in_6_57_in_data = data_store_6_56;
		end else begin
			data_in_6_57_in_data = 0;
		end
	end
	// controller for data_in_6_59.data_in_6_59_in_data
	always @(*) begin
		if (eq_250_out) begin 
			data_in_6_59_in_data = data_store_5_50;
		end else if (eq_251_out) begin 
			data_in_6_59_in_data = data_store_6_58;
		end else begin
			data_in_6_59_in_data = 0;
		end
	end
	// controller for data_in_6_61.data_in_6_61_in_data
	always @(*) begin
		if (eq_250_out) begin 
			data_in_6_61_in_data = data_store_5_52;
		end else if (eq_251_out) begin 
			data_in_6_61_in_data = data_store_6_60;
		end else begin
			data_in_6_61_in_data = 0;
		end
	end
	// controller for data_in_6_63.data_in_6_63_in_data
	always @(*) begin
		if (eq_250_out) begin 
			data_in_6_63_in_data = data_store_5_54;
		end else if (eq_251_out) begin 
			data_in_6_63_in_data = data_store_6_62;
		end else begin
			data_in_6_63_in_data = 0;
		end
	end
	// controller for data_in_7_65.data_in_7_65_in_data
	always @(*) begin
		if (eq_252_out) begin 
			data_in_7_65_in_data = data_store_1_8;
		end else if (eq_253_out) begin 
			data_in_7_65_in_data = data_store_6_56;
		end else if (eq_254_out) begin 
			data_in_7_65_in_data = data_store_7_64;
		end else begin
			data_in_7_65_in_data = 0;
		end
	end
	// controller for data_in_7_67.data_in_7_67_in_data
	always @(*) begin
		if (eq_252_out) begin 
			data_in_7_67_in_data = data_store_1_10;
		end else if (eq_253_out) begin 
			data_in_7_67_in_data = data_store_6_58;
		end else if (eq_254_out) begin 
			data_in_7_67_in_data = data_store_7_66;
		end else begin
			data_in_7_67_in_data = 0;
		end
	end
	// controller for data_in_7_69.data_in_7_69_in_data
	always @(*) begin
		if (eq_252_out) begin 
			data_in_7_69_in_data = data_store_1_12;
		end else if (eq_253_out) begin 
			data_in_7_69_in_data = data_store_6_60;
		end else if (eq_254_out) begin 
			data_in_7_69_in_data = data_store_7_68;
		end else begin
			data_in_7_69_in_data = 0;
		end
	end
	// controller for data_in_7_71.data_in_7_71_in_data
	always @(*) begin
		if (eq_252_out) begin 
			data_in_7_71_in_data = data_store_1_15;
		end else if (eq_253_out) begin 
			data_in_7_71_in_data = data_store_6_62;
		end else if (eq_254_out) begin 
			data_in_7_71_in_data = data_store_7_70;
		end else begin
			data_in_7_71_in_data = 0;
		end
	end
	// controller for eq_116.eq_116_in0
	// controller for eq_116.eq_116_in1
	// Insensitive connections
	assign eq_116_in0 = 32'd0;
	assign eq_116_in1 = state_0_entry_BB_reg;
	// controller for eq_117.eq_117_in0
	// controller for eq_117.eq_117_in1
	// Insensitive connections
	assign eq_117_in0 = 32'd1;
	assign eq_117_in1 = state_1_entry_BB_reg;
	// controller for eq_118.eq_118_in0
	// controller for eq_118.eq_118_in1
	// Insensitive connections
	assign eq_118_in0 = 32'd4;
	assign eq_118_in1 = state_1_entry_BB_reg;
	// controller for eq_120.eq_120_in0
	// controller for eq_120.eq_120_in1
	// Insensitive connections
	assign eq_120_in0 = 32'd4;
	assign eq_120_in1 = state_2_entry_BB_reg;
	// controller for eq_121.eq_121_in0
	// controller for eq_121.eq_121_in1
	// Insensitive connections
	assign eq_121_in0 = 32'd4;
	assign eq_121_in1 = state_3_entry_BB_reg;
	// controller for eq_122.eq_122_in0
	// controller for eq_122.eq_122_in1
	// Insensitive connections
	assign eq_122_in0 = 32'd4;
	assign eq_122_in1 = state_4_entry_BB_reg;
	// controller for eq_123.eq_123_in0
	// controller for eq_123.eq_123_in1
	// Insensitive connections
	assign eq_123_in0 = 32'd4;
	assign eq_123_in1 = state_5_entry_BB_reg;
	// controller for eq_124.eq_124_in0
	// controller for eq_124.eq_124_in1
	// Insensitive connections
	assign eq_124_in0 = 32'd4;
	assign eq_124_in1 = state_6_entry_BB_reg;
	// controller for eq_125.eq_125_in0
	// controller for eq_125.eq_125_in1
	// Insensitive connections
	assign eq_125_in0 = 32'd3;
	assign eq_125_in1 = state_7_entry_BB_reg;
	// controller for eq_127.eq_127_in0
	// controller for eq_127.eq_127_in1
	// Insensitive connections
	assign eq_127_in0 = 32'd4;
	assign eq_127_in1 = state_7_entry_BB_reg;
	// controller for eq_128.eq_128_in0
	// controller for eq_128.eq_128_in1
	// Insensitive connections
	assign eq_128_in0 = 32'd2;
	assign eq_128_in1 = state_8_entry_BB_reg;
	// controller for eq_129.eq_129_in0
	// controller for eq_129.eq_129_in1
	// Insensitive connections
	assign eq_129_in0 = 32'd0;
	assign eq_129_in1 = state_0_entry_BB_reg;
	// controller for eq_130.eq_130_in0
	// controller for eq_130.eq_130_in1
	// Insensitive connections
	assign eq_130_in0 = 32'd1;
	assign eq_130_in1 = state_1_entry_BB_reg;
	// controller for eq_131.eq_131_in0
	// controller for eq_131.eq_131_in1
	// Insensitive connections
	assign eq_131_in0 = 32'd4;
	assign eq_131_in1 = state_1_entry_BB_reg;
	// controller for eq_134.eq_134_in0
	// controller for eq_134.eq_134_in1
	// Insensitive connections
	assign eq_134_in0 = 32'd4;
	assign eq_134_in1 = state_2_entry_BB_reg;
	// controller for eq_135.eq_135_in0
	// controller for eq_135.eq_135_in1
	// Insensitive connections
	assign eq_135_in0 = 32'd4;
	assign eq_135_in1 = state_3_entry_BB_reg;
	// controller for eq_136.eq_136_in0
	// controller for eq_136.eq_136_in1
	// Insensitive connections
	assign eq_136_in0 = 32'd4;
	assign eq_136_in1 = state_4_entry_BB_reg;
	// controller for eq_137.eq_137_in0
	// controller for eq_137.eq_137_in1
	// Insensitive connections
	assign eq_137_in0 = 32'd4;
	assign eq_137_in1 = state_5_entry_BB_reg;
	// controller for eq_138.eq_138_in0
	// controller for eq_138.eq_138_in1
	// Insensitive connections
	assign eq_138_in0 = 32'd4;
	assign eq_138_in1 = state_6_entry_BB_reg;
	// controller for eq_139.eq_139_in0
	// controller for eq_139.eq_139_in1
	// Insensitive connections
	assign eq_139_in0 = 32'd3;
	assign eq_139_in1 = state_7_entry_BB_reg;
	// controller for eq_142.eq_142_in0
	// controller for eq_142.eq_142_in1
	// Insensitive connections
	assign eq_142_in0 = 32'd4;
	assign eq_142_in1 = state_7_entry_BB_reg;
	// controller for eq_143.eq_143_in0
	// controller for eq_143.eq_143_in1
	// Insensitive connections
	assign eq_143_in0 = 32'd2;
	assign eq_143_in1 = state_8_entry_BB_reg;
	// controller for eq_232.eq_232_in0
	// controller for eq_232.eq_232_in1
	// Insensitive connections
	assign eq_232_in0 = 32'd0;
	assign eq_232_in1 = state_0_last_state;
	// controller for eq_233.eq_233_in0
	// controller for eq_233.eq_233_in1
	// Insensitive connections
	assign eq_233_in0 = 32'd0;
	assign eq_233_in1 = state_1_last_state;
	// controller for eq_234.eq_234_in0
	// controller for eq_234.eq_234_in1
	// Insensitive connections
	assign eq_234_in0 = 32'd1;
	assign eq_234_in1 = state_1_last_state;
	// controller for eq_235.eq_235_in0
	// controller for eq_235.eq_235_in1
	// Insensitive connections
	assign eq_235_in0 = 32'd7;
	assign eq_235_in1 = state_1_last_state;
	// controller for eq_240.eq_240_in0
	// controller for eq_240.eq_240_in1
	// Insensitive connections
	assign eq_240_in0 = 32'd1;
	assign eq_240_in1 = state_2_last_state;
	// controller for eq_241.eq_241_in0
	// controller for eq_241.eq_241_in1
	// Insensitive connections
	assign eq_241_in0 = 32'd2;
	assign eq_241_in1 = state_2_last_state;
	// controller for eq_243.eq_243_in0
	// controller for eq_243.eq_243_in1
	// Insensitive connections
	assign eq_243_in0 = 32'd2;
	assign eq_243_in1 = state_3_last_state;
	// controller for eq_244.eq_244_in0
	// controller for eq_244.eq_244_in1
	// Insensitive connections
	assign eq_244_in0 = 32'd3;
	assign eq_244_in1 = state_3_last_state;
	// controller for eq_246.eq_246_in0
	// controller for eq_246.eq_246_in1
	// Insensitive connections
	assign eq_246_in0 = 32'd3;
	assign eq_246_in1 = state_4_last_state;
	// controller for eq_247.eq_247_in0
	// controller for eq_247.eq_247_in1
	// Insensitive connections
	assign eq_247_in0 = 32'd4;
	assign eq_247_in1 = state_4_last_state;
	// controller for eq_248.eq_248_in0
	// controller for eq_248.eq_248_in1
	// Insensitive connections
	assign eq_248_in0 = 32'd4;
	assign eq_248_in1 = state_5_last_state;
	// controller for eq_249.eq_249_in0
	// controller for eq_249.eq_249_in1
	// Insensitive connections
	assign eq_249_in0 = 32'd5;
	assign eq_249_in1 = state_5_last_state;
	// controller for eq_250.eq_250_in0
	// controller for eq_250.eq_250_in1
	// Insensitive connections
	assign eq_250_in0 = 32'd5;
	assign eq_250_in1 = state_6_last_state;
	// controller for eq_251.eq_251_in0
	// controller for eq_251.eq_251_in1
	// Insensitive connections
	assign eq_251_in0 = 32'd6;
	assign eq_251_in1 = state_6_last_state;
	// controller for eq_252.eq_252_in0
	// controller for eq_252.eq_252_in1
	// Insensitive connections
	assign eq_252_in0 = 32'd1;
	assign eq_252_in1 = state_7_last_state;
	// controller for eq_253.eq_253_in0
	// controller for eq_253.eq_253_in1
	// Insensitive connections
	assign eq_253_in0 = 32'd6;
	assign eq_253_in1 = state_7_last_state;
	// controller for eq_254.eq_254_in0
	// controller for eq_254.eq_254_in1
	// Insensitive connections
	assign eq_254_in0 = 32'd7;
	assign eq_254_in1 = state_7_last_state;
	// controller for eq_256.eq_256_in0
	// controller for eq_256.eq_256_in1
	// Insensitive connections
	assign eq_256_in0 = 32'd7;
	assign eq_256_in1 = state_8_last_state;
	// controller for eq_257.eq_257_in0
	// controller for eq_257.eq_257_in1
	// Insensitive connections
	assign eq_257_in0 = 32'd8;
	assign eq_257_in1 = state_8_last_state;
	// controller for icmp_icmp18.icmp_icmp18_in0
	// controller for icmp_icmp18.icmp_icmp18_in1
	// Insensitive connections
	assign icmp_icmp18_in0 = add_add17_out;
	assign icmp_icmp18_in1 = 32'd16;
	// controller for icmp_icmp7.icmp_icmp7_in0
	// controller for icmp_icmp7.icmp_icmp7_in1
	// Insensitive connections
	assign icmp_icmp7_in0 = add_add6_out;
	assign icmp_icmp7_in1 = 32'd16;
	// controller for in_pipeline_0.in_pipeline_0_in_data
	always @(*) begin
		if (1'd1) begin 
			in_pipeline_0_in_data = orOp_231_out;
		end else begin
			in_pipeline_0_in_data = 0;
		end
	end
	// controller for notOp_102.notOp_102_in0
	// Insensitive connections
	assign notOp_102_in0 = andOp_101_out;
	// controller for notOp_104.notOp_104_in0
	// Insensitive connections
	assign notOp_104_in0 = icmp_icmp7_out;
	// controller for notOp_107.notOp_107_in0
	// Insensitive connections
	assign notOp_107_in0 = andOp_106_out;
	// controller for notOp_109.notOp_109_in0
	// Insensitive connections
	assign notOp_109_in0 = icmp_icmp18_out;
	// controller for notOp_112.notOp_112_in0
	// Insensitive connections
	assign notOp_112_in0 = andOp_111_out;
	// controller for notOp_114.notOp_114_in0
	// Insensitive connections
	assign notOp_114_in0 = icmp_icmp7_out;
	// controller for notOp_132.notOp_132_in0
	// Insensitive connections
	assign notOp_132_in0 = eq_131_out;
	// controller for notOp_140.notOp_140_in0
	// Insensitive connections
	assign notOp_140_in0 = eq_139_out;
	// controller for notOp_171.notOp_171_in0
	// Insensitive connections
	assign notOp_171_in0 = state_1_is_active;
	// controller for notOp_173.notOp_173_in0
	// Insensitive connections
	assign notOp_173_in0 = state_2_is_active;
	// controller for notOp_175.notOp_175_in0
	// Insensitive connections
	assign notOp_175_in0 = state_3_is_active;
	// controller for notOp_177.notOp_177_in0
	// Insensitive connections
	assign notOp_177_in0 = state_4_is_active;
	// controller for notOp_179.notOp_179_in0
	// Insensitive connections
	assign notOp_179_in0 = state_5_is_active;
	// controller for notOp_181.notOp_181_in0
	// Insensitive connections
	assign notOp_181_in0 = state_6_is_active;
	// controller for notOp_186.notOp_186_in0
	// Insensitive connections
	assign notOp_186_in0 = state_1_is_active;
	// controller for notOp_188.notOp_188_in0
	// Insensitive connections
	assign notOp_188_in0 = state_2_is_active;
	// controller for notOp_190.notOp_190_in0
	// Insensitive connections
	assign notOp_190_in0 = state_3_is_active;
	// controller for notOp_192.notOp_192_in0
	// Insensitive connections
	assign notOp_192_in0 = state_4_is_active;
	// controller for notOp_194.notOp_194_in0
	// Insensitive connections
	assign notOp_194_in0 = state_5_is_active;
	// controller for notOp_196.notOp_196_in0
	// Insensitive connections
	assign notOp_196_in0 = state_6_is_active;
	// controller for notOp_201.notOp_201_in0
	// Insensitive connections
	assign notOp_201_in0 = andOp_110_out;
	// controller for notOp_203.notOp_203_in0
	// Insensitive connections
	assign notOp_203_in0 = andOp_72_out;
	// controller for notOp_205.notOp_205_in0
	// Insensitive connections
	assign notOp_205_in0 = andOp_80_out;
	// controller for notOp_207.notOp_207_in0
	// Insensitive connections
	assign notOp_207_in0 = andOp_165_out;
	// controller for notOp_209.notOp_209_in0
	// Insensitive connections
	assign notOp_209_in0 = andOp_166_out;
	// controller for notOp_211.notOp_211_in0
	// Insensitive connections
	assign notOp_211_in0 = andOp_167_out;
	// controller for notOp_213.notOp_213_in0
	// Insensitive connections
	assign notOp_213_in0 = andOp_168_out;
	// controller for notOp_215.notOp_215_in0
	// Insensitive connections
	assign notOp_215_in0 = andOp_169_out;
	// controller for notOp_217.notOp_217_in0
	// Insensitive connections
	assign notOp_217_in0 = andOp_170_out;
	// controller for notOp_219.notOp_219_in0
	// Insensitive connections
	assign notOp_219_in0 = andOp_78_out;
	// controller for notOp_221.notOp_221_in0
	// Insensitive connections
	assign notOp_221_in0 = andOp_185_out;
	// controller for notOp_223.notOp_223_in0
	// Insensitive connections
	assign notOp_223_in0 = andOp_200_out;
	// controller for notOp_73.notOp_73_in0
	// Insensitive connections
	assign notOp_73_in0 = andOp_72_out;
	// controller for notOp_75.notOp_75_in0
	// Insensitive connections
	assign notOp_75_in0 = andOp_74_out;
	// controller for notOp_77.notOp_77_in0
	// Insensitive connections
	assign notOp_77_in0 = andOp_76_out;
	// controller for notOp_79.notOp_79_in0
	// Insensitive connections
	assign notOp_79_in0 = icmp_icmp7_out;
	// controller for notOp_82.notOp_82_in0
	// Insensitive connections
	assign notOp_82_in0 = andOp_81_out;
	// controller for notOp_84.notOp_84_in0
	// Insensitive connections
	assign notOp_84_in0 = icmp_icmp7_out;
	// controller for notOp_87.notOp_87_in0
	// Insensitive connections
	assign notOp_87_in0 = andOp_86_out;
	// controller for notOp_89.notOp_89_in0
	// Insensitive connections
	assign notOp_89_in0 = icmp_icmp7_out;
	// controller for notOp_92.notOp_92_in0
	// Insensitive connections
	assign notOp_92_in0 = andOp_91_out;
	// controller for notOp_94.notOp_94_in0
	// Insensitive connections
	assign notOp_94_in0 = icmp_icmp7_out;
	// controller for notOp_97.notOp_97_in0
	// Insensitive connections
	assign notOp_97_in0 = andOp_96_out;
	// controller for notOp_99.notOp_99_in0
	// Insensitive connections
	assign notOp_99_in0 = icmp_icmp7_out;
	// controller for orOp_119.orOp_119_in0
	// controller for orOp_119.orOp_119_in1
	// Insensitive connections
	assign orOp_119_in0 = eq_118_out;
	assign orOp_119_in1 = andOp_74_out;
	// controller for orOp_126.orOp_126_in0
	// controller for orOp_126.orOp_126_in1
	// Insensitive connections
	assign orOp_126_in0 = eq_125_out;
	assign orOp_126_in1 = andOp_78_out;
	// controller for orOp_225.orOp_225_in0
	// controller for orOp_225.orOp_225_in1
	// Insensitive connections
	assign orOp_225_in0 = state_1_is_active;
	assign orOp_225_in1 = 1'd0;
	// controller for orOp_226.orOp_226_in0
	// controller for orOp_226.orOp_226_in1
	// Insensitive connections
	assign orOp_226_in0 = state_2_is_active;
	assign orOp_226_in1 = orOp_225_out;
	// controller for orOp_227.orOp_227_in0
	// controller for orOp_227.orOp_227_in1
	// Insensitive connections
	assign orOp_227_in0 = state_3_is_active;
	assign orOp_227_in1 = orOp_226_out;
	// controller for orOp_228.orOp_228_in0
	// controller for orOp_228.orOp_228_in1
	// Insensitive connections
	assign orOp_228_in0 = state_4_is_active;
	assign orOp_228_in1 = orOp_227_out;
	// controller for orOp_229.orOp_229_in0
	// controller for orOp_229.orOp_229_in1
	// Insensitive connections
	assign orOp_229_in0 = state_5_is_active;
	assign orOp_229_in1 = orOp_228_out;
	// controller for orOp_230.orOp_230_in0
	// controller for orOp_230.orOp_230_in1
	// Insensitive connections
	assign orOp_230_in0 = state_6_is_active;
	assign orOp_230_in1 = orOp_229_out;
	// controller for orOp_231.orOp_231_in0
	// controller for orOp_231.orOp_231_in1
	// Insensitive connections
	assign orOp_231_in0 = state_7_is_active;
	assign orOp_231_in1 = orOp_230_out;
	// controller for phi_phi3.phi_phi3_in
	// controller for phi_phi3.phi_phi3_last_block
	// controller for phi_phi3.phi_phi3_s
	// Insensitive connections
	assign phi_phi3_in = concat_146_out;
	assign phi_phi3_last_block = bb_1_predecessor_in_state_1_out_data;
	assign phi_phi3_s = concat_147_out;
	// controller for phi_phi4.phi_phi4_in
	// controller for phi_phi4.phi_phi4_last_block
	// controller for phi_phi4.phi_phi4_s
	// Insensitive connections
	assign phi_phi4_in = concat_149_out;
	assign phi_phi4_last_block = bb_4_predecessor_in_state_1_out_data;
	assign phi_phi4_s = concat_150_out;
	// controller for ret20.valid_reg
	always @(*) begin
		if (andOp_164_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// controller for shl_shl2.shl_shl2_in0
	// controller for shl_shl2.shl_shl2_in1
	// Insensitive connections
	assign shl_shl2_in0 = phi_phi3_out;
	assign shl_shl2_in1 = 32'd4;
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			data_store_0_0 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_0 <= data_in_0_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_2 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_2 <= data_in_0_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_4 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_4 <= data_in_0_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_6 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_6 <= data_in_0_7_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_10 <= 0;
		end else begin
			if (andOp_236_out) begin
				data_store_1_10 <= shl_shl2_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_12 <= 0;
		end else begin
			if (andOp_237_out) begin
				data_store_1_12 <= phi_phi3_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_14 <= 0;
		end else begin
			if (andOp_238_out) begin
				data_store_1_14 <= phi_phi4_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_15 <= 0;
		end else begin
			if (andOp_239_out) begin
				data_store_1_15 <= add_add6_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_8 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_8 <= data_in_1_9_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_17 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_17 <= data_in_2_18_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_19 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_19 <= data_in_2_20_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_21 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_21 <= data_in_2_22_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_24 <= 0;
		end else begin
			if (andOp_242_out) begin
				data_store_2_24 <= add_add8_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_25 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_25 <= data_in_2_26_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_27 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_27 <= data_in_3_28_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_29 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_29 <= data_in_3_30_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_31 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_31 <= data_in_3_32_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_33 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_33 <= data_in_3_34_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_35 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_35 <= data_in_3_36_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_37 <= 0;
		end else begin
			if (andOp_245_out) begin
				data_store_3_37 <= a_rdata_0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_38 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_38 <= data_in_4_39_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_40 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_40 <= data_in_4_41_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_42 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_42 <= data_in_4_43_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_45 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_45 <= data_in_4_46_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_48 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_48 <= data_in_5_49_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_50 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_50 <= data_in_5_51_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_52 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_52 <= data_in_5_53_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_54 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_54 <= data_in_5_55_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_56 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_56 <= data_in_6_57_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_58 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_58 <= data_in_6_59_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_60 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_60 <= data_in_6_61_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_62 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_62 <= data_in_6_63_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_7_64 <= 0;
		end else begin
			if (andOp_255_out) begin
				data_store_7_64 <= add_add17_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_7_66 <= 0;
		end else begin
			if (state_7_is_active) begin
				data_store_7_66 <= data_in_7_67_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_7_68 <= 0;
		end else begin
			if (state_7_is_active) begin
				data_store_7_68 <= data_in_7_69_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_7_70 <= 0;
		end else begin
			if (state_7_is_active) begin
				data_store_7_70 <= data_in_7_71_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_184_out) begin
				global_state <= 32'd8;
			end
			if (andOp_200_out) begin
				global_state <= 32'd8;
			end
			if (andOp_72_out) begin
				global_state <= 32'd200000;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			out_of_pipe_7_8 <= 0;
		end else begin
			if (andOp_108_out) begin
				out_of_pipe_7_8 <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			out_of_pipe_bb_7_8 <= 0;
		end else begin
			if (andOp_108_out) begin
				out_of_pipe_bb_7_8 <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (1'd1) begin
				state_0_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_110_out) begin
				state_1_entry_BB_reg <= 32'd1;
			end
			if (andOp_72_out) begin
				state_1_entry_BB_reg <= 32'd1;
			end
			if (andOp_80_out) begin
				state_1_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_110_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_206_out) begin
				state_1_is_active <= 1'd0;
			end
			if (andOp_72_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_80_out) begin
				state_1_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_110_out) begin
				state_1_last_BB_reg <= 32'd3;
			end
			if (andOp_72_out) begin
				state_1_last_BB_reg <= 32'd0;
			end
			if (andOp_80_out) begin
				state_1_last_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_110_out) begin
				state_1_last_state <= 32'd7;
			end
			if (andOp_72_out) begin
				state_1_last_state <= 32'd0;
			end
			if (andOp_80_out) begin
				state_1_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_165_out) begin
				state_2_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_165_out) begin
				state_2_is_active <= 1'd1;
			end
			if (andOp_208_out) begin
				state_2_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_165_out) begin
				state_2_last_BB_reg <= bb_4_predecessor_in_state_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_165_out) begin
				state_2_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_166_out) begin
				state_3_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_166_out) begin
				state_3_is_active <= 1'd1;
			end
			if (andOp_210_out) begin
				state_3_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_166_out) begin
				state_3_last_BB_reg <= bb_4_predecessor_in_state_2_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_state <= 0;
		end else begin
			if (andOp_166_out) begin
				state_3_last_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_167_out) begin
				state_4_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_167_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_212_out) begin
				state_4_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_167_out) begin
				state_4_last_BB_reg <= bb_4_predecessor_in_state_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_state <= 0;
		end else begin
			if (andOp_167_out) begin
				state_4_last_state <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_entry_BB_reg <= 0;
		end else begin
			if (andOp_168_out) begin
				state_5_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_is_active <= 0;
		end else begin
			if (andOp_168_out) begin
				state_5_is_active <= 1'd1;
			end
			if (andOp_214_out) begin
				state_5_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_last_BB_reg <= 0;
		end else begin
			if (andOp_168_out) begin
				state_5_last_BB_reg <= bb_4_predecessor_in_state_4_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_last_state <= 0;
		end else begin
			if (andOp_168_out) begin
				state_5_last_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_entry_BB_reg <= 0;
		end else begin
			if (andOp_169_out) begin
				state_6_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_is_active <= 0;
		end else begin
			if (andOp_169_out) begin
				state_6_is_active <= 1'd1;
			end
			if (andOp_216_out) begin
				state_6_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_last_BB_reg <= 0;
		end else begin
			if (andOp_169_out) begin
				state_6_last_BB_reg <= bb_4_predecessor_in_state_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_last_state <= 0;
		end else begin
			if (andOp_169_out) begin
				state_6_last_state <= 32'd5;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_entry_BB_reg <= 0;
		end else begin
			if (andOp_170_out) begin
				state_7_entry_BB_reg <= 32'd4;
			end
			if (andOp_78_out) begin
				state_7_entry_BB_reg <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_is_active <= 0;
		end else begin
			if (andOp_170_out) begin
				state_7_is_active <= 1'd1;
			end
			if (andOp_220_out) begin
				state_7_is_active <= 1'd0;
			end
			if (andOp_78_out) begin
				state_7_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_last_BB_reg <= 0;
		end else begin
			if (andOp_170_out) begin
				state_7_last_BB_reg <= bb_4_predecessor_in_state_6_out_data;
			end
			if (andOp_78_out) begin
				state_7_last_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_last_state <= 0;
		end else begin
			if (andOp_170_out) begin
				state_7_last_state <= 32'd6;
			end
			if (andOp_78_out) begin
				state_7_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_8_entry_BB_reg <= 0;
		end else begin
			if (andOp_199_out) begin
				state_8_entry_BB_reg <= 32'd2;
			end
			if (andOp_200_out) begin
				state_8_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_8_is_active <= 0;
		end else begin
			if (andOp_185_out) begin
				state_8_is_active <= 1'd1;
			end
			if (andOp_200_out) begin
				state_8_is_active <= 1'd1;
			end
			if (andOp_224_out) begin
				state_8_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_8_last_BB_reg <= 0;
		end else begin
			if (andOp_108_out) begin
				state_8_last_BB_reg <= 32'd3;
			end
			if (andOp_200_out) begin
				state_8_last_BB_reg <= bb_2_predecessor_in_state_8_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_8_last_state <= 0;
		end else begin
			if (andOp_108_out) begin
				state_8_last_state <= 32'd7;
			end
			if (andOp_200_out) begin
				state_8_last_state <= 32'd8;
			end
		end
	end

endmodule

