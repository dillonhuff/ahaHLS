module mvmul(input [0:0] clk, input [0:0] rst, output [0:0] valid, output [4:0] ram_debug_addr, input [31:0] ram_debug_data, output [4:0] ram_debug_write_addr, output [31:0] ram_debug_write_data, output [0:0] ram_debug_write_en, output [4:0] ram_raddr_0, output [4:0] ram_raddr_1, output [4:0] ram_raddr_2, input [31:0] ram_rdata_0, input [31:0] ram_rdata_1, input [31:0] ram_rdata_2, output [0:0] ram_rst, output [4:0] ram_waddr_0, output [31:0] ram_wdata_0, output [0:0] ram_wen_0);

	reg [0:0] valid_reg;
	reg [4:0] ram_debug_addr_reg;
	reg [4:0] ram_debug_write_addr_reg;
	reg [31:0] ram_debug_write_data_reg;
	reg [0:0] ram_debug_write_en_reg;
	reg [4:0] ram_raddr_0_reg;
	reg [4:0] ram_raddr_1_reg;
	reg [4:0] ram_raddr_2_reg;
	reg [0:0] ram_rst_reg;
	reg [4:0] ram_waddr_0_reg;
	reg [31:0] ram_wdata_0_reg;
	reg [0:0] ram_wen_0_reg;

	assign valid = valid_reg;
	assign ram_debug_addr = ram_debug_addr_reg;
	assign ram_debug_write_addr = ram_debug_write_addr_reg;
	assign ram_debug_write_data = ram_debug_write_data_reg;
	assign ram_debug_write_en = ram_debug_write_en_reg;
	assign ram_raddr_0 = ram_raddr_0_reg;
	assign ram_raddr_1 = ram_raddr_1_reg;
	assign ram_raddr_2 = ram_raddr_2_reg;
	assign ram_rst = ram_rst_reg;
	assign ram_waddr_0 = ram_waddr_0_reg;
	assign ram_wdata_0 = ram_wdata_0_reg;
	assign ram_wen_0 = ram_wen_0_reg;

	// Start debug wires and ports

	initial begin
	end






	// End debug wires and ports

	// Start Functional Units
	wire [63:0] phi_phi1_in;
	wire [31:0] phi_phi1_last_block;
	wire [63:0] phi_phi1_s;
	wire [31:0] phi_phi1_out;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_phi1(.in(phi_phi1_in), .last_block(phi_phi1_last_block), .out(phi_phi1_out), .s(phi_phi1_s));

	br_dummy br_unit();

	wire [31:0] add_add13_in0;
	wire [31:0] add_add13_in1;
	wire [31:0] add_add13_out;
	add #(.WIDTH(32)) add_add13(.in0(add_add13_in0), .in1(add_add13_in1), .out(add_add13_out));

	wire [31:0] add_add3_in0;
	wire [31:0] add_add3_in1;
	wire [31:0] add_add3_out;
	add #(.WIDTH(32)) add_add3(.in0(add_add3_in0), .in1(add_add3_in1), .out(add_add3_out));

	wire [31:0] icmp_icmp4_in0;
	wire [31:0] icmp_icmp4_in1;
	wire [0:0] icmp_icmp4_out;
	eq #(.WIDTH(32)) icmp_icmp4(.in0(icmp_icmp4_in0), .in1(icmp_icmp4_in1), .out(icmp_icmp4_out));

	wire [31:0] add_add20_in0;
	wire [31:0] add_add20_in1;
	wire [31:0] add_add20_out;
	add #(.WIDTH(32)) add_add20(.in0(add_add20_in0), .in1(add_add20_in1), .out(add_add20_out));

	wire [31:0] mul_mul5_in0;
	wire [31:0] mul_mul5_in1;
	wire [31:0] mul_mul5_out;
	mul #(.WIDTH(32)) mul_mul5(.in0(mul_mul5_in0), .in1(mul_mul5_in1), .out(mul_mul5_out));

	wire [31:0] add_add21_in0;
	wire [31:0] add_add21_in1;
	wire [31:0] add_add21_out;
	add #(.WIDTH(32)) add_add21(.in0(add_add21_in0), .in1(add_add21_in1), .out(add_add21_out));

	wire [31:0] icmp_icmp22_in0;
	wire [31:0] icmp_icmp22_in1;
	wire [0:0] icmp_icmp22_out;
	eq #(.WIDTH(32)) icmp_icmp22(.in0(icmp_icmp22_in0), .in1(icmp_icmp22_in1), .out(icmp_icmp22_out));

	wire [63:0] phi_phi6_in;
	wire [31:0] phi_phi6_last_block;
	wire [63:0] phi_phi6_s;
	wire [31:0] phi_phi6_out;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_phi6(.in(phi_phi6_in), .last_block(phi_phi6_last_block), .out(phi_phi6_out), .s(phi_phi6_s));

	wire [31:0] add_add7_in0;
	wire [31:0] add_add7_in1;
	wire [31:0] add_add7_out;
	add #(.WIDTH(32)) add_add7(.in0(add_add7_in0), .in1(add_add7_in1), .out(add_add7_out));

	wire [31:0] mul_mul16_in0;
	wire [31:0] mul_mul16_in1;
	wire [31:0] mul_mul16_out;
	mul #(.WIDTH(32)) mul_mul16(.in0(mul_mul16_in0), .in1(mul_mul16_in1), .out(mul_mul16_out));

	wire [63:0] phi_phi9_in;
	wire [31:0] phi_phi9_last_block;
	wire [63:0] phi_phi9_s;
	wire [31:0] phi_phi9_out;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_phi9(.in(phi_phi9_in), .last_block(phi_phi9_last_block), .out(phi_phi9_out), .s(phi_phi9_s));

	wire [31:0] add_add12_in0;
	wire [31:0] add_add12_in1;
	wire [31:0] add_add12_out;
	add #(.WIDTH(32)) add_add12(.in0(add_add12_in0), .in1(add_add12_in1), .out(add_add12_out));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] bb_1_active_in_state_0_in_data;
	wire [0:0] bb_1_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_0(.in_data(bb_1_active_in_state_0_in_data), .out_data(bb_1_active_in_state_0_out_data));

	reg [31:0] bb_1_predecessor_in_state_0_in_data;
	wire [31:0] bb_1_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_0(.in_data(bb_1_predecessor_in_state_0_in_data), .out_data(bb_1_predecessor_in_state_0_out_data));

	reg [0:0] br_1_happened_in_state_0_in_data;
	wire [0:0] br_1_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened_in_state_0(.in_data(br_1_happened_in_state_0_in_data), .out_data(br_1_happened_in_state_0_out_data));

	reg [0:0] bb_4_active_in_state_0_in_data;
	wire [0:0] bb_4_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_0(.in_data(bb_4_active_in_state_0_in_data), .out_data(bb_4_active_in_state_0_out_data));

	reg [31:0] bb_4_predecessor_in_state_0_in_data;
	wire [31:0] bb_4_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_0(.in_data(bb_4_predecessor_in_state_0_in_data), .out_data(bb_4_predecessor_in_state_0_out_data));

	reg [0:0] br_4_happened_in_state_0_in_data;
	wire [0:0] br_4_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_0(.in_data(br_4_happened_in_state_0_in_data), .out_data(br_4_happened_in_state_0_out_data));

	reg [0:0] bb_4_active_in_state_1_in_data;
	wire [0:0] bb_4_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_1(.in_data(bb_4_active_in_state_1_in_data), .out_data(bb_4_active_in_state_1_out_data));

	reg [31:0] bb_4_predecessor_in_state_1_in_data;
	wire [31:0] bb_4_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_1(.in_data(bb_4_predecessor_in_state_1_in_data), .out_data(bb_4_predecessor_in_state_1_out_data));

	reg [0:0] br_4_happened_in_state_1_in_data;
	wire [0:0] br_4_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_1(.in_data(br_4_happened_in_state_1_in_data), .out_data(br_4_happened_in_state_1_out_data));

	reg [0:0] bb_4_active_in_state_2_in_data;
	wire [0:0] bb_4_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_2(.in_data(bb_4_active_in_state_2_in_data), .out_data(bb_4_active_in_state_2_out_data));

	reg [31:0] bb_4_predecessor_in_state_2_in_data;
	wire [31:0] bb_4_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_2(.in_data(bb_4_predecessor_in_state_2_in_data), .out_data(bb_4_predecessor_in_state_2_out_data));

	reg [0:0] br_4_happened_in_state_2_in_data;
	wire [0:0] br_4_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_2(.in_data(br_4_happened_in_state_2_in_data), .out_data(br_4_happened_in_state_2_out_data));

	reg [0:0] bb_3_active_in_state_3_in_data;
	wire [0:0] bb_3_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_3(.in_data(bb_3_active_in_state_3_in_data), .out_data(bb_3_active_in_state_3_out_data));

	reg [31:0] bb_3_predecessor_in_state_3_in_data;
	wire [31:0] bb_3_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_3(.in_data(bb_3_predecessor_in_state_3_in_data), .out_data(bb_3_predecessor_in_state_3_out_data));

	reg [0:0] br_3_happened_in_state_3_in_data;
	wire [0:0] br_3_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_3(.in_data(br_3_happened_in_state_3_in_data), .out_data(br_3_happened_in_state_3_out_data));

	reg [0:0] bb_3_active_in_state_4_in_data;
	wire [0:0] bb_3_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_4(.in_data(bb_3_active_in_state_4_in_data), .out_data(bb_3_active_in_state_4_out_data));

	reg [31:0] bb_3_predecessor_in_state_4_in_data;
	wire [31:0] bb_3_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_4(.in_data(bb_3_predecessor_in_state_4_in_data), .out_data(bb_3_predecessor_in_state_4_out_data));

	reg [0:0] br_3_happened_in_state_4_in_data;
	wire [0:0] br_3_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_4(.in_data(br_3_happened_in_state_4_in_data), .out_data(br_3_happened_in_state_4_out_data));

	reg [0:0] bb_3_active_in_state_5_in_data;
	wire [0:0] bb_3_active_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_5(.in_data(bb_3_active_in_state_5_in_data), .out_data(bb_3_active_in_state_5_out_data));

	reg [31:0] bb_3_predecessor_in_state_5_in_data;
	wire [31:0] bb_3_predecessor_in_state_5_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_5(.in_data(bb_3_predecessor_in_state_5_in_data), .out_data(bb_3_predecessor_in_state_5_out_data));

	reg [0:0] br_3_happened_in_state_5_in_data;
	wire [0:0] br_3_happened_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_5(.in_data(br_3_happened_in_state_5_in_data), .out_data(br_3_happened_in_state_5_out_data));

	reg [0:0] bb_3_active_in_state_6_in_data;
	wire [0:0] bb_3_active_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_6(.in_data(bb_3_active_in_state_6_in_data), .out_data(bb_3_active_in_state_6_out_data));

	reg [31:0] bb_3_predecessor_in_state_6_in_data;
	wire [31:0] bb_3_predecessor_in_state_6_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_6(.in_data(bb_3_predecessor_in_state_6_in_data), .out_data(bb_3_predecessor_in_state_6_out_data));

	reg [0:0] br_3_happened_in_state_6_in_data;
	wire [0:0] br_3_happened_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_6(.in_data(br_3_happened_in_state_6_in_data), .out_data(br_3_happened_in_state_6_out_data));

	reg [0:0] bb_2_active_in_state_6_in_data;
	wire [0:0] bb_2_active_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_6(.in_data(bb_2_active_in_state_6_in_data), .out_data(bb_2_active_in_state_6_out_data));

	reg [31:0] bb_2_predecessor_in_state_6_in_data;
	wire [31:0] bb_2_predecessor_in_state_6_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_6(.in_data(bb_2_predecessor_in_state_6_in_data), .out_data(bb_2_predecessor_in_state_6_out_data));

	reg [31:0] data_in_0_1_in_data;
	wire [31:0] data_in_0_1_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_1(.in_data(data_in_0_1_in_data), .out_data(data_in_0_1_out_data));

	reg [31:0] data_in_0_2_in_data;
	wire [31:0] data_in_0_2_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_2(.in_data(data_in_0_2_in_data), .out_data(data_in_0_2_out_data));

	reg [31:0] data_in_0_4_in_data;
	wire [31:0] data_in_0_4_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_4(.in_data(data_in_0_4_in_data), .out_data(data_in_0_4_out_data));

	reg [31:0] data_in_0_7_in_data;
	wire [31:0] data_in_0_7_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_7(.in_data(data_in_0_7_in_data), .out_data(data_in_0_7_out_data));

	reg [31:0] data_in_0_9_in_data;
	wire [31:0] data_in_0_9_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_9(.in_data(data_in_0_9_in_data), .out_data(data_in_0_9_out_data));

	reg [31:0] data_in_1_14_in_data;
	wire [31:0] data_in_1_14_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_14(.in_data(data_in_1_14_in_data), .out_data(data_in_1_14_out_data));

	reg [31:0] data_in_1_16_in_data;
	wire [31:0] data_in_1_16_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_16(.in_data(data_in_1_16_in_data), .out_data(data_in_1_16_out_data));

	reg [0:0] data_in_1_18_in_data;
	wire [0:0] data_in_1_18_out_data;
	hls_wire #(.WIDTH(1)) data_in_1_18(.in_data(data_in_1_18_in_data), .out_data(data_in_1_18_out_data));

	reg [31:0] data_in_1_20_in_data;
	wire [31:0] data_in_1_20_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_20(.in_data(data_in_1_20_in_data), .out_data(data_in_1_20_out_data));

	reg [31:0] data_in_1_22_in_data;
	wire [31:0] data_in_1_22_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_22(.in_data(data_in_1_22_in_data), .out_data(data_in_1_22_out_data));

	reg [31:0] data_in_1_23_in_data;
	wire [31:0] data_in_1_23_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_23(.in_data(data_in_1_23_in_data), .out_data(data_in_1_23_out_data));

	reg [31:0] data_in_1_25_in_data;
	wire [31:0] data_in_1_25_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_25(.in_data(data_in_1_25_in_data), .out_data(data_in_1_25_out_data));

	reg [31:0] data_in_2_26_in_data;
	wire [31:0] data_in_2_26_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_26(.in_data(data_in_2_26_in_data), .out_data(data_in_2_26_out_data));

	reg [31:0] data_in_2_28_in_data;
	wire [31:0] data_in_2_28_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_28(.in_data(data_in_2_28_in_data), .out_data(data_in_2_28_out_data));

	reg [31:0] data_in_2_31_in_data;
	wire [31:0] data_in_2_31_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_31(.in_data(data_in_2_31_in_data), .out_data(data_in_2_31_out_data));

	reg [0:0] data_in_2_32_in_data;
	wire [0:0] data_in_2_32_out_data;
	hls_wire #(.WIDTH(1)) data_in_2_32(.in_data(data_in_2_32_in_data), .out_data(data_in_2_32_out_data));

	reg [31:0] data_in_2_34_in_data;
	wire [31:0] data_in_2_34_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_34(.in_data(data_in_2_34_in_data), .out_data(data_in_2_34_out_data));

	reg [31:0] data_in_2_36_in_data;
	wire [31:0] data_in_2_36_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_36(.in_data(data_in_2_36_in_data), .out_data(data_in_2_36_out_data));

	reg [31:0] data_in_2_37_in_data;
	wire [31:0] data_in_2_37_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_37(.in_data(data_in_2_37_in_data), .out_data(data_in_2_37_out_data));

	reg [31:0] data_in_3_39_in_data;
	wire [31:0] data_in_3_39_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_39(.in_data(data_in_3_39_in_data), .out_data(data_in_3_39_out_data));

	reg [31:0] data_in_3_41_in_data;
	wire [31:0] data_in_3_41_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_41(.in_data(data_in_3_41_in_data), .out_data(data_in_3_41_out_data));

	reg [31:0] data_in_3_43_in_data;
	wire [31:0] data_in_3_43_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_43(.in_data(data_in_3_43_in_data), .out_data(data_in_3_43_out_data));

	reg [31:0] data_in_3_45_in_data;
	wire [31:0] data_in_3_45_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_45(.in_data(data_in_3_45_in_data), .out_data(data_in_3_45_out_data));

	reg [31:0] data_in_4_49_in_data;
	wire [31:0] data_in_4_49_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_49(.in_data(data_in_4_49_in_data), .out_data(data_in_4_49_out_data));

	reg [31:0] data_in_4_51_in_data;
	wire [31:0] data_in_4_51_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_51(.in_data(data_in_4_51_in_data), .out_data(data_in_4_51_out_data));

	reg [31:0] data_in_4_53_in_data;
	wire [31:0] data_in_4_53_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_53(.in_data(data_in_4_53_in_data), .out_data(data_in_4_53_out_data));

	reg [31:0] data_in_4_55_in_data;
	wire [31:0] data_in_4_55_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_55(.in_data(data_in_4_55_in_data), .out_data(data_in_4_55_out_data));

	reg [31:0] data_in_4_57_in_data;
	wire [31:0] data_in_4_57_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_57(.in_data(data_in_4_57_in_data), .out_data(data_in_4_57_out_data));

	reg [0:0] data_in_4_59_in_data;
	wire [0:0] data_in_4_59_out_data;
	hls_wire #(.WIDTH(1)) data_in_4_59(.in_data(data_in_4_59_in_data), .out_data(data_in_4_59_out_data));

	reg [31:0] data_in_5_61_in_data;
	wire [31:0] data_in_5_61_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_61(.in_data(data_in_5_61_in_data), .out_data(data_in_5_61_out_data));

	reg [31:0] data_in_5_63_in_data;
	wire [31:0] data_in_5_63_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_63(.in_data(data_in_5_63_in_data), .out_data(data_in_5_63_out_data));

	reg [31:0] data_in_5_65_in_data;
	wire [31:0] data_in_5_65_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_65(.in_data(data_in_5_65_in_data), .out_data(data_in_5_65_out_data));

	reg [31:0] data_in_5_67_in_data;
	wire [31:0] data_in_5_67_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_67(.in_data(data_in_5_67_in_data), .out_data(data_in_5_67_out_data));

	reg [31:0] data_in_5_69_in_data;
	wire [31:0] data_in_5_69_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_69(.in_data(data_in_5_69_in_data), .out_data(data_in_5_69_out_data));

	reg [0:0] data_in_5_71_in_data;
	wire [0:0] data_in_5_71_out_data;
	hls_wire #(.WIDTH(1)) data_in_5_71(.in_data(data_in_5_71_in_data), .out_data(data_in_5_71_out_data));

	reg [31:0] data_in_6_73_in_data;
	wire [31:0] data_in_6_73_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_73(.in_data(data_in_6_73_in_data), .out_data(data_in_6_73_out_data));

	reg [31:0] data_in_6_75_in_data;
	wire [31:0] data_in_6_75_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_75(.in_data(data_in_6_75_in_data), .out_data(data_in_6_75_out_data));

	reg [31:0] data_in_6_77_in_data;
	wire [31:0] data_in_6_77_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_77(.in_data(data_in_6_77_in_data), .out_data(data_in_6_77_out_data));

	reg [31:0] data_in_6_79_in_data;
	wire [31:0] data_in_6_79_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_79(.in_data(data_in_6_79_in_data), .out_data(data_in_6_79_out_data));

	reg [31:0] data_in_6_81_in_data;
	wire [31:0] data_in_6_81_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_81(.in_data(data_in_6_81_in_data), .out_data(data_in_6_81_out_data));

	reg [0:0] data_in_6_82_in_data;
	wire [0:0] data_in_6_82_out_data;
	hls_wire #(.WIDTH(1)) data_in_6_82(.in_data(data_in_6_82_in_data), .out_data(data_in_6_82_out_data));

	wire [0:0] andOp_83_in0;
	wire [0:0] andOp_83_in1;
	wire [0:0] andOp_83_out;
	andOp #(.WIDTH(1)) andOp_83(.in0(andOp_83_in0), .in1(andOp_83_in1), .out(andOp_83_out));

	wire [0:0] notOp_84_in0;
	wire [0:0] notOp_84_out;
	notOp #(.WIDTH(1)) notOp_84(.in(notOp_84_in0), .out(notOp_84_out));

	wire [0:0] andOp_85_in0;
	wire [0:0] andOp_85_in1;
	wire [0:0] andOp_85_out;
	andOp #(.WIDTH(1)) andOp_85(.in0(andOp_85_in0), .in1(andOp_85_in1), .out(andOp_85_out));

	wire [0:0] notOp_86_in0;
	wire [0:0] notOp_86_out;
	notOp #(.WIDTH(1)) notOp_86(.in(notOp_86_in0), .out(notOp_86_out));

	wire [0:0] andOp_87_in0;
	wire [0:0] andOp_87_in1;
	wire [0:0] andOp_87_out;
	andOp #(.WIDTH(1)) andOp_87(.in0(andOp_87_in0), .in1(andOp_87_in1), .out(andOp_87_out));

	wire [0:0] notOp_88_in0;
	wire [0:0] notOp_88_out;
	notOp #(.WIDTH(1)) notOp_88(.in(notOp_88_in0), .out(notOp_88_out));

	wire [0:0] andOp_89_in0;
	wire [0:0] andOp_89_in1;
	wire [0:0] andOp_89_out;
	andOp #(.WIDTH(1)) andOp_89(.in0(andOp_89_in0), .in1(andOp_89_in1), .out(andOp_89_out));

	wire [0:0] notOp_90_in0;
	wire [0:0] notOp_90_out;
	notOp #(.WIDTH(1)) notOp_90(.in(notOp_90_in0), .out(notOp_90_out));

	wire [0:0] andOp_91_in0;
	wire [0:0] andOp_91_in1;
	wire [0:0] andOp_91_out;
	andOp #(.WIDTH(1)) andOp_91(.in0(andOp_91_in0), .in1(andOp_91_in1), .out(andOp_91_out));

	wire [0:0] andOp_92_in0;
	wire [0:0] andOp_92_in1;
	wire [0:0] andOp_92_out;
	andOp #(.WIDTH(1)) andOp_92(.in0(andOp_92_in0), .in1(andOp_92_in1), .out(andOp_92_out));

	wire [0:0] notOp_93_in0;
	wire [0:0] notOp_93_out;
	notOp #(.WIDTH(1)) notOp_93(.in(notOp_93_in0), .out(notOp_93_out));

	wire [0:0] andOp_94_in0;
	wire [0:0] andOp_94_in1;
	wire [0:0] andOp_94_out;
	andOp #(.WIDTH(1)) andOp_94(.in0(andOp_94_in0), .in1(andOp_94_in1), .out(andOp_94_out));

	wire [0:0] notOp_95_in0;
	wire [0:0] notOp_95_out;
	notOp #(.WIDTH(1)) notOp_95(.in(notOp_95_in0), .out(notOp_95_out));

	wire [0:0] andOp_96_in0;
	wire [0:0] andOp_96_in1;
	wire [0:0] andOp_96_out;
	andOp #(.WIDTH(1)) andOp_96(.in0(andOp_96_in0), .in1(andOp_96_in1), .out(andOp_96_out));

	wire [0:0] andOp_97_in0;
	wire [0:0] andOp_97_in1;
	wire [0:0] andOp_97_out;
	andOp #(.WIDTH(1)) andOp_97(.in0(andOp_97_in0), .in1(andOp_97_in1), .out(andOp_97_out));

	wire [0:0] notOp_98_in0;
	wire [0:0] notOp_98_out;
	notOp #(.WIDTH(1)) notOp_98(.in(notOp_98_in0), .out(notOp_98_out));

	wire [0:0] andOp_99_in0;
	wire [0:0] andOp_99_in1;
	wire [0:0] andOp_99_out;
	andOp #(.WIDTH(1)) andOp_99(.in0(andOp_99_in0), .in1(andOp_99_in1), .out(andOp_99_out));

	wire [0:0] notOp_100_in0;
	wire [0:0] notOp_100_out;
	notOp #(.WIDTH(1)) notOp_100(.in(notOp_100_in0), .out(notOp_100_out));

	wire [0:0] andOp_101_in0;
	wire [0:0] andOp_101_in1;
	wire [0:0] andOp_101_out;
	andOp #(.WIDTH(1)) andOp_101(.in0(andOp_101_in0), .in1(andOp_101_in1), .out(andOp_101_out));

	wire [0:0] andOp_102_in0;
	wire [0:0] andOp_102_in1;
	wire [0:0] andOp_102_out;
	andOp #(.WIDTH(1)) andOp_102(.in0(andOp_102_in0), .in1(andOp_102_in1), .out(andOp_102_out));

	wire [0:0] notOp_103_in0;
	wire [0:0] notOp_103_out;
	notOp #(.WIDTH(1)) notOp_103(.in(notOp_103_in0), .out(notOp_103_out));

	wire [0:0] andOp_104_in0;
	wire [0:0] andOp_104_in1;
	wire [0:0] andOp_104_out;
	andOp #(.WIDTH(1)) andOp_104(.in0(andOp_104_in0), .in1(andOp_104_in1), .out(andOp_104_out));

	wire [0:0] notOp_105_in0;
	wire [0:0] notOp_105_out;
	notOp #(.WIDTH(1)) notOp_105(.in(notOp_105_in0), .out(notOp_105_out));

	wire [0:0] andOp_106_in0;
	wire [0:0] andOp_106_in1;
	wire [0:0] andOp_106_out;
	andOp #(.WIDTH(1)) andOp_106(.in0(andOp_106_in0), .in1(andOp_106_in1), .out(andOp_106_out));

	wire [0:0] andOp_107_in0;
	wire [0:0] andOp_107_in1;
	wire [0:0] andOp_107_out;
	andOp #(.WIDTH(1)) andOp_107(.in0(andOp_107_in0), .in1(andOp_107_in1), .out(andOp_107_out));

	wire [0:0] notOp_108_in0;
	wire [0:0] notOp_108_out;
	notOp #(.WIDTH(1)) notOp_108(.in(notOp_108_in0), .out(notOp_108_out));

	wire [0:0] andOp_109_in0;
	wire [0:0] andOp_109_in1;
	wire [0:0] andOp_109_out;
	andOp #(.WIDTH(1)) andOp_109(.in0(andOp_109_in0), .in1(andOp_109_in1), .out(andOp_109_out));

	wire [0:0] notOp_110_in0;
	wire [0:0] notOp_110_out;
	notOp #(.WIDTH(1)) notOp_110(.in(notOp_110_in0), .out(notOp_110_out));

	wire [0:0] andOp_111_in0;
	wire [0:0] andOp_111_in1;
	wire [0:0] andOp_111_out;
	andOp #(.WIDTH(1)) andOp_111(.in0(andOp_111_in0), .in1(andOp_111_in1), .out(andOp_111_out));

	wire [0:0] andOp_112_in0;
	wire [0:0] andOp_112_in1;
	wire [0:0] andOp_112_out;
	andOp #(.WIDTH(1)) andOp_112(.in0(andOp_112_in0), .in1(andOp_112_in1), .out(andOp_112_out));

	wire [0:0] notOp_113_in0;
	wire [0:0] notOp_113_out;
	notOp #(.WIDTH(1)) notOp_113(.in(notOp_113_in0), .out(notOp_113_out));

	wire [0:0] andOp_114_in0;
	wire [0:0] andOp_114_in1;
	wire [0:0] andOp_114_out;
	andOp #(.WIDTH(1)) andOp_114(.in0(andOp_114_in0), .in1(andOp_114_in1), .out(andOp_114_out));

	wire [0:0] notOp_115_in0;
	wire [0:0] notOp_115_out;
	notOp #(.WIDTH(1)) notOp_115(.in(notOp_115_in0), .out(notOp_115_out));

	wire [0:0] andOp_116_in0;
	wire [0:0] andOp_116_in1;
	wire [0:0] andOp_116_out;
	andOp #(.WIDTH(1)) andOp_116(.in0(andOp_116_in0), .in1(andOp_116_in1), .out(andOp_116_out));

	wire [0:0] andOp_117_in0;
	wire [0:0] andOp_117_in1;
	wire [0:0] andOp_117_out;
	andOp #(.WIDTH(1)) andOp_117(.in0(andOp_117_in0), .in1(andOp_117_in1), .out(andOp_117_out));

	wire [0:0] notOp_118_in0;
	wire [0:0] notOp_118_out;
	notOp #(.WIDTH(1)) notOp_118(.in(notOp_118_in0), .out(notOp_118_out));

	wire [0:0] andOp_119_in0;
	wire [0:0] andOp_119_in1;
	wire [0:0] andOp_119_out;
	andOp #(.WIDTH(1)) andOp_119(.in0(andOp_119_in0), .in1(andOp_119_in1), .out(andOp_119_out));

	wire [0:0] notOp_120_in0;
	wire [0:0] notOp_120_out;
	notOp #(.WIDTH(1)) notOp_120(.in(notOp_120_in0), .out(notOp_120_out));

	wire [0:0] andOp_121_in0;
	wire [0:0] andOp_121_in1;
	wire [0:0] andOp_121_out;
	andOp #(.WIDTH(1)) andOp_121(.in0(andOp_121_in0), .in1(andOp_121_in1), .out(andOp_121_out));

	wire [31:0] eq_122_in0;
	wire [31:0] eq_122_in1;
	wire [0:0] eq_122_out;
	eq #(.WIDTH(32)) eq_122(.in0(eq_122_in0), .in1(eq_122_in1), .out(eq_122_out));

	wire [31:0] eq_123_in0;
	wire [31:0] eq_123_in1;
	wire [0:0] eq_123_out;
	eq #(.WIDTH(32)) eq_123(.in0(eq_123_in0), .in1(eq_123_in1), .out(eq_123_out));

	wire [0:0] orOp_124_in0;
	wire [0:0] orOp_124_in1;
	wire [0:0] orOp_124_out;
	orOp #(.WIDTH(1)) orOp_124(.in0(orOp_124_in0), .in1(orOp_124_in1), .out(orOp_124_out));

	wire [31:0] eq_125_in0;
	wire [31:0] eq_125_in1;
	wire [0:0] eq_125_out;
	eq #(.WIDTH(32)) eq_125(.in0(eq_125_in0), .in1(eq_125_in1), .out(eq_125_out));

	wire [0:0] orOp_126_in0;
	wire [0:0] orOp_126_in1;
	wire [0:0] orOp_126_out;
	orOp #(.WIDTH(1)) orOp_126(.in0(orOp_126_in0), .in1(orOp_126_in1), .out(orOp_126_out));

	wire [31:0] eq_127_in0;
	wire [31:0] eq_127_in1;
	wire [0:0] eq_127_out;
	eq #(.WIDTH(32)) eq_127(.in0(eq_127_in0), .in1(eq_127_in1), .out(eq_127_out));

	wire [31:0] eq_128_in0;
	wire [31:0] eq_128_in1;
	wire [0:0] eq_128_out;
	eq #(.WIDTH(32)) eq_128(.in0(eq_128_in0), .in1(eq_128_in1), .out(eq_128_out));

	wire [31:0] eq_129_in0;
	wire [31:0] eq_129_in1;
	wire [0:0] eq_129_out;
	eq #(.WIDTH(32)) eq_129(.in0(eq_129_in0), .in1(eq_129_in1), .out(eq_129_out));

	wire [31:0] eq_130_in0;
	wire [31:0] eq_130_in1;
	wire [0:0] eq_130_out;
	eq #(.WIDTH(32)) eq_130(.in0(eq_130_in0), .in1(eq_130_in1), .out(eq_130_out));

	wire [31:0] eq_131_in0;
	wire [31:0] eq_131_in1;
	wire [0:0] eq_131_out;
	eq #(.WIDTH(32)) eq_131(.in0(eq_131_in0), .in1(eq_131_in1), .out(eq_131_out));

	wire [31:0] eq_132_in0;
	wire [31:0] eq_132_in1;
	wire [0:0] eq_132_out;
	eq #(.WIDTH(32)) eq_132(.in0(eq_132_in0), .in1(eq_132_in1), .out(eq_132_out));

	wire [31:0] eq_133_in0;
	wire [31:0] eq_133_in1;
	wire [0:0] eq_133_out;
	eq #(.WIDTH(32)) eq_133(.in0(eq_133_in0), .in1(eq_133_in1), .out(eq_133_out));

	wire [0:0] orOp_134_in0;
	wire [0:0] orOp_134_in1;
	wire [0:0] orOp_134_out;
	orOp #(.WIDTH(1)) orOp_134(.in0(orOp_134_in0), .in1(orOp_134_in1), .out(orOp_134_out));

	wire [31:0] eq_135_in0;
	wire [31:0] eq_135_in1;
	wire [0:0] eq_135_out;
	eq #(.WIDTH(32)) eq_135(.in0(eq_135_in0), .in1(eq_135_in1), .out(eq_135_out));

	wire [31:0] eq_136_in0;
	wire [31:0] eq_136_in1;
	wire [0:0] eq_136_out;
	eq #(.WIDTH(32)) eq_136(.in0(eq_136_in0), .in1(eq_136_in1), .out(eq_136_out));

	wire [0:0] notOp_137_in0;
	wire [0:0] notOp_137_out;
	notOp #(.WIDTH(1)) notOp_137(.in(notOp_137_in0), .out(notOp_137_out));

	wire [0:0] andOp_138_in0;
	wire [0:0] andOp_138_in1;
	wire [0:0] andOp_138_out;
	andOp #(.WIDTH(1)) andOp_138(.in0(andOp_138_in0), .in1(andOp_138_in1), .out(andOp_138_out));

	wire [31:0] eq_139_in0;
	wire [31:0] eq_139_in1;
	wire [0:0] eq_139_out;
	eq #(.WIDTH(32)) eq_139(.in0(eq_139_in0), .in1(eq_139_in1), .out(eq_139_out));

	wire [0:0] notOp_140_in0;
	wire [0:0] notOp_140_out;
	notOp #(.WIDTH(1)) notOp_140(.in(notOp_140_in0), .out(notOp_140_out));

	wire [0:0] andOp_141_in0;
	wire [0:0] andOp_141_in1;
	wire [0:0] andOp_141_out;
	andOp #(.WIDTH(1)) andOp_141(.in0(andOp_141_in0), .in1(andOp_141_in1), .out(andOp_141_out));

	wire [31:0] eq_142_in0;
	wire [31:0] eq_142_in1;
	wire [0:0] eq_142_out;
	eq #(.WIDTH(32)) eq_142(.in0(eq_142_in0), .in1(eq_142_in1), .out(eq_142_out));

	wire [31:0] eq_143_in0;
	wire [31:0] eq_143_in1;
	wire [0:0] eq_143_out;
	eq #(.WIDTH(32)) eq_143(.in0(eq_143_in0), .in1(eq_143_in1), .out(eq_143_out));

	wire [31:0] eq_144_in0;
	wire [31:0] eq_144_in1;
	wire [0:0] eq_144_out;
	eq #(.WIDTH(32)) eq_144(.in0(eq_144_in0), .in1(eq_144_in1), .out(eq_144_out));

	wire [31:0] eq_145_in0;
	wire [31:0] eq_145_in1;
	wire [0:0] eq_145_out;
	eq #(.WIDTH(32)) eq_145(.in0(eq_145_in0), .in1(eq_145_in1), .out(eq_145_out));

	wire [31:0] eq_146_in0;
	wire [31:0] eq_146_in1;
	wire [0:0] eq_146_out;
	eq #(.WIDTH(32)) eq_146(.in0(eq_146_in0), .in1(eq_146_in1), .out(eq_146_out));

	wire [31:0] eq_147_in0;
	wire [31:0] eq_147_in1;
	wire [0:0] eq_147_out;
	eq #(.WIDTH(32)) eq_147(.in0(eq_147_in0), .in1(eq_147_in1), .out(eq_147_out));

	wire [31:0] eq_148_in0;
	wire [31:0] eq_148_in1;
	wire [0:0] eq_148_out;
	eq #(.WIDTH(32)) eq_148(.in0(eq_148_in0), .in1(eq_148_in1), .out(eq_148_out));

	wire [0:0] notOp_149_in0;
	wire [0:0] notOp_149_out;
	notOp #(.WIDTH(1)) notOp_149(.in(notOp_149_in0), .out(notOp_149_out));

	wire [0:0] andOp_150_in0;
	wire [0:0] andOp_150_in1;
	wire [0:0] andOp_150_out;
	andOp #(.WIDTH(1)) andOp_150(.in0(andOp_150_in0), .in1(andOp_150_in1), .out(andOp_150_out));

	wire [0:0] andOp_151_in0;
	wire [0:0] andOp_151_in1;
	wire [0:0] andOp_151_out;
	andOp #(.WIDTH(1)) andOp_151(.in0(andOp_151_in0), .in1(andOp_151_in1), .out(andOp_151_out));

	wire [0:0] andOp_152_in0;
	wire [0:0] andOp_152_in1;
	wire [0:0] andOp_152_out;
	andOp #(.WIDTH(1)) andOp_152(.in0(andOp_152_in0), .in1(andOp_152_in1), .out(andOp_152_out));

	wire [0:0] andOp_153_in0;
	wire [0:0] andOp_153_in1;
	wire [0:0] andOp_153_out;
	andOp #(.WIDTH(1)) andOp_153(.in0(andOp_153_in0), .in1(andOp_153_in1), .out(andOp_153_out));

	wire [0:0] andOp_154_in0;
	wire [0:0] andOp_154_in1;
	wire [0:0] andOp_154_out;
	andOp #(.WIDTH(1)) andOp_154(.in0(andOp_154_in0), .in1(andOp_154_in1), .out(andOp_154_out));

	wire [0:0] andOp_155_in0;
	wire [0:0] andOp_155_in1;
	wire [0:0] andOp_155_out;
	andOp #(.WIDTH(1)) andOp_155(.in0(andOp_155_in0), .in1(andOp_155_in1), .out(andOp_155_out));

	wire [0:0] andOp_156_in0;
	wire [0:0] andOp_156_in1;
	wire [0:0] andOp_156_out;
	andOp #(.WIDTH(1)) andOp_156(.in0(andOp_156_in0), .in1(andOp_156_in1), .out(andOp_156_out));

	wire [0:0] andOp_157_in0;
	wire [0:0] andOp_157_in1;
	wire [0:0] andOp_157_out;
	andOp #(.WIDTH(1)) andOp_157(.in0(andOp_157_in0), .in1(andOp_157_in1), .out(andOp_157_out));

	wire [0:0] andOp_158_in0;
	wire [0:0] andOp_158_in1;
	wire [0:0] andOp_158_out;
	andOp #(.WIDTH(1)) andOp_158(.in0(andOp_158_in0), .in1(andOp_158_in1), .out(andOp_158_out));

	wire [31:0] concat_159_in0;
	wire [31:0] concat_159_in1;
	wire [63:0] concat_159_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_159(.in0(concat_159_in0), .in1(concat_159_in1), .out(concat_159_out));

	wire [31:0] concat_160_in0;
	wire [31:0] concat_160_in1;
	wire [63:0] concat_160_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_160(.in0(concat_160_in0), .in1(concat_160_in1), .out(concat_160_out));

	wire [0:0] andOp_161_in0;
	wire [0:0] andOp_161_in1;
	wire [0:0] andOp_161_out;
	andOp #(.WIDTH(1)) andOp_161(.in0(andOp_161_in0), .in1(andOp_161_in1), .out(andOp_161_out));

	wire [0:0] andOp_162_in0;
	wire [0:0] andOp_162_in1;
	wire [0:0] andOp_162_out;
	andOp #(.WIDTH(1)) andOp_162(.in0(andOp_162_in0), .in1(andOp_162_in1), .out(andOp_162_out));

	wire [0:0] andOp_163_in0;
	wire [0:0] andOp_163_in1;
	wire [0:0] andOp_163_out;
	andOp #(.WIDTH(1)) andOp_163(.in0(andOp_163_in0), .in1(andOp_163_in1), .out(andOp_163_out));

	wire [0:0] andOp_164_in0;
	wire [0:0] andOp_164_in1;
	wire [0:0] andOp_164_out;
	andOp #(.WIDTH(1)) andOp_164(.in0(andOp_164_in0), .in1(andOp_164_in1), .out(andOp_164_out));

	wire [31:0] concat_165_in0;
	wire [31:0] concat_165_in1;
	wire [63:0] concat_165_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_165(.in0(concat_165_in0), .in1(concat_165_in1), .out(concat_165_out));

	wire [31:0] concat_166_in0;
	wire [31:0] concat_166_in1;
	wire [63:0] concat_166_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_166(.in0(concat_166_in0), .in1(concat_166_in1), .out(concat_166_out));

	wire [0:0] andOp_167_in0;
	wire [0:0] andOp_167_in1;
	wire [0:0] andOp_167_out;
	andOp #(.WIDTH(1)) andOp_167(.in0(andOp_167_in0), .in1(andOp_167_in1), .out(andOp_167_out));

	wire [0:0] andOp_168_in0;
	wire [0:0] andOp_168_in1;
	wire [0:0] andOp_168_out;
	andOp #(.WIDTH(1)) andOp_168(.in0(andOp_168_in0), .in1(andOp_168_in1), .out(andOp_168_out));

	wire [31:0] concat_169_in0;
	wire [31:0] concat_169_in1;
	wire [63:0] concat_169_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_169(.in0(concat_169_in0), .in1(concat_169_in1), .out(concat_169_out));

	wire [31:0] concat_170_in0;
	wire [31:0] concat_170_in1;
	wire [63:0] concat_170_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_170(.in0(concat_170_in0), .in1(concat_170_in1), .out(concat_170_out));

	wire [0:0] andOp_171_in0;
	wire [0:0] andOp_171_in1;
	wire [0:0] andOp_171_out;
	andOp #(.WIDTH(1)) andOp_171(.in0(andOp_171_in0), .in1(andOp_171_in1), .out(andOp_171_out));

	wire [0:0] andOp_172_in0;
	wire [0:0] andOp_172_in1;
	wire [0:0] andOp_172_out;
	andOp #(.WIDTH(1)) andOp_172(.in0(andOp_172_in0), .in1(andOp_172_in1), .out(andOp_172_out));

	wire [0:0] andOp_173_in0;
	wire [0:0] andOp_173_in1;
	wire [0:0] andOp_173_out;
	andOp #(.WIDTH(1)) andOp_173(.in0(andOp_173_in0), .in1(andOp_173_in1), .out(andOp_173_out));

	wire [0:0] andOp_174_in0;
	wire [0:0] andOp_174_in1;
	wire [0:0] andOp_174_out;
	andOp #(.WIDTH(1)) andOp_174(.in0(andOp_174_in0), .in1(andOp_174_in1), .out(andOp_174_out));

	wire [0:0] andOp_175_in0;
	wire [0:0] andOp_175_in1;
	wire [0:0] andOp_175_out;
	andOp #(.WIDTH(1)) andOp_175(.in0(andOp_175_in0), .in1(andOp_175_in1), .out(andOp_175_out));

	wire [0:0] andOp_176_in0;
	wire [0:0] andOp_176_in1;
	wire [0:0] andOp_176_out;
	andOp #(.WIDTH(1)) andOp_176(.in0(andOp_176_in0), .in1(andOp_176_in1), .out(andOp_176_out));

	wire [0:0] andOp_177_in0;
	wire [0:0] andOp_177_in1;
	wire [0:0] andOp_177_out;
	andOp #(.WIDTH(1)) andOp_177(.in0(andOp_177_in0), .in1(andOp_177_in1), .out(andOp_177_out));

	wire [0:0] andOp_178_in0;
	wire [0:0] andOp_178_in1;
	wire [0:0] andOp_178_out;
	andOp #(.WIDTH(1)) andOp_178(.in0(andOp_178_in0), .in1(andOp_178_in1), .out(andOp_178_out));

	wire [0:0] andOp_179_in0;
	wire [0:0] andOp_179_in1;
	wire [0:0] andOp_179_out;
	andOp #(.WIDTH(1)) andOp_179(.in0(andOp_179_in0), .in1(andOp_179_in1), .out(andOp_179_out));

	wire [0:0] andOp_180_in0;
	wire [0:0] andOp_180_in1;
	wire [0:0] andOp_180_out;
	andOp #(.WIDTH(1)) andOp_180(.in0(andOp_180_in0), .in1(andOp_180_in1), .out(andOp_180_out));

	wire [0:0] andOp_181_in0;
	wire [0:0] andOp_181_in1;
	wire [0:0] andOp_181_out;
	andOp #(.WIDTH(1)) andOp_181(.in0(andOp_181_in0), .in1(andOp_181_in1), .out(andOp_181_out));

	wire [0:0] andOp_182_in0;
	wire [0:0] andOp_182_in1;
	wire [0:0] andOp_182_out;
	andOp #(.WIDTH(1)) andOp_182(.in0(andOp_182_in0), .in1(andOp_182_in1), .out(andOp_182_out));

	wire [0:0] andOp_183_in0;
	wire [0:0] andOp_183_in1;
	wire [0:0] andOp_183_out;
	andOp #(.WIDTH(1)) andOp_183(.in0(andOp_183_in0), .in1(andOp_183_in1), .out(andOp_183_out));

	wire [0:0] notOp_184_in0;
	wire [0:0] notOp_184_out;
	notOp #(.WIDTH(1)) notOp_184(.in(notOp_184_in0), .out(notOp_184_out));

	wire [0:0] andOp_185_in0;
	wire [0:0] andOp_185_in1;
	wire [0:0] andOp_185_out;
	andOp #(.WIDTH(1)) andOp_185(.in0(andOp_185_in0), .in1(andOp_185_in1), .out(andOp_185_out));

	wire [0:0] notOp_186_in0;
	wire [0:0] notOp_186_out;
	notOp #(.WIDTH(1)) notOp_186(.in(notOp_186_in0), .out(notOp_186_out));

	wire [0:0] andOp_187_in0;
	wire [0:0] andOp_187_in1;
	wire [0:0] andOp_187_out;
	andOp #(.WIDTH(1)) andOp_187(.in0(andOp_187_in0), .in1(andOp_187_in1), .out(andOp_187_out));

	wire [0:0] notOp_188_in0;
	wire [0:0] notOp_188_out;
	notOp #(.WIDTH(1)) notOp_188(.in(notOp_188_in0), .out(notOp_188_out));

	wire [0:0] andOp_189_in0;
	wire [0:0] andOp_189_in1;
	wire [0:0] andOp_189_out;
	andOp #(.WIDTH(1)) andOp_189(.in0(andOp_189_in0), .in1(andOp_189_in1), .out(andOp_189_out));

	wire [0:0] notOp_190_in0;
	wire [0:0] notOp_190_out;
	notOp #(.WIDTH(1)) notOp_190(.in(notOp_190_in0), .out(notOp_190_out));

	wire [0:0] andOp_191_in0;
	wire [0:0] andOp_191_in1;
	wire [0:0] andOp_191_out;
	andOp #(.WIDTH(1)) andOp_191(.in0(andOp_191_in0), .in1(andOp_191_in1), .out(andOp_191_out));

	wire [0:0] notOp_192_in0;
	wire [0:0] notOp_192_out;
	notOp #(.WIDTH(1)) notOp_192(.in(notOp_192_in0), .out(notOp_192_out));

	wire [0:0] andOp_193_in0;
	wire [0:0] andOp_193_in1;
	wire [0:0] andOp_193_out;
	andOp #(.WIDTH(1)) andOp_193(.in0(andOp_193_in0), .in1(andOp_193_in1), .out(andOp_193_out));

	wire [0:0] notOp_194_in0;
	wire [0:0] notOp_194_out;
	notOp #(.WIDTH(1)) notOp_194(.in(notOp_194_in0), .out(notOp_194_out));

	wire [0:0] andOp_195_in0;
	wire [0:0] andOp_195_in1;
	wire [0:0] andOp_195_out;
	andOp #(.WIDTH(1)) andOp_195(.in0(andOp_195_in0), .in1(andOp_195_in1), .out(andOp_195_out));

	wire [0:0] notOp_196_in0;
	wire [0:0] notOp_196_out;
	notOp #(.WIDTH(1)) notOp_196(.in(notOp_196_in0), .out(notOp_196_out));

	wire [0:0] andOp_197_in0;
	wire [0:0] andOp_197_in1;
	wire [0:0] andOp_197_out;
	andOp #(.WIDTH(1)) andOp_197(.in0(andOp_197_in0), .in1(andOp_197_in1), .out(andOp_197_out));

	wire [0:0] notOp_198_in0;
	wire [0:0] notOp_198_out;
	notOp #(.WIDTH(1)) notOp_198(.in(notOp_198_in0), .out(notOp_198_out));

	wire [0:0] andOp_199_in0;
	wire [0:0] andOp_199_in1;
	wire [0:0] andOp_199_out;
	andOp #(.WIDTH(1)) andOp_199(.in0(andOp_199_in0), .in1(andOp_199_in1), .out(andOp_199_out));

	wire [0:0] notOp_200_in0;
	wire [0:0] notOp_200_out;
	notOp #(.WIDTH(1)) notOp_200(.in(notOp_200_in0), .out(notOp_200_out));

	wire [0:0] andOp_201_in0;
	wire [0:0] andOp_201_in1;
	wire [0:0] andOp_201_out;
	andOp #(.WIDTH(1)) andOp_201(.in0(andOp_201_in0), .in1(andOp_201_in1), .out(andOp_201_out));

	wire [31:0] eq_202_in0;
	wire [31:0] eq_202_in1;
	wire [0:0] eq_202_out;
	eq #(.WIDTH(32)) eq_202(.in0(eq_202_in0), .in1(eq_202_in1), .out(eq_202_out));

	wire [31:0] eq_203_in0;
	wire [31:0] eq_203_in1;
	wire [0:0] eq_203_out;
	eq #(.WIDTH(32)) eq_203(.in0(eq_203_in0), .in1(eq_203_in1), .out(eq_203_out));

	wire [31:0] eq_204_in0;
	wire [31:0] eq_204_in1;
	wire [0:0] eq_204_out;
	eq #(.WIDTH(32)) eq_204(.in0(eq_204_in0), .in1(eq_204_in1), .out(eq_204_out));

	wire [0:0] andOp_205_in0;
	wire [0:0] andOp_205_in1;
	wire [0:0] andOp_205_out;
	andOp #(.WIDTH(1)) andOp_205(.in0(andOp_205_in0), .in1(andOp_205_in1), .out(andOp_205_out));

	wire [0:0] andOp_206_in0;
	wire [0:0] andOp_206_in1;
	wire [0:0] andOp_206_out;
	andOp #(.WIDTH(1)) andOp_206(.in0(andOp_206_in0), .in1(andOp_206_in1), .out(andOp_206_out));

	wire [0:0] andOp_207_in0;
	wire [0:0] andOp_207_in1;
	wire [0:0] andOp_207_out;
	andOp #(.WIDTH(1)) andOp_207(.in0(andOp_207_in0), .in1(andOp_207_in1), .out(andOp_207_out));

	wire [0:0] andOp_208_in0;
	wire [0:0] andOp_208_in1;
	wire [0:0] andOp_208_out;
	andOp #(.WIDTH(1)) andOp_208(.in0(andOp_208_in0), .in1(andOp_208_in1), .out(andOp_208_out));

	wire [0:0] andOp_209_in0;
	wire [0:0] andOp_209_in1;
	wire [0:0] andOp_209_out;
	andOp #(.WIDTH(1)) andOp_209(.in0(andOp_209_in0), .in1(andOp_209_in1), .out(andOp_209_out));

	wire [0:0] andOp_210_in0;
	wire [0:0] andOp_210_in1;
	wire [0:0] andOp_210_out;
	andOp #(.WIDTH(1)) andOp_210(.in0(andOp_210_in0), .in1(andOp_210_in1), .out(andOp_210_out));

	wire [31:0] eq_211_in0;
	wire [31:0] eq_211_in1;
	wire [0:0] eq_211_out;
	eq #(.WIDTH(32)) eq_211(.in0(eq_211_in0), .in1(eq_211_in1), .out(eq_211_out));

	wire [31:0] eq_212_in0;
	wire [31:0] eq_212_in1;
	wire [0:0] eq_212_out;
	eq #(.WIDTH(32)) eq_212(.in0(eq_212_in0), .in1(eq_212_in1), .out(eq_212_out));

	wire [0:0] andOp_213_in0;
	wire [0:0] andOp_213_in1;
	wire [0:0] andOp_213_out;
	andOp #(.WIDTH(1)) andOp_213(.in0(andOp_213_in0), .in1(andOp_213_in1), .out(andOp_213_out));

	wire [31:0] eq_214_in0;
	wire [31:0] eq_214_in1;
	wire [0:0] eq_214_out;
	eq #(.WIDTH(32)) eq_214(.in0(eq_214_in0), .in1(eq_214_in1), .out(eq_214_out));

	wire [31:0] eq_215_in0;
	wire [31:0] eq_215_in1;
	wire [0:0] eq_215_out;
	eq #(.WIDTH(32)) eq_215(.in0(eq_215_in0), .in1(eq_215_in1), .out(eq_215_out));

	wire [0:0] andOp_216_in0;
	wire [0:0] andOp_216_in1;
	wire [0:0] andOp_216_out;
	andOp #(.WIDTH(1)) andOp_216(.in0(andOp_216_in0), .in1(andOp_216_in1), .out(andOp_216_out));

	wire [31:0] eq_217_in0;
	wire [31:0] eq_217_in1;
	wire [0:0] eq_217_out;
	eq #(.WIDTH(32)) eq_217(.in0(eq_217_in0), .in1(eq_217_in1), .out(eq_217_out));

	wire [31:0] eq_218_in0;
	wire [31:0] eq_218_in1;
	wire [0:0] eq_218_out;
	eq #(.WIDTH(32)) eq_218(.in0(eq_218_in0), .in1(eq_218_in1), .out(eq_218_out));

	wire [0:0] andOp_219_in0;
	wire [0:0] andOp_219_in1;
	wire [0:0] andOp_219_out;
	andOp #(.WIDTH(1)) andOp_219(.in0(andOp_219_in0), .in1(andOp_219_in1), .out(andOp_219_out));

	wire [0:0] andOp_220_in0;
	wire [0:0] andOp_220_in1;
	wire [0:0] andOp_220_out;
	andOp #(.WIDTH(1)) andOp_220(.in0(andOp_220_in0), .in1(andOp_220_in1), .out(andOp_220_out));

	wire [31:0] eq_221_in0;
	wire [31:0] eq_221_in1;
	wire [0:0] eq_221_out;
	eq #(.WIDTH(32)) eq_221(.in0(eq_221_in0), .in1(eq_221_in1), .out(eq_221_out));

	wire [31:0] eq_222_in0;
	wire [31:0] eq_222_in1;
	wire [0:0] eq_222_out;
	eq #(.WIDTH(32)) eq_222(.in0(eq_222_in0), .in1(eq_222_in1), .out(eq_222_out));

	wire [31:0] eq_223_in0;
	wire [31:0] eq_223_in1;
	wire [0:0] eq_223_out;
	eq #(.WIDTH(32)) eq_223(.in0(eq_223_in0), .in1(eq_223_in1), .out(eq_223_out));

	wire [31:0] eq_224_in0;
	wire [31:0] eq_224_in1;
	wire [0:0] eq_224_out;
	eq #(.WIDTH(32)) eq_224(.in0(eq_224_in0), .in1(eq_224_in1), .out(eq_224_out));

	wire [31:0] eq_225_in0;
	wire [31:0] eq_225_in1;
	wire [0:0] eq_225_out;
	eq #(.WIDTH(32)) eq_225(.in0(eq_225_in0), .in1(eq_225_in1), .out(eq_225_out));

	wire [31:0] eq_226_in0;
	wire [31:0] eq_226_in1;
	wire [0:0] eq_226_out;
	eq #(.WIDTH(32)) eq_226(.in0(eq_226_in0), .in1(eq_226_in1), .out(eq_226_out));

	// End Functional Units

	reg [31:0] data_store_0_0;
	reg [31:0] data_store_0_10;
	reg [31:0] data_store_0_11;
	reg [31:0] data_store_0_3;
	reg [0:0] data_store_0_5;
	reg [31:0] data_store_0_6;
	reg [31:0] data_store_0_8;
	reg [31:0] data_store_1_12;
	reg [31:0] data_store_1_13;
	reg [31:0] data_store_1_15;
	reg [0:0] data_store_1_17;
	reg [31:0] data_store_1_19;
	reg [31:0] data_store_1_21;
	reg [31:0] data_store_1_24;
	reg [31:0] data_store_2_27;
	reg [31:0] data_store_2_29;
	reg [31:0] data_store_2_30;
	reg [31:0] data_store_2_33;
	reg [31:0] data_store_2_35;
	reg [31:0] data_store_3_38;
	reg [31:0] data_store_3_40;
	reg [31:0] data_store_3_42;
	reg [31:0] data_store_3_44;
	reg [31:0] data_store_3_46;
	reg [0:0] data_store_3_47;
	reg [31:0] data_store_4_48;
	reg [31:0] data_store_4_50;
	reg [31:0] data_store_4_52;
	reg [31:0] data_store_4_54;
	reg [31:0] data_store_4_56;
	reg [0:0] data_store_4_58;
	reg [31:0] data_store_5_60;
	reg [31:0] data_store_5_62;
	reg [31:0] data_store_5_64;
	reg [31:0] data_store_5_66;
	reg [31:0] data_store_5_68;
	reg [0:0] data_store_5_70;
	reg [31:0] data_store_6_72;
	reg [31:0] data_store_6_74;
	reg [31:0] data_store_6_76;
	reg [31:0] data_store_6_78;
	reg [31:0] data_store_6_80;
	reg [31:0] global_state;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_3_last_state;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;
	reg [31:0] state_4_last_state;
	reg [31:0] state_5_entry_BB_reg;
	reg [0:0] state_5_is_active;
	reg [31:0] state_5_last_BB_reg;
	reg [31:0] state_5_last_state;
	reg [31:0] state_6_entry_BB_reg;
	reg [0:0] state_6_is_active;
	reg [31:0] state_6_last_BB_reg;
	reg [31:0] state_6_last_state;

	// controller for add_add12.add_add12_in0
	// controller for add_add12.add_add12_in1
	// Insensitive connections
	assign add_add12_in0 = data_in_1_23_out_data;
	assign add_add12_in1 = data_in_1_20_out_data;
	// controller for add_add13.add_add13_in0
	// controller for add_add13.add_add13_in1
	// Insensitive connections
	assign add_add13_in0 = mul_mul16_out;
	assign add_add13_in1 = data_in_2_37_out_data;
	// controller for add_add20.add_add20_in0
	// controller for add_add20.add_add20_in1
	// Insensitive connections
	assign add_add20_in0 = data_in_3_39_out_data;
	assign add_add20_in1 = 32'd12;
	// controller for add_add21.add_add21_in0
	// controller for add_add21.add_add21_in1
	// Insensitive connections
	assign add_add21_in0 = data_in_3_39_out_data;
	assign add_add21_in1 = 32'd1;
	// controller for add_add3.add_add3_in0
	// controller for add_add3.add_add3_in1
	// Insensitive connections
	assign add_add3_in0 = phi_phi6_out;
	assign add_add3_in1 = 32'd1;
	// controller for add_add7.add_add7_in0
	// controller for add_add7.add_add7_in1
	// Insensitive connections
	assign add_add7_in0 = phi_phi6_out;
	assign add_add7_in1 = 32'd9;
	// controller for andOp_101.andOp_101_in0
	// controller for andOp_101.andOp_101_in1
	// Insensitive connections
	assign andOp_101_in0 = andOp_97_out;
	assign andOp_101_in1 = notOp_100_out;
	// controller for andOp_102.andOp_102_in0
	// controller for andOp_102.andOp_102_in1
	// Insensitive connections
	assign andOp_102_in0 = bb_3_active_in_state_6_out_data;
	assign andOp_102_in1 = state_6_is_active;
	// controller for andOp_104.andOp_104_in0
	// controller for andOp_104.andOp_104_in1
	// Insensitive connections
	assign andOp_104_in0 = andOp_102_out;
	assign andOp_104_in1 = data_in_6_82_out_data;
	// controller for andOp_106.andOp_106_in0
	// controller for andOp_106.andOp_106_in1
	// Insensitive connections
	assign andOp_106_in0 = andOp_102_out;
	assign andOp_106_in1 = notOp_105_out;
	// controller for andOp_107.andOp_107_in0
	// controller for andOp_107.andOp_107_in1
	// Insensitive connections
	assign andOp_107_in0 = bb_3_active_in_state_6_out_data;
	assign andOp_107_in1 = state_6_is_active;
	// controller for andOp_109.andOp_109_in0
	// controller for andOp_109.andOp_109_in1
	// Insensitive connections
	assign andOp_109_in0 = andOp_107_out;
	assign andOp_109_in1 = data_in_6_82_out_data;
	// controller for andOp_111.andOp_111_in0
	// controller for andOp_111.andOp_111_in1
	// Insensitive connections
	assign andOp_111_in0 = andOp_107_out;
	assign andOp_111_in1 = notOp_110_out;
	// controller for andOp_112.andOp_112_in0
	// controller for andOp_112.andOp_112_in1
	// Insensitive connections
	assign andOp_112_in0 = bb_3_active_in_state_6_out_data;
	assign andOp_112_in1 = state_6_is_active;
	// controller for andOp_114.andOp_114_in0
	// controller for andOp_114.andOp_114_in1
	// Insensitive connections
	assign andOp_114_in0 = andOp_112_out;
	assign andOp_114_in1 = data_in_6_82_out_data;
	// controller for andOp_116.andOp_116_in0
	// controller for andOp_116.andOp_116_in1
	// Insensitive connections
	assign andOp_116_in0 = andOp_112_out;
	assign andOp_116_in1 = notOp_115_out;
	// controller for andOp_117.andOp_117_in0
	// controller for andOp_117.andOp_117_in1
	// Insensitive connections
	assign andOp_117_in0 = bb_3_active_in_state_6_out_data;
	assign andOp_117_in1 = state_6_is_active;
	// controller for andOp_119.andOp_119_in0
	// controller for andOp_119.andOp_119_in1
	// Insensitive connections
	assign andOp_119_in0 = andOp_117_out;
	assign andOp_119_in1 = data_in_6_82_out_data;
	// controller for andOp_121.andOp_121_in0
	// controller for andOp_121.andOp_121_in1
	// Insensitive connections
	assign andOp_121_in0 = andOp_117_out;
	assign andOp_121_in1 = notOp_120_out;
	// controller for andOp_138.andOp_138_in0
	// controller for andOp_138.andOp_138_in1
	// Insensitive connections
	assign andOp_138_in0 = notOp_137_out;
	assign andOp_138_in1 = andOp_83_out;
	// controller for andOp_141.andOp_141_in0
	// controller for andOp_141.andOp_141_in1
	// Insensitive connections
	assign andOp_141_in0 = notOp_140_out;
	assign andOp_141_in1 = andOp_85_out;
	// controller for andOp_150.andOp_150_in0
	// controller for andOp_150.andOp_150_in1
	// Insensitive connections
	assign andOp_150_in0 = notOp_149_out;
	assign andOp_150_in1 = andOp_104_out;
	// controller for andOp_151.andOp_151_in0
	// controller for andOp_151.andOp_151_in1
	// Insensitive connections
	assign andOp_151_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_151_in1 = state_0_is_active;
	// controller for andOp_152.andOp_152_in0
	// controller for andOp_152.andOp_152_in1
	// Insensitive connections
	assign andOp_152_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_152_in1 = state_1_is_active;
	// controller for andOp_153.andOp_153_in0
	// controller for andOp_153.andOp_153_in1
	// Insensitive connections
	assign andOp_153_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_153_in1 = state_1_is_active;
	// controller for andOp_154.andOp_154_in0
	// controller for andOp_154.andOp_154_in1
	// Insensitive connections
	assign andOp_154_in0 = bb_4_active_in_state_2_out_data;
	assign andOp_154_in1 = state_2_is_active;
	// controller for andOp_155.andOp_155_in0
	// controller for andOp_155.andOp_155_in1
	// Insensitive connections
	assign andOp_155_in0 = bb_3_active_in_state_3_out_data;
	assign andOp_155_in1 = state_3_is_active;
	// controller for andOp_156.andOp_156_in0
	// controller for andOp_156.andOp_156_in1
	// Insensitive connections
	assign andOp_156_in0 = bb_3_active_in_state_3_out_data;
	assign andOp_156_in1 = state_3_is_active;
	// controller for andOp_157.andOp_157_in0
	// controller for andOp_157.andOp_157_in1
	// Insensitive connections
	assign andOp_157_in0 = bb_3_active_in_state_3_out_data;
	assign andOp_157_in1 = state_3_is_active;
	// controller for andOp_158.andOp_158_in0
	// controller for andOp_158.andOp_158_in1
	// Insensitive connections
	assign andOp_158_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_158_in1 = state_0_is_active;
	// controller for andOp_161.andOp_161_in0
	// controller for andOp_161.andOp_161_in1
	// Insensitive connections
	assign andOp_161_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_161_in1 = state_0_is_active;
	// controller for andOp_162.andOp_162_in0
	// controller for andOp_162.andOp_162_in1
	// Insensitive connections
	assign andOp_162_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_162_in1 = state_0_is_active;
	// controller for andOp_163.andOp_163_in0
	// controller for andOp_163.andOp_163_in1
	// Insensitive connections
	assign andOp_163_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_163_in1 = state_0_is_active;
	// controller for andOp_164.andOp_164_in0
	// controller for andOp_164.andOp_164_in1
	// Insensitive connections
	assign andOp_164_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_164_in1 = state_0_is_active;
	// controller for andOp_167.andOp_167_in0
	// controller for andOp_167.andOp_167_in1
	// Insensitive connections
	assign andOp_167_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_167_in1 = state_0_is_active;
	// controller for andOp_168.andOp_168_in0
	// controller for andOp_168.andOp_168_in1
	// Insensitive connections
	assign andOp_168_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_168_in1 = state_0_is_active;
	// controller for andOp_171.andOp_171_in0
	// controller for andOp_171.andOp_171_in1
	// Insensitive connections
	assign andOp_171_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_171_in1 = state_1_is_active;
	// controller for andOp_172.andOp_172_in0
	// controller for andOp_172.andOp_172_in1
	// Insensitive connections
	assign andOp_172_in0 = bb_4_active_in_state_2_out_data;
	assign andOp_172_in1 = state_2_is_active;
	// controller for andOp_173.andOp_173_in0
	// controller for andOp_173.andOp_173_in1
	// Insensitive connections
	assign andOp_173_in0 = bb_4_active_in_state_2_out_data;
	assign andOp_173_in1 = state_2_is_active;
	// controller for andOp_174.andOp_174_in0
	// controller for andOp_174.andOp_174_in1
	// Insensitive connections
	assign andOp_174_in0 = bb_3_active_in_state_3_out_data;
	assign andOp_174_in1 = state_3_is_active;
	// controller for andOp_175.andOp_175_in0
	// controller for andOp_175.andOp_175_in1
	// Insensitive connections
	assign andOp_175_in0 = bb_3_active_in_state_3_out_data;
	assign andOp_175_in1 = state_3_is_active;
	// controller for andOp_176.andOp_176_in0
	// controller for andOp_176.andOp_176_in1
	// Insensitive connections
	assign andOp_176_in0 = bb_3_active_in_state_3_out_data;
	assign andOp_176_in1 = state_3_is_active;
	// controller for andOp_177.andOp_177_in0
	// controller for andOp_177.andOp_177_in1
	// Insensitive connections
	assign andOp_177_in0 = bb_2_active_in_state_6_out_data;
	assign andOp_177_in1 = state_6_is_active;
	// controller for andOp_178.andOp_178_in0
	// controller for andOp_178.andOp_178_in1
	// Insensitive connections
	assign andOp_178_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_178_in1 = state_0_is_active;
	// controller for andOp_179.andOp_179_in0
	// controller for andOp_179.andOp_179_in1
	// Insensitive connections
	assign andOp_179_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_179_in1 = state_1_is_active;
	// controller for andOp_180.andOp_180_in0
	// controller for andOp_180.andOp_180_in1
	// Insensitive connections
	assign andOp_180_in0 = bb_3_active_in_state_3_out_data;
	assign andOp_180_in1 = state_3_is_active;
	// controller for andOp_181.andOp_181_in0
	// controller for andOp_181.andOp_181_in1
	// Insensitive connections
	assign andOp_181_in0 = bb_3_active_in_state_4_out_data;
	assign andOp_181_in1 = state_4_is_active;
	// controller for andOp_182.andOp_182_in0
	// controller for andOp_182.andOp_182_in1
	// Insensitive connections
	assign andOp_182_in0 = bb_3_active_in_state_5_out_data;
	assign andOp_182_in1 = state_5_is_active;
	// controller for andOp_183.andOp_183_in0
	// controller for andOp_183.andOp_183_in1
	// Insensitive connections
	assign andOp_183_in0 = bb_2_active_in_state_6_out_data;
	assign andOp_183_in1 = state_6_is_active;
	// controller for andOp_185.andOp_185_in0
	// controller for andOp_185.andOp_185_in1
	// Insensitive connections
	assign andOp_185_in0 = notOp_184_out;
	assign andOp_185_in1 = 1'd1;
	// controller for andOp_187.andOp_187_in0
	// controller for andOp_187.andOp_187_in1
	// Insensitive connections
	assign andOp_187_in0 = notOp_186_out;
	assign andOp_187_in1 = andOp_185_out;
	// controller for andOp_189.andOp_189_in0
	// controller for andOp_189.andOp_189_in1
	// Insensitive connections
	assign andOp_189_in0 = notOp_188_out;
	assign andOp_189_in1 = 1'd1;
	// controller for andOp_191.andOp_191_in0
	// controller for andOp_191.andOp_191_in1
	// Insensitive connections
	assign andOp_191_in0 = notOp_190_out;
	assign andOp_191_in1 = 1'd1;
	// controller for andOp_193.andOp_193_in0
	// controller for andOp_193.andOp_193_in1
	// Insensitive connections
	assign andOp_193_in0 = notOp_192_out;
	assign andOp_193_in1 = 1'd1;
	// controller for andOp_195.andOp_195_in0
	// controller for andOp_195.andOp_195_in1
	// Insensitive connections
	assign andOp_195_in0 = notOp_194_out;
	assign andOp_195_in1 = 1'd1;
	// controller for andOp_197.andOp_197_in0
	// controller for andOp_197.andOp_197_in1
	// Insensitive connections
	assign andOp_197_in0 = notOp_196_out;
	assign andOp_197_in1 = 1'd1;
	// controller for andOp_199.andOp_199_in0
	// controller for andOp_199.andOp_199_in1
	// Insensitive connections
	assign andOp_199_in0 = notOp_198_out;
	assign andOp_199_in1 = 1'd1;
	// controller for andOp_201.andOp_201_in0
	// controller for andOp_201.andOp_201_in1
	// Insensitive connections
	assign andOp_201_in0 = notOp_200_out;
	assign andOp_201_in1 = andOp_199_out;
	// controller for andOp_205.andOp_205_in0
	// controller for andOp_205.andOp_205_in1
	// Insensitive connections
	assign andOp_205_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_205_in1 = state_0_is_active;
	// controller for andOp_206.andOp_206_in0
	// controller for andOp_206.andOp_206_in1
	// Insensitive connections
	assign andOp_206_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_206_in1 = state_0_is_active;
	// controller for andOp_207.andOp_207_in0
	// controller for andOp_207.andOp_207_in1
	// Insensitive connections
	assign andOp_207_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_207_in1 = state_0_is_active;
	// controller for andOp_208.andOp_208_in0
	// controller for andOp_208.andOp_208_in1
	// Insensitive connections
	assign andOp_208_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_208_in1 = state_0_is_active;
	// controller for andOp_209.andOp_209_in0
	// controller for andOp_209.andOp_209_in1
	// Insensitive connections
	assign andOp_209_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_209_in1 = state_0_is_active;
	// controller for andOp_210.andOp_210_in0
	// controller for andOp_210.andOp_210_in1
	// Insensitive connections
	assign andOp_210_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_210_in1 = state_0_is_active;
	// controller for andOp_213.andOp_213_in0
	// controller for andOp_213.andOp_213_in1
	// Insensitive connections
	assign andOp_213_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_213_in1 = state_1_is_active;
	// controller for andOp_216.andOp_216_in0
	// controller for andOp_216.andOp_216_in1
	// Insensitive connections
	assign andOp_216_in0 = bb_4_active_in_state_2_out_data;
	assign andOp_216_in1 = state_2_is_active;
	// controller for andOp_219.andOp_219_in0
	// controller for andOp_219.andOp_219_in1
	// Insensitive connections
	assign andOp_219_in0 = bb_3_active_in_state_3_out_data;
	assign andOp_219_in1 = state_3_is_active;
	// controller for andOp_220.andOp_220_in0
	// controller for andOp_220.andOp_220_in1
	// Insensitive connections
	assign andOp_220_in0 = bb_3_active_in_state_3_out_data;
	assign andOp_220_in1 = state_3_is_active;
	// controller for andOp_83.andOp_83_in0
	// controller for andOp_83.andOp_83_in1
	// Insensitive connections
	assign andOp_83_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_83_in1 = state_0_is_active;
	// controller for andOp_85.andOp_85_in0
	// controller for andOp_85.andOp_85_in1
	// Insensitive connections
	assign andOp_85_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_85_in1 = state_0_is_active;
	// controller for andOp_87.andOp_87_in0
	// controller for andOp_87.andOp_87_in1
	// Insensitive connections
	assign andOp_87_in0 = bb_4_active_in_state_2_out_data;
	assign andOp_87_in1 = state_2_is_active;
	// controller for andOp_89.andOp_89_in0
	// controller for andOp_89.andOp_89_in1
	// Insensitive connections
	assign andOp_89_in0 = andOp_87_out;
	assign andOp_89_in1 = data_in_2_32_out_data;
	// controller for andOp_91.andOp_91_in0
	// controller for andOp_91.andOp_91_in1
	// Insensitive connections
	assign andOp_91_in0 = andOp_87_out;
	assign andOp_91_in1 = notOp_90_out;
	// controller for andOp_92.andOp_92_in0
	// controller for andOp_92.andOp_92_in1
	// Insensitive connections
	assign andOp_92_in0 = bb_4_active_in_state_2_out_data;
	assign andOp_92_in1 = state_2_is_active;
	// controller for andOp_94.andOp_94_in0
	// controller for andOp_94.andOp_94_in1
	// Insensitive connections
	assign andOp_94_in0 = andOp_92_out;
	assign andOp_94_in1 = data_in_2_32_out_data;
	// controller for andOp_96.andOp_96_in0
	// controller for andOp_96.andOp_96_in1
	// Insensitive connections
	assign andOp_96_in0 = andOp_92_out;
	assign andOp_96_in1 = notOp_95_out;
	// controller for andOp_97.andOp_97_in0
	// controller for andOp_97.andOp_97_in1
	// Insensitive connections
	assign andOp_97_in0 = bb_4_active_in_state_2_out_data;
	assign andOp_97_in1 = state_2_is_active;
	// controller for andOp_99.andOp_99_in0
	// controller for andOp_99.andOp_99_in1
	// Insensitive connections
	assign andOp_99_in0 = andOp_97_out;
	assign andOp_99_in1 = data_in_2_32_out_data;
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_122_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_135_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_0.bb_1_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_0_in_data = orOp_124_out;
		end else begin
			bb_1_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_0.bb_1_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_138_out) begin 
			bb_1_predecessor_in_state_0_in_data = 32'd0;
		end else if (eq_136_out) begin 
			bb_1_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_6.bb_2_active_in_state_6_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_6_in_data = orOp_134_out;
		end else begin
			bb_2_active_in_state_6_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_6.bb_2_predecessor_in_state_6_in_data
	always @(*) begin
		if (andOp_150_out) begin 
			bb_2_predecessor_in_state_6_in_data = 32'd3;
		end else if (eq_148_out) begin 
			bb_2_predecessor_in_state_6_in_data = state_6_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_6_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_3.bb_3_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_3_in_data = eq_129_out;
		end else begin
			bb_3_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_4.bb_3_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_4_in_data = eq_130_out;
		end else begin
			bb_3_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_5.bb_3_active_in_state_5_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_5_in_data = eq_131_out;
		end else begin
			bb_3_active_in_state_5_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_6.bb_3_active_in_state_6_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_6_in_data = eq_132_out;
		end else begin
			bb_3_active_in_state_6_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_3.bb_3_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_144_out) begin 
			bb_3_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_4.bb_3_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_145_out) begin 
			bb_3_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_5.bb_3_predecessor_in_state_5_in_data
	always @(*) begin
		if (eq_146_out) begin 
			bb_3_predecessor_in_state_5_in_data = state_5_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_5_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_6.bb_3_predecessor_in_state_6_in_data
	always @(*) begin
		if (eq_147_out) begin 
			bb_3_predecessor_in_state_6_in_data = state_6_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_6_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_0.bb_4_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_0_in_data = orOp_126_out;
		end else begin
			bb_4_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_1.bb_4_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_1_in_data = eq_127_out;
		end else begin
			bb_4_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_2.bb_4_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_2_in_data = eq_128_out;
		end else begin
			bb_4_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_0.bb_4_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_141_out) begin 
			bb_4_predecessor_in_state_0_in_data = 32'd1;
		end else if (eq_139_out) begin 
			bb_4_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_1.bb_4_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_142_out) begin 
			bb_4_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_2.bb_4_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_143_out) begin 
			bb_4_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_83_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_84_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_1_happened_in_state_0.br_1_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_85_out) begin 
			br_1_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_86_out) begin 
			br_1_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_1_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_3.br_3_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_102_out) begin 
			br_3_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_103_out) begin 
			br_3_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_4.br_3_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_107_out) begin 
			br_3_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_108_out) begin 
			br_3_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_5.br_3_happened_in_state_5_in_data
	always @(*) begin
		if (andOp_112_out) begin 
			br_3_happened_in_state_5_in_data = 1'd1;
		end else if (notOp_113_out) begin 
			br_3_happened_in_state_5_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_5_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_6.br_3_happened_in_state_6_in_data
	always @(*) begin
		if (andOp_117_out) begin 
			br_3_happened_in_state_6_in_data = 1'd1;
		end else if (notOp_118_out) begin 
			br_3_happened_in_state_6_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_6_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_0.br_4_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_87_out) begin 
			br_4_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_88_out) begin 
			br_4_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_1.br_4_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_92_out) begin 
			br_4_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_93_out) begin 
			br_4_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_2.br_4_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_97_out) begin 
			br_4_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_98_out) begin 
			br_4_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_2_in_data = 0;
		end
	end
	// controller for concat_159.concat_159_in0
	// controller for concat_159.concat_159_in1
	// Insensitive connections
	assign concat_159_in0 = data_in_0_9_out_data;
	assign concat_159_in1 = 32'd0;
	// controller for concat_160.concat_160_in0
	// controller for concat_160.concat_160_in1
	// Insensitive connections
	assign concat_160_in0 = 32'd3;
	assign concat_160_in1 = 32'd0;
	// controller for concat_165.concat_165_in0
	// controller for concat_165.concat_165_in1
	// Insensitive connections
	assign concat_165_in0 = data_in_0_4_out_data;
	assign concat_165_in1 = 32'd0;
	// controller for concat_166.concat_166_in0
	// controller for concat_166.concat_166_in1
	// Insensitive connections
	assign concat_166_in0 = 32'd4;
	assign concat_166_in1 = 32'd1;
	// controller for concat_169.concat_169_in0
	// controller for concat_169.concat_169_in1
	// Insensitive connections
	assign concat_169_in0 = data_in_0_2_out_data;
	assign concat_169_in1 = 32'd0;
	// controller for concat_170.concat_170_in0
	// controller for concat_170.concat_170_in1
	// Insensitive connections
	assign concat_170_in0 = 32'd4;
	assign concat_170_in1 = 32'd1;
	// controller for data_in_0_1.data_in_0_1_in_data
	always @(*) begin
		if (eq_202_out) begin 
			data_in_0_1_in_data = data_store_0_0;
		end else if (eq_203_out) begin 
			data_in_0_1_in_data = data_store_2_27;
		end else if (eq_204_out) begin 
			data_in_0_1_in_data = data_store_6_72;
		end else begin
			data_in_0_1_in_data = 0;
		end
	end
	// controller for data_in_0_2.data_in_0_2_in_data
	always @(*) begin
		if (eq_202_out) begin 
			data_in_0_2_in_data = 32'd0;
		end else if (eq_203_out) begin 
			data_in_0_2_in_data = data_store_2_29;
		end else if (eq_204_out) begin 
			data_in_0_2_in_data = data_store_6_74;
		end else begin
			data_in_0_2_in_data = 0;
		end
	end
	// controller for data_in_0_4.data_in_0_4_in_data
	always @(*) begin
		if (eq_202_out) begin 
			data_in_0_4_in_data = data_store_0_3;
		end else if (eq_203_out) begin 
			data_in_0_4_in_data = data_store_2_30;
		end else if (eq_204_out) begin 
			data_in_0_4_in_data = data_store_6_76;
		end else begin
			data_in_0_4_in_data = 0;
		end
	end
	// controller for data_in_0_7.data_in_0_7_in_data
	always @(*) begin
		if (eq_202_out) begin 
			data_in_0_7_in_data = data_store_0_6;
		end else if (eq_203_out) begin 
			data_in_0_7_in_data = data_store_2_33;
		end else if (eq_204_out) begin 
			data_in_0_7_in_data = data_store_6_78;
		end else begin
			data_in_0_7_in_data = 0;
		end
	end
	// controller for data_in_0_9.data_in_0_9_in_data
	always @(*) begin
		if (eq_202_out) begin 
			data_in_0_9_in_data = data_store_0_8;
		end else if (eq_203_out) begin 
			data_in_0_9_in_data = data_store_2_35;
		end else if (eq_204_out) begin 
			data_in_0_9_in_data = data_store_6_80;
		end else begin
			data_in_0_9_in_data = 0;
		end
	end
	// controller for data_in_1_14.data_in_1_14_in_data
	always @(*) begin
		if (eq_211_out) begin 
			data_in_1_14_in_data = data_store_0_0;
		end else if (eq_212_out) begin 
			data_in_1_14_in_data = data_store_1_13;
		end else begin
			data_in_1_14_in_data = 0;
		end
	end
	// controller for data_in_1_16.data_in_1_16_in_data
	always @(*) begin
		if (eq_211_out) begin 
			data_in_1_16_in_data = data_store_0_3;
		end else if (eq_212_out) begin 
			data_in_1_16_in_data = data_store_1_15;
		end else begin
			data_in_1_16_in_data = 0;
		end
	end
	// controller for data_in_1_18.data_in_1_18_in_data
	always @(*) begin
		if (eq_211_out) begin 
			data_in_1_18_in_data = data_store_0_5;
		end else if (eq_212_out) begin 
			data_in_1_18_in_data = data_store_1_17;
		end else begin
			data_in_1_18_in_data = 0;
		end
	end
	// controller for data_in_1_20.data_in_1_20_in_data
	always @(*) begin
		if (eq_211_out) begin 
			data_in_1_20_in_data = data_store_0_6;
		end else if (eq_212_out) begin 
			data_in_1_20_in_data = data_store_1_19;
		end else begin
			data_in_1_20_in_data = 0;
		end
	end
	// controller for data_in_1_22.data_in_1_22_in_data
	always @(*) begin
		if (eq_211_out) begin 
			data_in_1_22_in_data = data_store_0_8;
		end else if (eq_212_out) begin 
			data_in_1_22_in_data = data_store_1_21;
		end else begin
			data_in_1_22_in_data = 0;
		end
	end
	// controller for data_in_1_23.data_in_1_23_in_data
	always @(*) begin
		if (eq_211_out) begin 
			data_in_1_23_in_data = data_store_0_10;
		end else if (eq_212_out) begin 
			data_in_1_23_in_data = 32'd0;
		end else begin
			data_in_1_23_in_data = 0;
		end
	end
	// controller for data_in_1_25.data_in_1_25_in_data
	always @(*) begin
		if (eq_211_out) begin 
			data_in_1_25_in_data = data_store_0_11;
		end else if (eq_212_out) begin 
			data_in_1_25_in_data = data_store_1_24;
		end else begin
			data_in_1_25_in_data = 0;
		end
	end
	// controller for data_in_2_26.data_in_2_26_in_data
	always @(*) begin
		if (eq_214_out) begin 
			data_in_2_26_in_data = data_store_1_12;
		end else if (eq_215_out) begin 
			data_in_2_26_in_data = 32'd0;
		end else begin
			data_in_2_26_in_data = 0;
		end
	end
	// controller for data_in_2_28.data_in_2_28_in_data
	always @(*) begin
		if (eq_214_out) begin 
			data_in_2_28_in_data = data_store_1_13;
		end else if (eq_215_out) begin 
			data_in_2_28_in_data = data_store_2_27;
		end else begin
			data_in_2_28_in_data = 0;
		end
	end
	// controller for data_in_2_31.data_in_2_31_in_data
	always @(*) begin
		if (eq_214_out) begin 
			data_in_2_31_in_data = data_store_1_15;
		end else if (eq_215_out) begin 
			data_in_2_31_in_data = data_store_2_30;
		end else begin
			data_in_2_31_in_data = 0;
		end
	end
	// controller for data_in_2_32.data_in_2_32_in_data
	always @(*) begin
		if (eq_214_out) begin 
			data_in_2_32_in_data = data_store_1_17;
		end else if (eq_215_out) begin 
			data_in_2_32_in_data = 1'd0;
		end else begin
			data_in_2_32_in_data = 0;
		end
	end
	// controller for data_in_2_34.data_in_2_34_in_data
	always @(*) begin
		if (eq_214_out) begin 
			data_in_2_34_in_data = data_store_1_19;
		end else if (eq_215_out) begin 
			data_in_2_34_in_data = data_store_2_33;
		end else begin
			data_in_2_34_in_data = 0;
		end
	end
	// controller for data_in_2_36.data_in_2_36_in_data
	always @(*) begin
		if (eq_214_out) begin 
			data_in_2_36_in_data = data_store_1_21;
		end else if (eq_215_out) begin 
			data_in_2_36_in_data = data_store_2_35;
		end else begin
			data_in_2_36_in_data = 0;
		end
	end
	// controller for data_in_2_37.data_in_2_37_in_data
	always @(*) begin
		if (eq_214_out) begin 
			data_in_2_37_in_data = data_store_1_24;
		end else if (eq_215_out) begin 
			data_in_2_37_in_data = 32'd0;
		end else begin
			data_in_2_37_in_data = 0;
		end
	end
	// controller for data_in_3_39.data_in_3_39_in_data
	always @(*) begin
		if (eq_217_out) begin 
			data_in_3_39_in_data = data_store_2_27;
		end else if (eq_218_out) begin 
			data_in_3_39_in_data = data_store_3_38;
		end else begin
			data_in_3_39_in_data = 0;
		end
	end
	// controller for data_in_3_41.data_in_3_41_in_data
	always @(*) begin
		if (eq_217_out) begin 
			data_in_3_41_in_data = data_store_2_29;
		end else if (eq_218_out) begin 
			data_in_3_41_in_data = data_store_3_40;
		end else begin
			data_in_3_41_in_data = 0;
		end
	end
	// controller for data_in_3_43.data_in_3_43_in_data
	always @(*) begin
		if (eq_217_out) begin 
			data_in_3_43_in_data = data_store_2_30;
		end else if (eq_218_out) begin 
			data_in_3_43_in_data = data_store_3_42;
		end else begin
			data_in_3_43_in_data = 0;
		end
	end
	// controller for data_in_3_45.data_in_3_45_in_data
	always @(*) begin
		if (eq_217_out) begin 
			data_in_3_45_in_data = data_store_2_33;
		end else if (eq_218_out) begin 
			data_in_3_45_in_data = data_store_3_44;
		end else begin
			data_in_3_45_in_data = 0;
		end
	end
	// controller for data_in_4_49.data_in_4_49_in_data
	always @(*) begin
		if (eq_221_out) begin 
			data_in_4_49_in_data = data_store_3_38;
		end else if (eq_222_out) begin 
			data_in_4_49_in_data = data_store_4_48;
		end else begin
			data_in_4_49_in_data = 0;
		end
	end
	// controller for data_in_4_51.data_in_4_51_in_data
	always @(*) begin
		if (eq_221_out) begin 
			data_in_4_51_in_data = data_store_3_40;
		end else if (eq_222_out) begin 
			data_in_4_51_in_data = data_store_4_50;
		end else begin
			data_in_4_51_in_data = 0;
		end
	end
	// controller for data_in_4_53.data_in_4_53_in_data
	always @(*) begin
		if (eq_221_out) begin 
			data_in_4_53_in_data = data_store_3_42;
		end else if (eq_222_out) begin 
			data_in_4_53_in_data = data_store_4_52;
		end else begin
			data_in_4_53_in_data = 0;
		end
	end
	// controller for data_in_4_55.data_in_4_55_in_data
	always @(*) begin
		if (eq_221_out) begin 
			data_in_4_55_in_data = data_store_3_44;
		end else if (eq_222_out) begin 
			data_in_4_55_in_data = data_store_4_54;
		end else begin
			data_in_4_55_in_data = 0;
		end
	end
	// controller for data_in_4_57.data_in_4_57_in_data
	always @(*) begin
		if (eq_221_out) begin 
			data_in_4_57_in_data = data_store_3_46;
		end else if (eq_222_out) begin 
			data_in_4_57_in_data = data_store_4_56;
		end else begin
			data_in_4_57_in_data = 0;
		end
	end
	// controller for data_in_4_59.data_in_4_59_in_data
	always @(*) begin
		if (eq_221_out) begin 
			data_in_4_59_in_data = data_store_3_47;
		end else if (eq_222_out) begin 
			data_in_4_59_in_data = data_store_4_58;
		end else begin
			data_in_4_59_in_data = 0;
		end
	end
	// controller for data_in_5_61.data_in_5_61_in_data
	always @(*) begin
		if (eq_223_out) begin 
			data_in_5_61_in_data = data_store_4_48;
		end else if (eq_224_out) begin 
			data_in_5_61_in_data = data_store_5_60;
		end else begin
			data_in_5_61_in_data = 0;
		end
	end
	// controller for data_in_5_63.data_in_5_63_in_data
	always @(*) begin
		if (eq_223_out) begin 
			data_in_5_63_in_data = data_store_4_50;
		end else if (eq_224_out) begin 
			data_in_5_63_in_data = data_store_5_62;
		end else begin
			data_in_5_63_in_data = 0;
		end
	end
	// controller for data_in_5_65.data_in_5_65_in_data
	always @(*) begin
		if (eq_223_out) begin 
			data_in_5_65_in_data = data_store_4_52;
		end else if (eq_224_out) begin 
			data_in_5_65_in_data = data_store_5_64;
		end else begin
			data_in_5_65_in_data = 0;
		end
	end
	// controller for data_in_5_67.data_in_5_67_in_data
	always @(*) begin
		if (eq_223_out) begin 
			data_in_5_67_in_data = data_store_4_54;
		end else if (eq_224_out) begin 
			data_in_5_67_in_data = data_store_5_66;
		end else begin
			data_in_5_67_in_data = 0;
		end
	end
	// controller for data_in_5_69.data_in_5_69_in_data
	always @(*) begin
		if (eq_223_out) begin 
			data_in_5_69_in_data = data_store_4_56;
		end else if (eq_224_out) begin 
			data_in_5_69_in_data = data_store_5_68;
		end else begin
			data_in_5_69_in_data = 0;
		end
	end
	// controller for data_in_5_71.data_in_5_71_in_data
	always @(*) begin
		if (eq_223_out) begin 
			data_in_5_71_in_data = data_store_4_58;
		end else if (eq_224_out) begin 
			data_in_5_71_in_data = data_store_5_70;
		end else begin
			data_in_5_71_in_data = 0;
		end
	end
	// controller for data_in_6_73.data_in_6_73_in_data
	always @(*) begin
		if (eq_225_out) begin 
			data_in_6_73_in_data = data_store_5_60;
		end else if (eq_226_out) begin 
			data_in_6_73_in_data = data_store_6_72;
		end else begin
			data_in_6_73_in_data = 0;
		end
	end
	// controller for data_in_6_75.data_in_6_75_in_data
	always @(*) begin
		if (eq_225_out) begin 
			data_in_6_75_in_data = data_store_5_62;
		end else if (eq_226_out) begin 
			data_in_6_75_in_data = data_store_6_74;
		end else begin
			data_in_6_75_in_data = 0;
		end
	end
	// controller for data_in_6_77.data_in_6_77_in_data
	always @(*) begin
		if (eq_225_out) begin 
			data_in_6_77_in_data = data_store_5_64;
		end else if (eq_226_out) begin 
			data_in_6_77_in_data = data_store_6_76;
		end else begin
			data_in_6_77_in_data = 0;
		end
	end
	// controller for data_in_6_79.data_in_6_79_in_data
	always @(*) begin
		if (eq_225_out) begin 
			data_in_6_79_in_data = data_store_5_66;
		end else if (eq_226_out) begin 
			data_in_6_79_in_data = data_store_6_78;
		end else begin
			data_in_6_79_in_data = 0;
		end
	end
	// controller for data_in_6_81.data_in_6_81_in_data
	always @(*) begin
		if (eq_225_out) begin 
			data_in_6_81_in_data = data_store_5_68;
		end else if (eq_226_out) begin 
			data_in_6_81_in_data = data_store_6_80;
		end else begin
			data_in_6_81_in_data = 0;
		end
	end
	// controller for data_in_6_82.data_in_6_82_in_data
	always @(*) begin
		if (eq_225_out) begin 
			data_in_6_82_in_data = data_store_5_70;
		end else if (eq_226_out) begin 
			data_in_6_82_in_data = 1'd0;
		end else begin
			data_in_6_82_in_data = 0;
		end
	end
	// controller for eq_122.eq_122_in0
	// controller for eq_122.eq_122_in1
	// Insensitive connections
	assign eq_122_in0 = 32'd0;
	assign eq_122_in1 = state_0_entry_BB_reg;
	// controller for eq_123.eq_123_in0
	// controller for eq_123.eq_123_in1
	// Insensitive connections
	assign eq_123_in0 = 32'd1;
	assign eq_123_in1 = state_0_entry_BB_reg;
	// controller for eq_125.eq_125_in0
	// controller for eq_125.eq_125_in1
	// Insensitive connections
	assign eq_125_in0 = 32'd4;
	assign eq_125_in1 = state_0_entry_BB_reg;
	// controller for eq_127.eq_127_in0
	// controller for eq_127.eq_127_in1
	// Insensitive connections
	assign eq_127_in0 = 32'd4;
	assign eq_127_in1 = state_1_entry_BB_reg;
	// controller for eq_128.eq_128_in0
	// controller for eq_128.eq_128_in1
	// Insensitive connections
	assign eq_128_in0 = 32'd4;
	assign eq_128_in1 = state_2_entry_BB_reg;
	// controller for eq_129.eq_129_in0
	// controller for eq_129.eq_129_in1
	// Insensitive connections
	assign eq_129_in0 = 32'd3;
	assign eq_129_in1 = state_3_entry_BB_reg;
	// controller for eq_130.eq_130_in0
	// controller for eq_130.eq_130_in1
	// Insensitive connections
	assign eq_130_in0 = 32'd3;
	assign eq_130_in1 = state_4_entry_BB_reg;
	// controller for eq_131.eq_131_in0
	// controller for eq_131.eq_131_in1
	// Insensitive connections
	assign eq_131_in0 = 32'd3;
	assign eq_131_in1 = state_5_entry_BB_reg;
	// controller for eq_132.eq_132_in0
	// controller for eq_132.eq_132_in1
	// Insensitive connections
	assign eq_132_in0 = 32'd3;
	assign eq_132_in1 = state_6_entry_BB_reg;
	// controller for eq_133.eq_133_in0
	// controller for eq_133.eq_133_in1
	// Insensitive connections
	assign eq_133_in0 = 32'd2;
	assign eq_133_in1 = state_6_entry_BB_reg;
	// controller for eq_135.eq_135_in0
	// controller for eq_135.eq_135_in1
	// Insensitive connections
	assign eq_135_in0 = 32'd0;
	assign eq_135_in1 = state_0_entry_BB_reg;
	// controller for eq_136.eq_136_in0
	// controller for eq_136.eq_136_in1
	// Insensitive connections
	assign eq_136_in0 = 32'd1;
	assign eq_136_in1 = state_0_entry_BB_reg;
	// controller for eq_139.eq_139_in0
	// controller for eq_139.eq_139_in1
	// Insensitive connections
	assign eq_139_in0 = 32'd4;
	assign eq_139_in1 = state_0_entry_BB_reg;
	// controller for eq_142.eq_142_in0
	// controller for eq_142.eq_142_in1
	// Insensitive connections
	assign eq_142_in0 = 32'd4;
	assign eq_142_in1 = state_1_entry_BB_reg;
	// controller for eq_143.eq_143_in0
	// controller for eq_143.eq_143_in1
	// Insensitive connections
	assign eq_143_in0 = 32'd4;
	assign eq_143_in1 = state_2_entry_BB_reg;
	// controller for eq_144.eq_144_in0
	// controller for eq_144.eq_144_in1
	// Insensitive connections
	assign eq_144_in0 = 32'd3;
	assign eq_144_in1 = state_3_entry_BB_reg;
	// controller for eq_145.eq_145_in0
	// controller for eq_145.eq_145_in1
	// Insensitive connections
	assign eq_145_in0 = 32'd3;
	assign eq_145_in1 = state_4_entry_BB_reg;
	// controller for eq_146.eq_146_in0
	// controller for eq_146.eq_146_in1
	// Insensitive connections
	assign eq_146_in0 = 32'd3;
	assign eq_146_in1 = state_5_entry_BB_reg;
	// controller for eq_147.eq_147_in0
	// controller for eq_147.eq_147_in1
	// Insensitive connections
	assign eq_147_in0 = 32'd3;
	assign eq_147_in1 = state_6_entry_BB_reg;
	// controller for eq_148.eq_148_in0
	// controller for eq_148.eq_148_in1
	// Insensitive connections
	assign eq_148_in0 = 32'd2;
	assign eq_148_in1 = state_6_entry_BB_reg;
	// controller for eq_202.eq_202_in0
	// controller for eq_202.eq_202_in1
	// Insensitive connections
	assign eq_202_in0 = 32'd0;
	assign eq_202_in1 = state_0_last_state;
	// controller for eq_203.eq_203_in0
	// controller for eq_203.eq_203_in1
	// Insensitive connections
	assign eq_203_in0 = 32'd2;
	assign eq_203_in1 = state_0_last_state;
	// controller for eq_204.eq_204_in0
	// controller for eq_204.eq_204_in1
	// Insensitive connections
	assign eq_204_in0 = 32'd6;
	assign eq_204_in1 = state_0_last_state;
	// controller for eq_211.eq_211_in0
	// controller for eq_211.eq_211_in1
	// Insensitive connections
	assign eq_211_in0 = 32'd0;
	assign eq_211_in1 = state_1_last_state;
	// controller for eq_212.eq_212_in0
	// controller for eq_212.eq_212_in1
	// Insensitive connections
	assign eq_212_in0 = 32'd1;
	assign eq_212_in1 = state_1_last_state;
	// controller for eq_214.eq_214_in0
	// controller for eq_214.eq_214_in1
	// Insensitive connections
	assign eq_214_in0 = 32'd1;
	assign eq_214_in1 = state_2_last_state;
	// controller for eq_215.eq_215_in0
	// controller for eq_215.eq_215_in1
	// Insensitive connections
	assign eq_215_in0 = 32'd2;
	assign eq_215_in1 = state_2_last_state;
	// controller for eq_217.eq_217_in0
	// controller for eq_217.eq_217_in1
	// Insensitive connections
	assign eq_217_in0 = 32'd2;
	assign eq_217_in1 = state_3_last_state;
	// controller for eq_218.eq_218_in0
	// controller for eq_218.eq_218_in1
	// Insensitive connections
	assign eq_218_in0 = 32'd3;
	assign eq_218_in1 = state_3_last_state;
	// controller for eq_221.eq_221_in0
	// controller for eq_221.eq_221_in1
	// Insensitive connections
	assign eq_221_in0 = 32'd3;
	assign eq_221_in1 = state_4_last_state;
	// controller for eq_222.eq_222_in0
	// controller for eq_222.eq_222_in1
	// Insensitive connections
	assign eq_222_in0 = 32'd4;
	assign eq_222_in1 = state_4_last_state;
	// controller for eq_223.eq_223_in0
	// controller for eq_223.eq_223_in1
	// Insensitive connections
	assign eq_223_in0 = 32'd4;
	assign eq_223_in1 = state_5_last_state;
	// controller for eq_224.eq_224_in0
	// controller for eq_224.eq_224_in1
	// Insensitive connections
	assign eq_224_in0 = 32'd5;
	assign eq_224_in1 = state_5_last_state;
	// controller for eq_225.eq_225_in0
	// controller for eq_225.eq_225_in1
	// Insensitive connections
	assign eq_225_in0 = 32'd5;
	assign eq_225_in1 = state_6_last_state;
	// controller for eq_226.eq_226_in0
	// controller for eq_226.eq_226_in1
	// Insensitive connections
	assign eq_226_in0 = 32'd6;
	assign eq_226_in1 = state_6_last_state;
	// controller for icmp_icmp22.icmp_icmp22_in0
	// controller for icmp_icmp22.icmp_icmp22_in1
	// Insensitive connections
	assign icmp_icmp22_in0 = add_add21_out;
	assign icmp_icmp22_in1 = 32'd3;
	// controller for icmp_icmp4.icmp_icmp4_in0
	// controller for icmp_icmp4.icmp_icmp4_in1
	// Insensitive connections
	assign icmp_icmp4_in0 = add_add3_out;
	assign icmp_icmp4_in1 = 32'd3;
	// controller for mul_mul16.mul_mul16_in0
	// controller for mul_mul16.mul_mul16_in1
	// Insensitive connections
	assign mul_mul16_in0 = data_in_2_26_out_data;
	assign mul_mul16_in1 = ram_rdata_1;
	// controller for mul_mul5.mul_mul5_in0
	// controller for mul_mul5.mul_mul5_in1
	// Insensitive connections
	assign mul_mul5_in0 = phi_phi1_out;
	assign mul_mul5_in1 = 32'd3;
	// controller for notOp_100.notOp_100_in0
	// Insensitive connections
	assign notOp_100_in0 = data_in_2_32_out_data;
	// controller for notOp_103.notOp_103_in0
	// Insensitive connections
	assign notOp_103_in0 = andOp_102_out;
	// controller for notOp_105.notOp_105_in0
	// Insensitive connections
	assign notOp_105_in0 = data_in_6_82_out_data;
	// controller for notOp_108.notOp_108_in0
	// Insensitive connections
	assign notOp_108_in0 = andOp_107_out;
	// controller for notOp_110.notOp_110_in0
	// Insensitive connections
	assign notOp_110_in0 = data_in_6_82_out_data;
	// controller for notOp_113.notOp_113_in0
	// Insensitive connections
	assign notOp_113_in0 = andOp_112_out;
	// controller for notOp_115.notOp_115_in0
	// Insensitive connections
	assign notOp_115_in0 = data_in_6_82_out_data;
	// controller for notOp_118.notOp_118_in0
	// Insensitive connections
	assign notOp_118_in0 = andOp_117_out;
	// controller for notOp_120.notOp_120_in0
	// Insensitive connections
	assign notOp_120_in0 = data_in_6_82_out_data;
	// controller for notOp_137.notOp_137_in0
	// Insensitive connections
	assign notOp_137_in0 = eq_136_out;
	// controller for notOp_140.notOp_140_in0
	// Insensitive connections
	assign notOp_140_in0 = eq_139_out;
	// controller for notOp_149.notOp_149_in0
	// Insensitive connections
	assign notOp_149_in0 = eq_148_out;
	// controller for notOp_184.notOp_184_in0
	// Insensitive connections
	assign notOp_184_in0 = andOp_106_out;
	// controller for notOp_186.notOp_186_in0
	// Insensitive connections
	assign notOp_186_in0 = andOp_91_out;
	// controller for notOp_188.notOp_188_in0
	// Insensitive connections
	assign notOp_188_in0 = andOp_178_out;
	// controller for notOp_190.notOp_190_in0
	// Insensitive connections
	assign notOp_190_in0 = andOp_179_out;
	// controller for notOp_192.notOp_192_in0
	// Insensitive connections
	assign notOp_192_in0 = andOp_89_out;
	// controller for notOp_194.notOp_194_in0
	// Insensitive connections
	assign notOp_194_in0 = andOp_180_out;
	// controller for notOp_196.notOp_196_in0
	// Insensitive connections
	assign notOp_196_in0 = andOp_181_out;
	// controller for notOp_198.notOp_198_in0
	// Insensitive connections
	assign notOp_198_in0 = andOp_182_out;
	// controller for notOp_200.notOp_200_in0
	// Insensitive connections
	assign notOp_200_in0 = andOp_183_out;
	// controller for notOp_84.notOp_84_in0
	// Insensitive connections
	assign notOp_84_in0 = andOp_83_out;
	// controller for notOp_86.notOp_86_in0
	// Insensitive connections
	assign notOp_86_in0 = andOp_85_out;
	// controller for notOp_88.notOp_88_in0
	// Insensitive connections
	assign notOp_88_in0 = andOp_87_out;
	// controller for notOp_90.notOp_90_in0
	// Insensitive connections
	assign notOp_90_in0 = data_in_2_32_out_data;
	// controller for notOp_93.notOp_93_in0
	// Insensitive connections
	assign notOp_93_in0 = andOp_92_out;
	// controller for notOp_95.notOp_95_in0
	// Insensitive connections
	assign notOp_95_in0 = data_in_2_32_out_data;
	// controller for notOp_98.notOp_98_in0
	// Insensitive connections
	assign notOp_98_in0 = andOp_97_out;
	// controller for orOp_124.orOp_124_in0
	// controller for orOp_124.orOp_124_in1
	// Insensitive connections
	assign orOp_124_in0 = eq_123_out;
	assign orOp_124_in1 = andOp_83_out;
	// controller for orOp_126.orOp_126_in0
	// controller for orOp_126.orOp_126_in1
	// Insensitive connections
	assign orOp_126_in0 = eq_125_out;
	assign orOp_126_in1 = andOp_85_out;
	// controller for orOp_134.orOp_134_in0
	// controller for orOp_134.orOp_134_in1
	// Insensitive connections
	assign orOp_134_in0 = eq_133_out;
	assign orOp_134_in1 = andOp_104_out;
	// controller for phi_phi1.phi_phi1_in
	// controller for phi_phi1.phi_phi1_last_block
	// controller for phi_phi1.phi_phi1_s
	// Insensitive connections
	assign phi_phi1_in = concat_159_out;
	assign phi_phi1_last_block = bb_1_predecessor_in_state_0_out_data;
	assign phi_phi1_s = concat_160_out;
	// controller for phi_phi6.phi_phi6_in
	// controller for phi_phi6.phi_phi6_last_block
	// controller for phi_phi6.phi_phi6_s
	// Insensitive connections
	assign phi_phi6_in = concat_165_out;
	assign phi_phi6_last_block = bb_4_predecessor_in_state_0_out_data;
	assign phi_phi6_s = concat_166_out;
	// controller for phi_phi9.phi_phi9_in
	// controller for phi_phi9.phi_phi9_last_block
	// controller for phi_phi9.phi_phi9_s
	// Insensitive connections
	assign phi_phi9_in = concat_169_out;
	assign phi_phi9_last_block = bb_4_predecessor_in_state_0_out_data;
	assign phi_phi9_s = concat_170_out;
	// controller for ram.ram_raddr_1_reg
	always @(*) begin
		if (andOp_153_out) begin 
			ram_raddr_1_reg = add_add12_out;
		end else begin
			ram_raddr_1_reg = 0;
		end
	end
	// controller for ram.ram_raddr_2_reg
	always @(*) begin
		if (andOp_151_out) begin 
			ram_raddr_2_reg = add_add7_out;
		end else begin
			ram_raddr_2_reg = 0;
		end
	end
	// controller for ram.ram_waddr_0_reg
	always @(*) begin
		if (andOp_156_out) begin 
			ram_waddr_0_reg = add_add20_out;
		end else begin
			ram_waddr_0_reg = 0;
		end
	end
	// controller for ram.ram_wdata_0_reg
	always @(*) begin
		if (andOp_157_out) begin 
			ram_wdata_0_reg = data_in_3_41_out_data;
		end else begin
			ram_wdata_0_reg = 0;
		end
	end
	// controller for ram.ram_wen_0_reg
	always @(*) begin
		if (andOp_155_out) begin 
			ram_wen_0_reg = -(1'd1);
		end else begin
			ram_wen_0_reg = 0;
		end
	end
	// controller for ret24.valid_reg
	always @(*) begin
		if (andOp_177_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			data_store_0_0 <= 0;
		end else begin
			if (andOp_205_out) begin
				data_store_0_0 <= phi_phi1_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_10 <= 0;
		end else begin
			if (andOp_209_out) begin
				data_store_0_10 <= phi_phi6_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_11 <= 0;
		end else begin
			if (andOp_210_out) begin
				data_store_0_11 <= phi_phi9_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_3 <= 0;
		end else begin
			if (andOp_206_out) begin
				data_store_0_3 <= add_add3_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_5 <= 0;
		end else begin
			if (andOp_207_out) begin
				data_store_0_5 <= icmp_icmp4_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_6 <= 0;
		end else begin
			if (andOp_208_out) begin
				data_store_0_6 <= mul_mul5_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_8 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_8 <= data_in_0_9_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_12 <= 0;
		end else begin
			if (andOp_213_out) begin
				data_store_1_12 <= ram_rdata_2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_13 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_13 <= data_in_1_14_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_15 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_15 <= data_in_1_16_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_17 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_17 <= data_in_1_18_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_19 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_19 <= data_in_1_20_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_21 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_21 <= data_in_1_22_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_24 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_24 <= data_in_1_25_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_27 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_27 <= data_in_2_28_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_29 <= 0;
		end else begin
			if (andOp_216_out) begin
				data_store_2_29 <= add_add13_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_30 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_30 <= data_in_2_31_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_33 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_33 <= data_in_2_34_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_35 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_35 <= data_in_2_36_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_38 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_38 <= data_in_3_39_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_40 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_40 <= data_in_3_41_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_42 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_42 <= data_in_3_43_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_44 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_44 <= data_in_3_45_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_46 <= 0;
		end else begin
			if (andOp_219_out) begin
				data_store_3_46 <= add_add21_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_47 <= 0;
		end else begin
			if (andOp_220_out) begin
				data_store_3_47 <= icmp_icmp22_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_48 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_48 <= data_in_4_49_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_50 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_50 <= data_in_4_51_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_52 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_52 <= data_in_4_53_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_54 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_54 <= data_in_4_55_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_56 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_56 <= data_in_4_57_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_58 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_58 <= data_in_4_59_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_60 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_60 <= data_in_5_61_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_62 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_62 <= data_in_5_63_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_64 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_64 <= data_in_5_65_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_66 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_66 <= data_in_5_67_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_68 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_68 <= data_in_5_69_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_70 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_70 <= data_in_5_71_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_72 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_72 <= data_in_6_73_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_74 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_74 <= data_in_6_75_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_76 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_76 <= data_in_6_77_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_78 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_78 <= data_in_6_79_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_80 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_80 <= data_in_6_81_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_106_out) begin
				global_state <= 32'd0;
			end
			if (andOp_178_out) begin
				global_state <= 32'd1;
			end
			if (andOp_179_out) begin
				global_state <= 32'd2;
			end
			if (andOp_180_out) begin
				global_state <= 32'd4;
			end
			if (andOp_181_out) begin
				global_state <= 32'd5;
			end
			if (andOp_182_out) begin
				global_state <= 32'd6;
			end
			if (andOp_183_out) begin
				global_state <= 32'd6;
			end
			if (andOp_89_out) begin
				global_state <= 32'd3;
			end
			if (andOp_91_out) begin
				global_state <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
			if (andOp_106_out) begin
				state_0_entry_BB_reg <= 32'd1;
			end
			if (andOp_91_out) begin
				state_0_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (andOp_106_out) begin
				state_0_is_active <= 1'd1;
			end
			if (andOp_187_out) begin
				state_0_is_active <= 1'd0;
			end
			if (andOp_91_out) begin
				state_0_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
			if (andOp_106_out) begin
				state_0_last_BB_reg <= 32'd3;
			end
			if (andOp_91_out) begin
				state_0_last_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
			if (andOp_106_out) begin
				state_0_last_state <= 32'd6;
			end
			if (andOp_91_out) begin
				state_0_last_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_178_out) begin
				state_1_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_178_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_189_out) begin
				state_1_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_178_out) begin
				state_1_last_BB_reg <= bb_4_predecessor_in_state_0_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_178_out) begin
				state_1_last_state <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_179_out) begin
				state_2_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_179_out) begin
				state_2_is_active <= 1'd1;
			end
			if (andOp_191_out) begin
				state_2_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_179_out) begin
				state_2_last_BB_reg <= bb_4_predecessor_in_state_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_179_out) begin
				state_2_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_89_out) begin
				state_3_entry_BB_reg <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_193_out) begin
				state_3_is_active <= 1'd0;
			end
			if (andOp_89_out) begin
				state_3_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_89_out) begin
				state_3_last_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_state <= 0;
		end else begin
			if (andOp_89_out) begin
				state_3_last_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_180_out) begin
				state_4_entry_BB_reg <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_180_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_195_out) begin
				state_4_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_180_out) begin
				state_4_last_BB_reg <= bb_3_predecessor_in_state_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_state <= 0;
		end else begin
			if (andOp_180_out) begin
				state_4_last_state <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_entry_BB_reg <= 0;
		end else begin
			if (andOp_181_out) begin
				state_5_entry_BB_reg <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_is_active <= 0;
		end else begin
			if (andOp_181_out) begin
				state_5_is_active <= 1'd1;
			end
			if (andOp_197_out) begin
				state_5_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_last_BB_reg <= 0;
		end else begin
			if (andOp_181_out) begin
				state_5_last_BB_reg <= bb_3_predecessor_in_state_4_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_last_state <= 0;
		end else begin
			if (andOp_181_out) begin
				state_5_last_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_entry_BB_reg <= 0;
		end else begin
			if (andOp_182_out) begin
				state_6_entry_BB_reg <= 32'd3;
			end
			if (andOp_183_out) begin
				state_6_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_is_active <= 0;
		end else begin
			if (andOp_182_out) begin
				state_6_is_active <= 1'd1;
			end
			if (andOp_183_out) begin
				state_6_is_active <= 1'd1;
			end
			if (andOp_201_out) begin
				state_6_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_last_BB_reg <= 0;
		end else begin
			if (andOp_182_out) begin
				state_6_last_BB_reg <= bb_3_predecessor_in_state_5_out_data;
			end
			if (andOp_183_out) begin
				state_6_last_BB_reg <= bb_2_predecessor_in_state_6_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_last_state <= 0;
		end else begin
			if (andOp_182_out) begin
				state_6_last_state <= 32'd5;
			end
			if (andOp_183_out) begin
				state_6_last_state <= 32'd6;
			end
		end
	end

endmodule

