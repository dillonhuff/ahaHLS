module temp_storage_pipe(input [0:0] clk, input [0:0] rst, output [0:0] valid, output [3:0] arg_0_debug_addr, input [31:0] arg_0_debug_data, output [3:0] arg_0_debug_write_addr, output [31:0] arg_0_debug_write_data, output [0:0] arg_0_debug_write_en, output [3:0] arg_0_raddr_0, input [31:0] arg_0_rdata_0, output [0:0] arg_0_rst, output [3:0] arg_0_waddr_0, output [31:0] arg_0_wdata_0, output [0:0] arg_0_wen_0, output [3:0] arg_1_debug_addr, input [31:0] arg_1_debug_data, output [3:0] arg_1_debug_write_addr, output [31:0] arg_1_debug_write_data, output [0:0] arg_1_debug_write_en, output [3:0] arg_1_raddr_0, input [31:0] arg_1_rdata_0, output [0:0] arg_1_rst, output [3:0] arg_1_waddr_0, output [31:0] arg_1_wdata_0, output [0:0] arg_1_wen_0);

	reg [0:0] valid_reg;
	reg [3:0] arg_0_debug_addr_reg;
	reg [3:0] arg_0_debug_write_addr_reg;
	reg [31:0] arg_0_debug_write_data_reg;
	reg [0:0] arg_0_debug_write_en_reg;
	reg [3:0] arg_0_raddr_0_reg;
	reg [0:0] arg_0_rst_reg;
	reg [3:0] arg_0_waddr_0_reg;
	reg [31:0] arg_0_wdata_0_reg;
	reg [0:0] arg_0_wen_0_reg;
	reg [3:0] arg_1_debug_addr_reg;
	reg [3:0] arg_1_debug_write_addr_reg;
	reg [31:0] arg_1_debug_write_data_reg;
	reg [0:0] arg_1_debug_write_en_reg;
	reg [3:0] arg_1_raddr_0_reg;
	reg [0:0] arg_1_rst_reg;
	reg [3:0] arg_1_waddr_0_reg;
	reg [31:0] arg_1_wdata_0_reg;
	reg [0:0] arg_1_wen_0_reg;

	assign valid = valid_reg;
	assign arg_0_debug_addr = arg_0_debug_addr_reg;
	assign arg_0_debug_write_addr = arg_0_debug_write_addr_reg;
	assign arg_0_debug_write_data = arg_0_debug_write_data_reg;
	assign arg_0_debug_write_en = arg_0_debug_write_en_reg;
	assign arg_0_raddr_0 = arg_0_raddr_0_reg;
	assign arg_0_rst = arg_0_rst_reg;
	assign arg_0_waddr_0 = arg_0_waddr_0_reg;
	assign arg_0_wdata_0 = arg_0_wdata_0_reg;
	assign arg_0_wen_0 = arg_0_wen_0_reg;
	assign arg_1_debug_addr = arg_1_debug_addr_reg;
	assign arg_1_debug_write_addr = arg_1_debug_write_addr_reg;
	assign arg_1_debug_write_data = arg_1_debug_write_data_reg;
	assign arg_1_debug_write_en = arg_1_debug_write_en_reg;
	assign arg_1_raddr_0 = arg_1_raddr_0_reg;
	assign arg_1_rst = arg_1_rst_reg;
	assign arg_1_waddr_0 = arg_1_waddr_0_reg;
	assign arg_1_wdata_0 = arg_1_wdata_0_reg;
	assign arg_1_wen_0 = arg_1_wen_0_reg;

	// Start debug wires and ports

	initial begin
	end



	always @(posedge clk) begin
		if (!((!(andOp_12_out === 1) || andOp_16_out !== 1))) begin $display("assertion((!(andOp_12_out === 1) || andOp_16_out !== 1))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_16_out === 1) || andOp_12_out !== 1))) begin $display("assertion((!(andOp_16_out === 1) || andOp_12_out !== 1))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_111_out === 1) || andOp_18_out !== 1))) begin $display("assertion((!(andOp_111_out === 1) || andOp_18_out !== 1))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_18_out === 1) || andOp_111_out !== 1))) begin $display("assertion((!(andOp_18_out === 1) || andOp_111_out !== 1))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_12_out === 1) || andOp_16_out !== 1))) begin $display("assertion((!(andOp_12_out === 1) || andOp_16_out !== 1))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_16_out === 1) || andOp_12_out !== 1))) begin $display("assertion((!(andOp_16_out === 1) || andOp_12_out !== 1))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_111_out === 1) || andOp_98_out !== 1))) begin $display("assertion((!(andOp_111_out === 1) || andOp_98_out !== 1))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_98_out === 1) || andOp_111_out !== 1))) begin $display("assertion((!(andOp_98_out === 1) || andOp_111_out !== 1))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_105_out === 1) || andOp_115_out !== 1))) begin $display("assertion((!(andOp_105_out === 1) || andOp_115_out !== 1)) failed: Overlapping state active transition for state 1"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_105_out === 1) || andOp_12_out !== 1))) begin $display("assertion((!(andOp_105_out === 1) || andOp_12_out !== 1)) failed: Overlapping state active transition for state 1"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_115_out === 1) || andOp_105_out !== 1))) begin $display("assertion((!(andOp_115_out === 1) || andOp_105_out !== 1)) failed: Overlapping state active transition for state 1"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_115_out === 1) || andOp_12_out !== 1))) begin $display("assertion((!(andOp_115_out === 1) || andOp_12_out !== 1)) failed: Overlapping state active transition for state 1"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_12_out === 1) || andOp_105_out !== 1))) begin $display("assertion((!(andOp_12_out === 1) || andOp_105_out !== 1)) failed: Overlapping state active transition for state 1"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_12_out === 1) || andOp_115_out !== 1))) begin $display("assertion((!(andOp_12_out === 1) || andOp_115_out !== 1)) failed: Overlapping state active transition for state 1"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_106_out === 1) || andOp_117_out !== 1))) begin $display("assertion((!(andOp_106_out === 1) || andOp_117_out !== 1)) failed: Overlapping state active transition for state 2"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_117_out === 1) || andOp_106_out !== 1))) begin $display("assertion((!(andOp_117_out === 1) || andOp_106_out !== 1)) failed: Overlapping state active transition for state 2"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_107_out === 1) || andOp_119_out !== 1))) begin $display("assertion((!(andOp_107_out === 1) || andOp_119_out !== 1)) failed: Overlapping state active transition for state 3"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_119_out === 1) || andOp_107_out !== 1))) begin $display("assertion((!(andOp_119_out === 1) || andOp_107_out !== 1)) failed: Overlapping state active transition for state 3"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_108_out === 1) || andOp_121_out !== 1))) begin $display("assertion((!(andOp_108_out === 1) || andOp_121_out !== 1)) failed: Overlapping state active transition for state 4"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_121_out === 1) || andOp_108_out !== 1))) begin $display("assertion((!(andOp_121_out === 1) || andOp_108_out !== 1)) failed: Overlapping state active transition for state 4"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_109_out === 1) || andOp_123_out !== 1))) begin $display("assertion((!(andOp_109_out === 1) || andOp_123_out !== 1)) failed: Overlapping state active transition for state 5"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_123_out === 1) || andOp_109_out !== 1))) begin $display("assertion((!(andOp_123_out === 1) || andOp_109_out !== 1)) failed: Overlapping state active transition for state 5"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_110_out === 1) || andOp_125_out !== 1))) begin $display("assertion((!(andOp_110_out === 1) || andOp_125_out !== 1)) failed: Overlapping state active transition for state 6"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_125_out === 1) || andOp_110_out !== 1))) begin $display("assertion((!(andOp_125_out === 1) || andOp_110_out !== 1)) failed: Overlapping state active transition for state 6"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_111_out === 1) || andOp_129_out !== 1))) begin $display("assertion((!(andOp_111_out === 1) || andOp_129_out !== 1)) failed: Overlapping state active transition for state 7"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_111_out === 1) || andOp_86_out !== 1))) begin $display("assertion((!(andOp_111_out === 1) || andOp_86_out !== 1)) failed: Overlapping state active transition for state 7"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_129_out === 1) || andOp_111_out !== 1))) begin $display("assertion((!(andOp_129_out === 1) || andOp_111_out !== 1)) failed: Overlapping state active transition for state 7"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_129_out === 1) || andOp_86_out !== 1))) begin $display("assertion((!(andOp_129_out === 1) || andOp_86_out !== 1)) failed: Overlapping state active transition for state 7"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_86_out === 1) || andOp_111_out !== 1))) begin $display("assertion((!(andOp_86_out === 1) || andOp_111_out !== 1)) failed: Overlapping state active transition for state 7"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_86_out === 1) || andOp_129_out !== 1))) begin $display("assertion((!(andOp_86_out === 1) || andOp_129_out !== 1)) failed: Overlapping state active transition for state 7"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_1_is_active) || !(1'd0)))) begin $display("assertion((!(state_1_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_2_is_active) || !(1'd0)))) begin $display("assertion((!(state_2_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_3_is_active) || !(1'd0)))) begin $display("assertion((!(state_3_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_4_is_active) || !(1'd0)))) begin $display("assertion((!(state_4_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_5_is_active) || !(1'd0)))) begin $display("assertion((!(state_5_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_6_is_active) || !(1'd0)))) begin $display("assertion((!(state_6_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_7_is_active) || !(1'd0)))) begin $display("assertion((!(state_7_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_0_is_active) || !(1'd0)))) begin $display("assertion((!(state_0_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_1_is_active) || !(1'd0)))) begin $display("assertion((!(state_1_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_2_is_active) || !(1'd0)))) begin $display("assertion((!(state_2_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_3_is_active) || !(1'd0)))) begin $display("assertion((!(state_3_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_4_is_active) || !(1'd0)))) begin $display("assertion((!(state_4_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_5_is_active) || !(1'd0)))) begin $display("assertion((!(state_5_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_6_is_active) || !(1'd0)))) begin $display("assertion((!(state_6_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_0_is_active) || !(1'd0)))) begin $display("assertion((!(state_0_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_7_is_active) || !(1'd0)))) begin $display("assertion((!(state_7_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(notOp_156_out || icmp_icmp3_in0 !== 32'dx)) begin $display("assertion(notOp_156_out || icmp_icmp3_in0 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(notOp_157_out || icmp_icmp3_in1 !== 32'dx)) begin $display("assertion(notOp_157_out || icmp_icmp3_in1 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_158_out) || add_add2_in0 !== 32'dx)) begin $display("assertion(!(andOp_158_out) || add_add2_in0 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_158_out) || add_add2_in1 !== 32'dx)) begin $display("assertion(!(andOp_158_out) || add_add2_in1 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_159_out) || add_add10_in0 !== 32'dx)) begin $display("assertion(!(andOp_159_out) || add_add10_in0 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_159_out) || add_add10_in1 !== 32'dx)) begin $display("assertion(!(andOp_159_out) || add_add10_in1 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_160_out) || mul_mul6_in0 !== 32'dx)) begin $display("assertion(!(andOp_160_out) || mul_mul6_in0 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_160_out) || mul_mul6_in1 !== 32'dx)) begin $display("assertion(!(andOp_160_out) || mul_mul6_in1 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_161_out) || mul_mul9_in0 !== 32'dx)) begin $display("assertion(!(andOp_161_out) || mul_mul9_in0 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_161_out) || mul_mul9_in1 !== 32'dx)) begin $display("assertion(!(andOp_161_out) || mul_mul9_in1 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_162_out) || phi_phi1_out !== 'dx))) begin $display("assertion((!(andOp_162_out) || phi_phi1_out !== 'dx))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_163_out) || data_in_3_9_out_data !== 32'dx))) begin $display("assertion((!(andOp_163_out) || data_in_3_9_out_data !== 32'dx))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_164_out) || add_add10_out !== 32'dx))) begin $display("assertion((!(andOp_164_out) || add_add10_out !== 32'dx))"); $finish(); end
	end




	// End debug wires and ports

	// Start Functional Units
	wire [63:0] phi_phi1_in;
	wire [31:0] phi_phi1_last_block;
	wire [63:0] phi_phi1_s;
	wire [31:0] phi_phi1_out;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_phi1(.in(phi_phi1_in), .last_block(phi_phi1_last_block), .out(phi_phi1_out), .s(phi_phi1_s));

	wire [31:0] add_add2_in0;
	wire [31:0] add_add2_in1;
	wire [31:0] add_add2_out;
	add #(.WIDTH(32)) add_add2(.in0(add_add2_in0), .in1(add_add2_in1), .out(add_add2_out));

	wire [31:0] mul_mul6_in0;
	wire [31:0] mul_mul6_in1;
	wire [31:0] mul_mul6_out;
	mul #(.WIDTH(32)) mul_mul6(.in0(mul_mul6_in0), .in1(mul_mul6_in1), .out(mul_mul6_out));

	wire [31:0] mul_mul9_in0;
	wire [31:0] mul_mul9_in1;
	wire [31:0] mul_mul9_out;
	mul #(.WIDTH(32)) mul_mul9(.in0(mul_mul9_in0), .in1(mul_mul9_in1), .out(mul_mul9_out));

	wire [31:0] add_add10_in0;
	wire [31:0] add_add10_in1;
	wire [31:0] add_add10_out;
	add #(.WIDTH(32)) add_add10(.in0(add_add10_in0), .in1(add_add10_in1), .out(add_add10_out));

	wire [31:0] icmp_icmp3_in0;
	wire [31:0] icmp_icmp3_in1;
	wire [0:0] icmp_icmp3_out;
	ne #(.WIDTH(32)) icmp_icmp3(.in0(icmp_icmp3_in0), .in1(icmp_icmp3_in1), .out(icmp_icmp3_out));

	br_dummy br_unit();

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] bb_2_active_in_state_1_in_data;
	wire [0:0] bb_2_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_1(.in_data(bb_2_active_in_state_1_in_data), .out_data(bb_2_active_in_state_1_out_data));

	reg [31:0] bb_2_predecessor_in_state_1_in_data;
	wire [31:0] bb_2_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_1(.in_data(bb_2_predecessor_in_state_1_in_data), .out_data(bb_2_predecessor_in_state_1_out_data));

	reg [0:0] br_2_happened_in_state_1_in_data;
	wire [0:0] br_2_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_2_happened_in_state_1(.in_data(br_2_happened_in_state_1_in_data), .out_data(br_2_happened_in_state_1_out_data));

	reg [0:0] bb_2_active_in_state_2_in_data;
	wire [0:0] bb_2_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_2(.in_data(bb_2_active_in_state_2_in_data), .out_data(bb_2_active_in_state_2_out_data));

	reg [31:0] bb_2_predecessor_in_state_2_in_data;
	wire [31:0] bb_2_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_2(.in_data(bb_2_predecessor_in_state_2_in_data), .out_data(bb_2_predecessor_in_state_2_out_data));

	reg [0:0] br_2_happened_in_state_2_in_data;
	wire [0:0] br_2_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_2_happened_in_state_2(.in_data(br_2_happened_in_state_2_in_data), .out_data(br_2_happened_in_state_2_out_data));

	reg [0:0] bb_2_active_in_state_3_in_data;
	wire [0:0] bb_2_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_3(.in_data(bb_2_active_in_state_3_in_data), .out_data(bb_2_active_in_state_3_out_data));

	reg [31:0] bb_2_predecessor_in_state_3_in_data;
	wire [31:0] bb_2_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_3(.in_data(bb_2_predecessor_in_state_3_in_data), .out_data(bb_2_predecessor_in_state_3_out_data));

	reg [0:0] br_2_happened_in_state_3_in_data;
	wire [0:0] br_2_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_2_happened_in_state_3(.in_data(br_2_happened_in_state_3_in_data), .out_data(br_2_happened_in_state_3_out_data));

	reg [0:0] bb_2_active_in_state_4_in_data;
	wire [0:0] bb_2_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_4(.in_data(bb_2_active_in_state_4_in_data), .out_data(bb_2_active_in_state_4_out_data));

	reg [31:0] bb_2_predecessor_in_state_4_in_data;
	wire [31:0] bb_2_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_4(.in_data(bb_2_predecessor_in_state_4_in_data), .out_data(bb_2_predecessor_in_state_4_out_data));

	reg [0:0] br_2_happened_in_state_4_in_data;
	wire [0:0] br_2_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_2_happened_in_state_4(.in_data(br_2_happened_in_state_4_in_data), .out_data(br_2_happened_in_state_4_out_data));

	reg [0:0] bb_2_active_in_state_5_in_data;
	wire [0:0] bb_2_active_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_5(.in_data(bb_2_active_in_state_5_in_data), .out_data(bb_2_active_in_state_5_out_data));

	reg [31:0] bb_2_predecessor_in_state_5_in_data;
	wire [31:0] bb_2_predecessor_in_state_5_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_5(.in_data(bb_2_predecessor_in_state_5_in_data), .out_data(bb_2_predecessor_in_state_5_out_data));

	reg [0:0] br_2_happened_in_state_5_in_data;
	wire [0:0] br_2_happened_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) br_2_happened_in_state_5(.in_data(br_2_happened_in_state_5_in_data), .out_data(br_2_happened_in_state_5_out_data));

	reg [0:0] bb_2_active_in_state_6_in_data;
	wire [0:0] bb_2_active_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_6(.in_data(bb_2_active_in_state_6_in_data), .out_data(bb_2_active_in_state_6_out_data));

	reg [31:0] bb_2_predecessor_in_state_6_in_data;
	wire [31:0] bb_2_predecessor_in_state_6_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_6(.in_data(bb_2_predecessor_in_state_6_in_data), .out_data(bb_2_predecessor_in_state_6_out_data));

	reg [0:0] br_2_happened_in_state_6_in_data;
	wire [0:0] br_2_happened_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) br_2_happened_in_state_6(.in_data(br_2_happened_in_state_6_in_data), .out_data(br_2_happened_in_state_6_out_data));

	reg [0:0] bb_1_active_in_state_7_in_data;
	wire [0:0] bb_1_active_in_state_7_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_7(.in_data(bb_1_active_in_state_7_in_data), .out_data(bb_1_active_in_state_7_out_data));

	reg [31:0] bb_1_predecessor_in_state_7_in_data;
	wire [31:0] bb_1_predecessor_in_state_7_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_7(.in_data(bb_1_predecessor_in_state_7_in_data), .out_data(bb_1_predecessor_in_state_7_out_data));

	reg [31:0] data_in_0_1_in_data;
	wire [31:0] data_in_0_1_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_1(.in_data(data_in_0_1_in_data), .out_data(data_in_0_1_out_data));

	reg [31:0] data_in_1_4_in_data;
	wire [31:0] data_in_1_4_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_4(.in_data(data_in_1_4_in_data), .out_data(data_in_1_4_out_data));

	reg [31:0] data_in_2_6_in_data;
	wire [31:0] data_in_2_6_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_6(.in_data(data_in_2_6_in_data), .out_data(data_in_2_6_out_data));

	reg [31:0] data_in_3_9_in_data;
	wire [31:0] data_in_3_9_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_9(.in_data(data_in_3_9_in_data), .out_data(data_in_3_9_out_data));

	reg [31:0] data_in_3_10_in_data;
	wire [31:0] data_in_3_10_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_10(.in_data(data_in_3_10_in_data), .out_data(data_in_3_10_out_data));

	reg [31:0] data_in_3_11_in_data;
	wire [31:0] data_in_3_11_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_11(.in_data(data_in_3_11_in_data), .out_data(data_in_3_11_out_data));

	wire [0:0] andOp_12_in0;
	wire [0:0] andOp_12_in1;
	wire [0:0] andOp_12_out;
	andOp #(.WIDTH(1)) andOp_12(.in0(andOp_12_in0), .in1(andOp_12_in1), .out(andOp_12_out));

	wire [0:0] notOp_13_in0;
	wire [0:0] notOp_13_out;
	notOp #(.WIDTH(1)) notOp_13(.in(notOp_13_in0), .out(notOp_13_out));

	wire [0:0] andOp_14_in0;
	wire [0:0] andOp_14_in1;
	wire [0:0] andOp_14_out;
	andOp #(.WIDTH(1)) andOp_14(.in0(andOp_14_in0), .in1(andOp_14_in1), .out(andOp_14_out));

	wire [0:0] notOp_15_in0;
	wire [0:0] notOp_15_out;
	notOp #(.WIDTH(1)) notOp_15(.in(notOp_15_in0), .out(notOp_15_out));

	wire [0:0] andOp_16_in0;
	wire [0:0] andOp_16_in1;
	wire [0:0] andOp_16_out;
	andOp #(.WIDTH(1)) andOp_16(.in0(andOp_16_in0), .in1(andOp_16_in1), .out(andOp_16_out));

	wire [0:0] notOp_17_in0;
	wire [0:0] notOp_17_out;
	notOp #(.WIDTH(1)) notOp_17(.in(notOp_17_in0), .out(notOp_17_out));

	wire [0:0] andOp_18_in0;
	wire [0:0] andOp_18_in1;
	wire [0:0] andOp_18_out;
	andOp #(.WIDTH(1)) andOp_18(.in0(andOp_18_in0), .in1(andOp_18_in1), .out(andOp_18_out));

	wire [0:0] andOp_19_in0;
	wire [0:0] andOp_19_in1;
	wire [0:0] andOp_19_out;
	andOp #(.WIDTH(1)) andOp_19(.in0(andOp_19_in0), .in1(andOp_19_in1), .out(andOp_19_out));

	wire [0:0] notOp_20_in0;
	wire [0:0] notOp_20_out;
	notOp #(.WIDTH(1)) notOp_20(.in(notOp_20_in0), .out(notOp_20_out));

	wire [0:0] andOp_21_in0;
	wire [0:0] andOp_21_in1;
	wire [0:0] andOp_21_out;
	andOp #(.WIDTH(1)) andOp_21(.in0(andOp_21_in0), .in1(andOp_21_in1), .out(andOp_21_out));

	wire [0:0] notOp_22_in0;
	wire [0:0] notOp_22_out;
	notOp #(.WIDTH(1)) notOp_22(.in(notOp_22_in0), .out(notOp_22_out));

	wire [0:0] andOp_23_in0;
	wire [0:0] andOp_23_in1;
	wire [0:0] andOp_23_out;
	andOp #(.WIDTH(1)) andOp_23(.in0(andOp_23_in0), .in1(andOp_23_in1), .out(andOp_23_out));

	wire [0:0] andOp_24_in0;
	wire [0:0] andOp_24_in1;
	wire [0:0] andOp_24_out;
	andOp #(.WIDTH(1)) andOp_24(.in0(andOp_24_in0), .in1(andOp_24_in1), .out(andOp_24_out));

	wire [0:0] notOp_25_in0;
	wire [0:0] notOp_25_out;
	notOp #(.WIDTH(1)) notOp_25(.in(notOp_25_in0), .out(notOp_25_out));

	wire [0:0] andOp_26_in0;
	wire [0:0] andOp_26_in1;
	wire [0:0] andOp_26_out;
	andOp #(.WIDTH(1)) andOp_26(.in0(andOp_26_in0), .in1(andOp_26_in1), .out(andOp_26_out));

	wire [0:0] notOp_27_in0;
	wire [0:0] notOp_27_out;
	notOp #(.WIDTH(1)) notOp_27(.in(notOp_27_in0), .out(notOp_27_out));

	wire [0:0] andOp_28_in0;
	wire [0:0] andOp_28_in1;
	wire [0:0] andOp_28_out;
	andOp #(.WIDTH(1)) andOp_28(.in0(andOp_28_in0), .in1(andOp_28_in1), .out(andOp_28_out));

	wire [0:0] andOp_29_in0;
	wire [0:0] andOp_29_in1;
	wire [0:0] andOp_29_out;
	andOp #(.WIDTH(1)) andOp_29(.in0(andOp_29_in0), .in1(andOp_29_in1), .out(andOp_29_out));

	wire [0:0] notOp_30_in0;
	wire [0:0] notOp_30_out;
	notOp #(.WIDTH(1)) notOp_30(.in(notOp_30_in0), .out(notOp_30_out));

	wire [0:0] andOp_31_in0;
	wire [0:0] andOp_31_in1;
	wire [0:0] andOp_31_out;
	andOp #(.WIDTH(1)) andOp_31(.in0(andOp_31_in0), .in1(andOp_31_in1), .out(andOp_31_out));

	wire [0:0] notOp_32_in0;
	wire [0:0] notOp_32_out;
	notOp #(.WIDTH(1)) notOp_32(.in(notOp_32_in0), .out(notOp_32_out));

	wire [0:0] andOp_33_in0;
	wire [0:0] andOp_33_in1;
	wire [0:0] andOp_33_out;
	andOp #(.WIDTH(1)) andOp_33(.in0(andOp_33_in0), .in1(andOp_33_in1), .out(andOp_33_out));

	wire [0:0] andOp_34_in0;
	wire [0:0] andOp_34_in1;
	wire [0:0] andOp_34_out;
	andOp #(.WIDTH(1)) andOp_34(.in0(andOp_34_in0), .in1(andOp_34_in1), .out(andOp_34_out));

	wire [0:0] notOp_35_in0;
	wire [0:0] notOp_35_out;
	notOp #(.WIDTH(1)) notOp_35(.in(notOp_35_in0), .out(notOp_35_out));

	wire [0:0] andOp_36_in0;
	wire [0:0] andOp_36_in1;
	wire [0:0] andOp_36_out;
	andOp #(.WIDTH(1)) andOp_36(.in0(andOp_36_in0), .in1(andOp_36_in1), .out(andOp_36_out));

	wire [0:0] notOp_37_in0;
	wire [0:0] notOp_37_out;
	notOp #(.WIDTH(1)) notOp_37(.in(notOp_37_in0), .out(notOp_37_out));

	wire [0:0] andOp_38_in0;
	wire [0:0] andOp_38_in1;
	wire [0:0] andOp_38_out;
	andOp #(.WIDTH(1)) andOp_38(.in0(andOp_38_in0), .in1(andOp_38_in1), .out(andOp_38_out));

	wire [0:0] andOp_39_in0;
	wire [0:0] andOp_39_in1;
	wire [0:0] andOp_39_out;
	andOp #(.WIDTH(1)) andOp_39(.in0(andOp_39_in0), .in1(andOp_39_in1), .out(andOp_39_out));

	wire [0:0] notOp_40_in0;
	wire [0:0] notOp_40_out;
	notOp #(.WIDTH(1)) notOp_40(.in(notOp_40_in0), .out(notOp_40_out));

	wire [0:0] andOp_41_in0;
	wire [0:0] andOp_41_in1;
	wire [0:0] andOp_41_out;
	andOp #(.WIDTH(1)) andOp_41(.in0(andOp_41_in0), .in1(andOp_41_in1), .out(andOp_41_out));

	wire [0:0] notOp_42_in0;
	wire [0:0] notOp_42_out;
	notOp #(.WIDTH(1)) notOp_42(.in(notOp_42_in0), .out(notOp_42_out));

	wire [0:0] andOp_43_in0;
	wire [0:0] andOp_43_in1;
	wire [0:0] andOp_43_out;
	andOp #(.WIDTH(1)) andOp_43(.in0(andOp_43_in0), .in1(andOp_43_in1), .out(andOp_43_out));

	wire [31:0] eq_44_in0;
	wire [31:0] eq_44_in1;
	wire [0:0] eq_44_out;
	eq #(.WIDTH(32)) eq_44(.in0(eq_44_in0), .in1(eq_44_in1), .out(eq_44_out));

	wire [31:0] eq_45_in0;
	wire [31:0] eq_45_in1;
	wire [0:0] eq_45_out;
	eq #(.WIDTH(32)) eq_45(.in0(eq_45_in0), .in1(eq_45_in1), .out(eq_45_out));

	wire [31:0] eq_46_in0;
	wire [31:0] eq_46_in1;
	wire [0:0] eq_46_out;
	eq #(.WIDTH(32)) eq_46(.in0(eq_46_in0), .in1(eq_46_in1), .out(eq_46_out));

	wire [31:0] eq_47_in0;
	wire [31:0] eq_47_in1;
	wire [0:0] eq_47_out;
	eq #(.WIDTH(32)) eq_47(.in0(eq_47_in0), .in1(eq_47_in1), .out(eq_47_out));

	wire [31:0] eq_48_in0;
	wire [31:0] eq_48_in1;
	wire [0:0] eq_48_out;
	eq #(.WIDTH(32)) eq_48(.in0(eq_48_in0), .in1(eq_48_in1), .out(eq_48_out));

	wire [31:0] eq_49_in0;
	wire [31:0] eq_49_in1;
	wire [0:0] eq_49_out;
	eq #(.WIDTH(32)) eq_49(.in0(eq_49_in0), .in1(eq_49_in1), .out(eq_49_out));

	wire [31:0] eq_50_in0;
	wire [31:0] eq_50_in1;
	wire [0:0] eq_50_out;
	eq #(.WIDTH(32)) eq_50(.in0(eq_50_in0), .in1(eq_50_in1), .out(eq_50_out));

	wire [31:0] eq_51_in0;
	wire [31:0] eq_51_in1;
	wire [0:0] eq_51_out;
	eq #(.WIDTH(32)) eq_51(.in0(eq_51_in0), .in1(eq_51_in1), .out(eq_51_out));

	wire [31:0] eq_52_in0;
	wire [31:0] eq_52_in1;
	wire [0:0] eq_52_out;
	eq #(.WIDTH(32)) eq_52(.in0(eq_52_in0), .in1(eq_52_in1), .out(eq_52_out));

	wire [31:0] eq_53_in0;
	wire [31:0] eq_53_in1;
	wire [0:0] eq_53_out;
	eq #(.WIDTH(32)) eq_53(.in0(eq_53_in0), .in1(eq_53_in1), .out(eq_53_out));

	wire [31:0] eq_54_in0;
	wire [31:0] eq_54_in1;
	wire [0:0] eq_54_out;
	eq #(.WIDTH(32)) eq_54(.in0(eq_54_in0), .in1(eq_54_in1), .out(eq_54_out));

	wire [31:0] eq_55_in0;
	wire [31:0] eq_55_in1;
	wire [0:0] eq_55_out;
	eq #(.WIDTH(32)) eq_55(.in0(eq_55_in0), .in1(eq_55_in1), .out(eq_55_out));

	wire [31:0] eq_56_in0;
	wire [31:0] eq_56_in1;
	wire [0:0] eq_56_out;
	eq #(.WIDTH(32)) eq_56(.in0(eq_56_in0), .in1(eq_56_in1), .out(eq_56_out));

	wire [31:0] eq_57_in0;
	wire [31:0] eq_57_in1;
	wire [0:0] eq_57_out;
	eq #(.WIDTH(32)) eq_57(.in0(eq_57_in0), .in1(eq_57_in1), .out(eq_57_out));

	wire [31:0] eq_58_in0;
	wire [31:0] eq_58_in1;
	wire [0:0] eq_58_out;
	eq #(.WIDTH(32)) eq_58(.in0(eq_58_in0), .in1(eq_58_in1), .out(eq_58_out));

	wire [31:0] eq_59_in0;
	wire [31:0] eq_59_in1;
	wire [0:0] eq_59_out;
	eq #(.WIDTH(32)) eq_59(.in0(eq_59_in0), .in1(eq_59_in1), .out(eq_59_out));

	wire [0:0] andOp_60_in0;
	wire [0:0] andOp_60_in1;
	wire [0:0] andOp_60_out;
	andOp #(.WIDTH(1)) andOp_60(.in0(andOp_60_in0), .in1(andOp_60_in1), .out(andOp_60_out));

	wire [31:0] concat_61_in0;
	wire [31:0] concat_61_in1;
	wire [63:0] concat_61_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_61(.in0(concat_61_in0), .in1(concat_61_in1), .out(concat_61_out));

	wire [31:0] concat_62_in0;
	wire [31:0] concat_62_in1;
	wire [63:0] concat_62_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_62(.in0(concat_62_in0), .in1(concat_62_in1), .out(concat_62_out));

	wire [0:0] andOp_63_in0;
	wire [0:0] andOp_63_in1;
	wire [0:0] andOp_63_out;
	andOp #(.WIDTH(1)) andOp_63(.in0(andOp_63_in0), .in1(andOp_63_in1), .out(andOp_63_out));

	wire [0:0] andOp_64_in0;
	wire [0:0] andOp_64_in1;
	wire [0:0] andOp_64_out;
	andOp #(.WIDTH(1)) andOp_64(.in0(andOp_64_in0), .in1(andOp_64_in1), .out(andOp_64_out));

	wire [0:0] andOp_65_in0;
	wire [0:0] andOp_65_in1;
	wire [0:0] andOp_65_out;
	andOp #(.WIDTH(1)) andOp_65(.in0(andOp_65_in0), .in1(andOp_65_in1), .out(andOp_65_out));

	wire [0:0] andOp_66_in0;
	wire [0:0] andOp_66_in1;
	wire [0:0] andOp_66_out;
	andOp #(.WIDTH(1)) andOp_66(.in0(andOp_66_in0), .in1(andOp_66_in1), .out(andOp_66_out));

	wire [0:0] andOp_67_in0;
	wire [0:0] andOp_67_in1;
	wire [0:0] andOp_67_out;
	andOp #(.WIDTH(1)) andOp_67(.in0(andOp_67_in0), .in1(andOp_67_in1), .out(andOp_67_out));

	wire [0:0] andOp_68_in0;
	wire [0:0] andOp_68_in1;
	wire [0:0] andOp_68_out;
	andOp #(.WIDTH(1)) andOp_68(.in0(andOp_68_in0), .in1(andOp_68_in1), .out(andOp_68_out));

	wire [0:0] andOp_69_in0;
	wire [0:0] andOp_69_in1;
	wire [0:0] andOp_69_out;
	andOp #(.WIDTH(1)) andOp_69(.in0(andOp_69_in0), .in1(andOp_69_in1), .out(andOp_69_out));

	wire [0:0] andOp_70_in0;
	wire [0:0] andOp_70_in1;
	wire [0:0] andOp_70_out;
	andOp #(.WIDTH(1)) andOp_70(.in0(andOp_70_in0), .in1(andOp_70_in1), .out(andOp_70_out));

	wire [0:0] andOp_71_in0;
	wire [0:0] andOp_71_in1;
	wire [0:0] andOp_71_out;
	andOp #(.WIDTH(1)) andOp_71(.in0(andOp_71_in0), .in1(andOp_71_in1), .out(andOp_71_out));

	wire [0:0] andOp_72_in0;
	wire [0:0] andOp_72_in1;
	wire [0:0] andOp_72_out;
	andOp #(.WIDTH(1)) andOp_72(.in0(andOp_72_in0), .in1(andOp_72_in1), .out(andOp_72_out));

	wire [0:0] andOp_73_in0;
	wire [0:0] andOp_73_in1;
	wire [0:0] andOp_73_out;
	andOp #(.WIDTH(1)) andOp_73(.in0(andOp_73_in0), .in1(andOp_73_in1), .out(andOp_73_out));

	wire [0:0] notOp_74_in0;
	wire [0:0] notOp_74_out;
	notOp #(.WIDTH(1)) notOp_74(.in(notOp_74_in0), .out(notOp_74_out));

	wire [0:0] andOp_75_in0;
	wire [0:0] andOp_75_in1;
	wire [0:0] andOp_75_out;
	andOp #(.WIDTH(1)) andOp_75(.in0(andOp_75_in0), .in1(andOp_75_in1), .out(andOp_75_out));

	wire [0:0] notOp_76_in0;
	wire [0:0] notOp_76_out;
	notOp #(.WIDTH(1)) notOp_76(.in(notOp_76_in0), .out(notOp_76_out));

	wire [0:0] andOp_77_in0;
	wire [0:0] andOp_77_in1;
	wire [0:0] andOp_77_out;
	andOp #(.WIDTH(1)) andOp_77(.in0(andOp_77_in0), .in1(andOp_77_in1), .out(andOp_77_out));

	wire [0:0] notOp_78_in0;
	wire [0:0] notOp_78_out;
	notOp #(.WIDTH(1)) notOp_78(.in(notOp_78_in0), .out(notOp_78_out));

	wire [0:0] andOp_79_in0;
	wire [0:0] andOp_79_in1;
	wire [0:0] andOp_79_out;
	andOp #(.WIDTH(1)) andOp_79(.in0(andOp_79_in0), .in1(andOp_79_in1), .out(andOp_79_out));

	wire [0:0] notOp_80_in0;
	wire [0:0] notOp_80_out;
	notOp #(.WIDTH(1)) notOp_80(.in(notOp_80_in0), .out(notOp_80_out));

	wire [0:0] andOp_81_in0;
	wire [0:0] andOp_81_in1;
	wire [0:0] andOp_81_out;
	andOp #(.WIDTH(1)) andOp_81(.in0(andOp_81_in0), .in1(andOp_81_in1), .out(andOp_81_out));

	wire [0:0] notOp_82_in0;
	wire [0:0] notOp_82_out;
	notOp #(.WIDTH(1)) notOp_82(.in(notOp_82_in0), .out(notOp_82_out));

	wire [0:0] andOp_83_in0;
	wire [0:0] andOp_83_in1;
	wire [0:0] andOp_83_out;
	andOp #(.WIDTH(1)) andOp_83(.in0(andOp_83_in0), .in1(andOp_83_in1), .out(andOp_83_out));

	wire [0:0] andOp_84_in0;
	wire [0:0] andOp_84_in1;
	wire [0:0] andOp_84_out;
	andOp #(.WIDTH(1)) andOp_84(.in0(andOp_84_in0), .in1(andOp_84_in1), .out(andOp_84_out));

	wire [0:0] andOp_85_in0;
	wire [0:0] andOp_85_in1;
	wire [0:0] andOp_85_out;
	andOp #(.WIDTH(1)) andOp_85(.in0(andOp_85_in0), .in1(andOp_85_in1), .out(andOp_85_out));

	wire [0:0] andOp_86_in0;
	wire [0:0] andOp_86_in1;
	wire [0:0] andOp_86_out;
	andOp #(.WIDTH(1)) andOp_86(.in0(andOp_86_in0), .in1(andOp_86_in1), .out(andOp_86_out));

	wire [0:0] notOp_87_in0;
	wire [0:0] notOp_87_out;
	notOp #(.WIDTH(1)) notOp_87(.in(notOp_87_in0), .out(notOp_87_out));

	wire [0:0] andOp_88_in0;
	wire [0:0] andOp_88_in1;
	wire [0:0] andOp_88_out;
	andOp #(.WIDTH(1)) andOp_88(.in0(andOp_88_in0), .in1(andOp_88_in1), .out(andOp_88_out));

	wire [0:0] notOp_89_in0;
	wire [0:0] notOp_89_out;
	notOp #(.WIDTH(1)) notOp_89(.in(notOp_89_in0), .out(notOp_89_out));

	wire [0:0] andOp_90_in0;
	wire [0:0] andOp_90_in1;
	wire [0:0] andOp_90_out;
	andOp #(.WIDTH(1)) andOp_90(.in0(andOp_90_in0), .in1(andOp_90_in1), .out(andOp_90_out));

	wire [0:0] notOp_91_in0;
	wire [0:0] notOp_91_out;
	notOp #(.WIDTH(1)) notOp_91(.in(notOp_91_in0), .out(notOp_91_out));

	wire [0:0] andOp_92_in0;
	wire [0:0] andOp_92_in1;
	wire [0:0] andOp_92_out;
	andOp #(.WIDTH(1)) andOp_92(.in0(andOp_92_in0), .in1(andOp_92_in1), .out(andOp_92_out));

	wire [0:0] notOp_93_in0;
	wire [0:0] notOp_93_out;
	notOp #(.WIDTH(1)) notOp_93(.in(notOp_93_in0), .out(notOp_93_out));

	wire [0:0] andOp_94_in0;
	wire [0:0] andOp_94_in1;
	wire [0:0] andOp_94_out;
	andOp #(.WIDTH(1)) andOp_94(.in0(andOp_94_in0), .in1(andOp_94_in1), .out(andOp_94_out));

	wire [0:0] notOp_95_in0;
	wire [0:0] notOp_95_out;
	notOp #(.WIDTH(1)) notOp_95(.in(notOp_95_in0), .out(notOp_95_out));

	wire [0:0] andOp_96_in0;
	wire [0:0] andOp_96_in1;
	wire [0:0] andOp_96_out;
	andOp #(.WIDTH(1)) andOp_96(.in0(andOp_96_in0), .in1(andOp_96_in1), .out(andOp_96_out));

	wire [0:0] andOp_97_in0;
	wire [0:0] andOp_97_in1;
	wire [0:0] andOp_97_out;
	andOp #(.WIDTH(1)) andOp_97(.in0(andOp_97_in0), .in1(andOp_97_in1), .out(andOp_97_out));

	wire [0:0] andOp_98_in0;
	wire [0:0] andOp_98_in1;
	wire [0:0] andOp_98_out;
	andOp #(.WIDTH(1)) andOp_98(.in0(andOp_98_in0), .in1(andOp_98_in1), .out(andOp_98_out));

	wire [31:0] add_100_in0;
	wire [31:0] add_100_in1;
	wire [31:0] add_100_out;
	add #(.WIDTH(32)) add_100(.in0(add_100_in0), .in1(add_100_in1), .out(add_100_out));

	wire [0:0] notOp_101_in0;
	wire [0:0] notOp_101_out;
	notOp #(.WIDTH(1)) notOp_101(.in(notOp_101_in0), .out(notOp_101_out));

	wire [0:0] andOp_102_in0;
	wire [0:0] andOp_102_in1;
	wire [0:0] andOp_102_out;
	andOp #(.WIDTH(1)) andOp_102(.in0(andOp_102_in0), .in1(andOp_102_in1), .out(andOp_102_out));

	wire [31:0] eq_103_in0;
	wire [31:0] eq_103_in1;
	wire [0:0] eq_103_out;
	eq #(.WIDTH(32)) eq_103(.in0(eq_103_in0), .in1(eq_103_in1), .out(eq_103_out));

	wire [0:0] andOp_105_in0;
	wire [0:0] andOp_105_in1;
	wire [0:0] andOp_105_out;
	andOp #(.WIDTH(1)) andOp_105(.in0(andOp_105_in0), .in1(andOp_105_in1), .out(andOp_105_out));

	wire [0:0] andOp_106_in0;
	wire [0:0] andOp_106_in1;
	wire [0:0] andOp_106_out;
	andOp #(.WIDTH(1)) andOp_106(.in0(andOp_106_in0), .in1(andOp_106_in1), .out(andOp_106_out));

	wire [0:0] andOp_107_in0;
	wire [0:0] andOp_107_in1;
	wire [0:0] andOp_107_out;
	andOp #(.WIDTH(1)) andOp_107(.in0(andOp_107_in0), .in1(andOp_107_in1), .out(andOp_107_out));

	wire [0:0] andOp_108_in0;
	wire [0:0] andOp_108_in1;
	wire [0:0] andOp_108_out;
	andOp #(.WIDTH(1)) andOp_108(.in0(andOp_108_in0), .in1(andOp_108_in1), .out(andOp_108_out));

	wire [0:0] andOp_109_in0;
	wire [0:0] andOp_109_in1;
	wire [0:0] andOp_109_out;
	andOp #(.WIDTH(1)) andOp_109(.in0(andOp_109_in0), .in1(andOp_109_in1), .out(andOp_109_out));

	wire [0:0] andOp_110_in0;
	wire [0:0] andOp_110_in1;
	wire [0:0] andOp_110_out;
	andOp #(.WIDTH(1)) andOp_110(.in0(andOp_110_in0), .in1(andOp_110_in1), .out(andOp_110_out));

	wire [0:0] andOp_111_in0;
	wire [0:0] andOp_111_in1;
	wire [0:0] andOp_111_out;
	andOp #(.WIDTH(1)) andOp_111(.in0(andOp_111_in0), .in1(andOp_111_in1), .out(andOp_111_out));

	wire [0:0] notOp_112_in0;
	wire [0:0] notOp_112_out;
	notOp #(.WIDTH(1)) notOp_112(.in(notOp_112_in0), .out(notOp_112_out));

	wire [0:0] andOp_113_in0;
	wire [0:0] andOp_113_in1;
	wire [0:0] andOp_113_out;
	andOp #(.WIDTH(1)) andOp_113(.in0(andOp_113_in0), .in1(andOp_113_in1), .out(andOp_113_out));

	wire [0:0] notOp_114_in0;
	wire [0:0] notOp_114_out;
	notOp #(.WIDTH(1)) notOp_114(.in(notOp_114_in0), .out(notOp_114_out));

	wire [0:0] andOp_115_in0;
	wire [0:0] andOp_115_in1;
	wire [0:0] andOp_115_out;
	andOp #(.WIDTH(1)) andOp_115(.in0(andOp_115_in0), .in1(andOp_115_in1), .out(andOp_115_out));

	wire [0:0] notOp_116_in0;
	wire [0:0] notOp_116_out;
	notOp #(.WIDTH(1)) notOp_116(.in(notOp_116_in0), .out(notOp_116_out));

	wire [0:0] andOp_117_in0;
	wire [0:0] andOp_117_in1;
	wire [0:0] andOp_117_out;
	andOp #(.WIDTH(1)) andOp_117(.in0(andOp_117_in0), .in1(andOp_117_in1), .out(andOp_117_out));

	wire [0:0] notOp_118_in0;
	wire [0:0] notOp_118_out;
	notOp #(.WIDTH(1)) notOp_118(.in(notOp_118_in0), .out(notOp_118_out));

	wire [0:0] andOp_119_in0;
	wire [0:0] andOp_119_in1;
	wire [0:0] andOp_119_out;
	andOp #(.WIDTH(1)) andOp_119(.in0(andOp_119_in0), .in1(andOp_119_in1), .out(andOp_119_out));

	wire [0:0] notOp_120_in0;
	wire [0:0] notOp_120_out;
	notOp #(.WIDTH(1)) notOp_120(.in(notOp_120_in0), .out(notOp_120_out));

	wire [0:0] andOp_121_in0;
	wire [0:0] andOp_121_in1;
	wire [0:0] andOp_121_out;
	andOp #(.WIDTH(1)) andOp_121(.in0(andOp_121_in0), .in1(andOp_121_in1), .out(andOp_121_out));

	wire [0:0] notOp_122_in0;
	wire [0:0] notOp_122_out;
	notOp #(.WIDTH(1)) notOp_122(.in(notOp_122_in0), .out(notOp_122_out));

	wire [0:0] andOp_123_in0;
	wire [0:0] andOp_123_in1;
	wire [0:0] andOp_123_out;
	andOp #(.WIDTH(1)) andOp_123(.in0(andOp_123_in0), .in1(andOp_123_in1), .out(andOp_123_out));

	wire [0:0] notOp_124_in0;
	wire [0:0] notOp_124_out;
	notOp #(.WIDTH(1)) notOp_124(.in(notOp_124_in0), .out(notOp_124_out));

	wire [0:0] andOp_125_in0;
	wire [0:0] andOp_125_in1;
	wire [0:0] andOp_125_out;
	andOp #(.WIDTH(1)) andOp_125(.in0(andOp_125_in0), .in1(andOp_125_in1), .out(andOp_125_out));

	wire [0:0] notOp_126_in0;
	wire [0:0] notOp_126_out;
	notOp #(.WIDTH(1)) notOp_126(.in(notOp_126_in0), .out(notOp_126_out));

	wire [0:0] andOp_127_in0;
	wire [0:0] andOp_127_in1;
	wire [0:0] andOp_127_out;
	andOp #(.WIDTH(1)) andOp_127(.in0(andOp_127_in0), .in1(andOp_127_in1), .out(andOp_127_out));

	wire [0:0] notOp_128_in0;
	wire [0:0] notOp_128_out;
	notOp #(.WIDTH(1)) notOp_128(.in(notOp_128_in0), .out(notOp_128_out));

	wire [0:0] andOp_129_in0;
	wire [0:0] andOp_129_in1;
	wire [0:0] andOp_129_out;
	andOp #(.WIDTH(1)) andOp_129(.in0(andOp_129_in0), .in1(andOp_129_in1), .out(andOp_129_out));

	reg [0:0] in_pipeline_0_in_data;
	wire [0:0] in_pipeline_0_out_data;
	hls_wire #(.WIDTH(1)) in_pipeline_0(.in_data(in_pipeline_0_in_data), .out_data(in_pipeline_0_out_data));

	wire [0:0] orOp_130_in0;
	wire [0:0] orOp_130_in1;
	wire [0:0] orOp_130_out;
	orOp #(.WIDTH(1)) orOp_130(.in0(orOp_130_in0), .in1(orOp_130_in1), .out(orOp_130_out));

	wire [0:0] orOp_131_in0;
	wire [0:0] orOp_131_in1;
	wire [0:0] orOp_131_out;
	orOp #(.WIDTH(1)) orOp_131(.in0(orOp_131_in0), .in1(orOp_131_in1), .out(orOp_131_out));

	wire [0:0] orOp_132_in0;
	wire [0:0] orOp_132_in1;
	wire [0:0] orOp_132_out;
	orOp #(.WIDTH(1)) orOp_132(.in0(orOp_132_in0), .in1(orOp_132_in1), .out(orOp_132_out));

	wire [0:0] orOp_133_in0;
	wire [0:0] orOp_133_in1;
	wire [0:0] orOp_133_out;
	orOp #(.WIDTH(1)) orOp_133(.in0(orOp_133_in0), .in1(orOp_133_in1), .out(orOp_133_out));

	wire [0:0] orOp_134_in0;
	wire [0:0] orOp_134_in1;
	wire [0:0] orOp_134_out;
	orOp #(.WIDTH(1)) orOp_134(.in0(orOp_134_in0), .in1(orOp_134_in1), .out(orOp_134_out));

	wire [0:0] orOp_135_in0;
	wire [0:0] orOp_135_in1;
	wire [0:0] orOp_135_out;
	orOp #(.WIDTH(1)) orOp_135(.in0(orOp_135_in0), .in1(orOp_135_in1), .out(orOp_135_out));

	wire [31:0] eq_136_in0;
	wire [31:0] eq_136_in1;
	wire [0:0] eq_136_out;
	eq #(.WIDTH(32)) eq_136(.in0(eq_136_in0), .in1(eq_136_in1), .out(eq_136_out));

	wire [31:0] eq_137_in0;
	wire [31:0] eq_137_in1;
	wire [0:0] eq_137_out;
	eq #(.WIDTH(32)) eq_137(.in0(eq_137_in0), .in1(eq_137_in1), .out(eq_137_out));

	wire [31:0] eq_138_in0;
	wire [31:0] eq_138_in1;
	wire [0:0] eq_138_out;
	eq #(.WIDTH(32)) eq_138(.in0(eq_138_in0), .in1(eq_138_in1), .out(eq_138_out));

	wire [0:0] andOp_139_in0;
	wire [0:0] andOp_139_in1;
	wire [0:0] andOp_139_out;
	andOp #(.WIDTH(1)) andOp_139(.in0(andOp_139_in0), .in1(andOp_139_in1), .out(andOp_139_out));

	wire [0:0] andOp_140_in0;
	wire [0:0] andOp_140_in1;
	wire [0:0] andOp_140_out;
	andOp #(.WIDTH(1)) andOp_140(.in0(andOp_140_in0), .in1(andOp_140_in1), .out(andOp_140_out));

	wire [31:0] eq_141_in0;
	wire [31:0] eq_141_in1;
	wire [0:0] eq_141_out;
	eq #(.WIDTH(32)) eq_141(.in0(eq_141_in0), .in1(eq_141_in1), .out(eq_141_out));

	wire [31:0] eq_142_in0;
	wire [31:0] eq_142_in1;
	wire [0:0] eq_142_out;
	eq #(.WIDTH(32)) eq_142(.in0(eq_142_in0), .in1(eq_142_in1), .out(eq_142_out));

	wire [0:0] andOp_143_in0;
	wire [0:0] andOp_143_in1;
	wire [0:0] andOp_143_out;
	andOp #(.WIDTH(1)) andOp_143(.in0(andOp_143_in0), .in1(andOp_143_in1), .out(andOp_143_out));

	wire [0:0] andOp_144_in0;
	wire [0:0] andOp_144_in1;
	wire [0:0] andOp_144_out;
	andOp #(.WIDTH(1)) andOp_144(.in0(andOp_144_in0), .in1(andOp_144_in1), .out(andOp_144_out));

	wire [31:0] eq_145_in0;
	wire [31:0] eq_145_in1;
	wire [0:0] eq_145_out;
	eq #(.WIDTH(32)) eq_145(.in0(eq_145_in0), .in1(eq_145_in1), .out(eq_145_out));

	wire [31:0] eq_146_in0;
	wire [31:0] eq_146_in1;
	wire [0:0] eq_146_out;
	eq #(.WIDTH(32)) eq_146(.in0(eq_146_in0), .in1(eq_146_in1), .out(eq_146_out));

	wire [31:0] eq_147_in0;
	wire [31:0] eq_147_in1;
	wire [0:0] eq_147_out;
	eq #(.WIDTH(32)) eq_147(.in0(eq_147_in0), .in1(eq_147_in1), .out(eq_147_out));

	wire [31:0] eq_148_in0;
	wire [31:0] eq_148_in1;
	wire [0:0] eq_148_out;
	eq #(.WIDTH(32)) eq_148(.in0(eq_148_in0), .in1(eq_148_in1), .out(eq_148_out));

	wire [31:0] eq_149_in0;
	wire [31:0] eq_149_in1;
	wire [0:0] eq_149_out;
	eq #(.WIDTH(32)) eq_149(.in0(eq_149_in0), .in1(eq_149_in1), .out(eq_149_out));

	wire [31:0] eq_150_in0;
	wire [31:0] eq_150_in1;
	wire [0:0] eq_150_out;
	eq #(.WIDTH(32)) eq_150(.in0(eq_150_in0), .in1(eq_150_in1), .out(eq_150_out));

	wire [31:0] eq_151_in0;
	wire [31:0] eq_151_in1;
	wire [0:0] eq_151_out;
	eq #(.WIDTH(32)) eq_151(.in0(eq_151_in0), .in1(eq_151_in1), .out(eq_151_out));

	wire [31:0] eq_152_in0;
	wire [31:0] eq_152_in1;
	wire [0:0] eq_152_out;
	eq #(.WIDTH(32)) eq_152(.in0(eq_152_in0), .in1(eq_152_in1), .out(eq_152_out));

	wire [31:0] eq_153_in0;
	wire [31:0] eq_153_in1;
	wire [0:0] eq_153_out;
	eq #(.WIDTH(32)) eq_153(.in0(eq_153_in0), .in1(eq_153_in1), .out(eq_153_out));

	wire [31:0] eq_154_in0;
	wire [31:0] eq_154_in1;
	wire [0:0] eq_154_out;
	eq #(.WIDTH(32)) eq_154(.in0(eq_154_in0), .in1(eq_154_in1), .out(eq_154_out));

	wire [31:0] eq_155_in0;
	wire [31:0] eq_155_in1;
	wire [0:0] eq_155_out;
	eq #(.WIDTH(32)) eq_155(.in0(eq_155_in0), .in1(eq_155_in1), .out(eq_155_out));

	wire [0:0] notOp_156_in0;
	wire [0:0] notOp_156_out;
	notOp #(.WIDTH(1)) notOp_156(.in(notOp_156_in0), .out(notOp_156_out));

	wire [0:0] notOp_157_in0;
	wire [0:0] notOp_157_out;
	notOp #(.WIDTH(1)) notOp_157(.in(notOp_157_in0), .out(notOp_157_out));

	wire [0:0] andOp_158_in0;
	wire [0:0] andOp_158_in1;
	wire [0:0] andOp_158_out;
	andOp #(.WIDTH(1)) andOp_158(.in0(andOp_158_in0), .in1(andOp_158_in1), .out(andOp_158_out));

	wire [0:0] andOp_159_in0;
	wire [0:0] andOp_159_in1;
	wire [0:0] andOp_159_out;
	andOp #(.WIDTH(1)) andOp_159(.in0(andOp_159_in0), .in1(andOp_159_in1), .out(andOp_159_out));

	wire [0:0] andOp_160_in0;
	wire [0:0] andOp_160_in1;
	wire [0:0] andOp_160_out;
	andOp #(.WIDTH(1)) andOp_160(.in0(andOp_160_in0), .in1(andOp_160_in1), .out(andOp_160_out));

	wire [0:0] andOp_161_in0;
	wire [0:0] andOp_161_in1;
	wire [0:0] andOp_161_out;
	andOp #(.WIDTH(1)) andOp_161(.in0(andOp_161_in0), .in1(andOp_161_in1), .out(andOp_161_out));

	wire [0:0] andOp_162_in0;
	wire [0:0] andOp_162_in1;
	wire [0:0] andOp_162_out;
	andOp #(.WIDTH(1)) andOp_162(.in0(andOp_162_in0), .in1(andOp_162_in1), .out(andOp_162_out));

	wire [0:0] andOp_163_in0;
	wire [0:0] andOp_163_in1;
	wire [0:0] andOp_163_out;
	andOp #(.WIDTH(1)) andOp_163(.in0(andOp_163_in0), .in1(andOp_163_in1), .out(andOp_163_out));

	wire [0:0] andOp_164_in0;
	wire [0:0] andOp_164_in1;
	wire [0:0] andOp_164_out;
	andOp #(.WIDTH(1)) andOp_164(.in0(andOp_164_in0), .in1(andOp_164_in1), .out(andOp_164_out));

	// End Functional Units

	reg [31:0] counter__99;
	reg [31:0] data_store_0_0;
	reg [31:0] data_store_1_2;
	reg [31:0] data_store_1_3;
	reg [31:0] data_store_2_5;
	reg [31:0] data_store_2_7;
	reg [31:0] data_store_2_8;
	reg [0:0] delayed_signal__104;
	reg [31:0] global_state;
	reg [0:0] out_of_pipe_1_7;
	reg [0:0] out_of_pipe_bb_1_7;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_3_last_state;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;
	reg [31:0] state_4_last_state;
	reg [31:0] state_5_entry_BB_reg;
	reg [0:0] state_5_is_active;
	reg [31:0] state_5_last_BB_reg;
	reg [31:0] state_5_last_state;
	reg [31:0] state_6_entry_BB_reg;
	reg [0:0] state_6_is_active;
	reg [31:0] state_6_last_BB_reg;
	reg [31:0] state_6_last_state;
	reg [31:0] state_7_entry_BB_reg;
	reg [0:0] state_7_is_active;
	reg [31:0] state_7_last_BB_reg;
	reg [31:0] state_7_last_state;

	// controller for add_100.add_100_in0
	// controller for add_100.add_100_in1
	// Insensitive connections
	assign add_100_in0 = counter__99;
	assign add_100_in1 = 32'd1;
	// controller for add_add10.add_add10_in0
	// controller for add_add10.add_add10_in1
	// Insensitive connections
	assign add_add10_in0 = data_in_3_10_out_data;
	assign add_add10_in1 = mul_mul9_out;
	// controller for add_add2.add_add2_in0
	// controller for add_add2.add_add2_in1
	// Insensitive connections
	assign add_add2_in0 = phi_phi1_out;
	assign add_add2_in1 = 32'd1;
	// controller for andOp_102.andOp_102_in0
	// controller for andOp_102.andOp_102_in1
	// Insensitive connections
	assign andOp_102_in0 = notOp_101_out;
	assign andOp_102_in1 = 1'd1;
	// controller for andOp_105.andOp_105_in0
	// controller for andOp_105.andOp_105_in1
	// Insensitive connections
	assign andOp_105_in0 = delayed_signal__104;
	assign andOp_105_in1 = eq_103_out;
	// controller for andOp_106.andOp_106_in0
	// controller for andOp_106.andOp_106_in1
	// Insensitive connections
	assign andOp_106_in0 = bb_2_active_in_state_1_out_data;
	assign andOp_106_in1 = state_1_is_active;
	// controller for andOp_107.andOp_107_in0
	// controller for andOp_107.andOp_107_in1
	// Insensitive connections
	assign andOp_107_in0 = bb_2_active_in_state_2_out_data;
	assign andOp_107_in1 = state_2_is_active;
	// controller for andOp_108.andOp_108_in0
	// controller for andOp_108.andOp_108_in1
	// Insensitive connections
	assign andOp_108_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_108_in1 = state_3_is_active;
	// controller for andOp_109.andOp_109_in0
	// controller for andOp_109.andOp_109_in1
	// Insensitive connections
	assign andOp_109_in0 = bb_2_active_in_state_4_out_data;
	assign andOp_109_in1 = state_4_is_active;
	// controller for andOp_110.andOp_110_in0
	// controller for andOp_110.andOp_110_in1
	// Insensitive connections
	assign andOp_110_in0 = bb_2_active_in_state_5_out_data;
	assign andOp_110_in1 = state_5_is_active;
	// controller for andOp_111.andOp_111_in0
	// controller for andOp_111.andOp_111_in1
	// Insensitive connections
	assign andOp_111_in0 = bb_1_active_in_state_7_out_data;
	assign andOp_111_in1 = state_7_is_active;
	// controller for andOp_113.andOp_113_in0
	// controller for andOp_113.andOp_113_in1
	// Insensitive connections
	assign andOp_113_in0 = notOp_112_out;
	assign andOp_113_in1 = 1'd1;
	// controller for andOp_115.andOp_115_in0
	// controller for andOp_115.andOp_115_in1
	// Insensitive connections
	assign andOp_115_in0 = notOp_114_out;
	assign andOp_115_in1 = andOp_113_out;
	// controller for andOp_117.andOp_117_in0
	// controller for andOp_117.andOp_117_in1
	// Insensitive connections
	assign andOp_117_in0 = notOp_116_out;
	assign andOp_117_in1 = 1'd1;
	// controller for andOp_119.andOp_119_in0
	// controller for andOp_119.andOp_119_in1
	// Insensitive connections
	assign andOp_119_in0 = notOp_118_out;
	assign andOp_119_in1 = 1'd1;
	// controller for andOp_12.andOp_12_in0
	// controller for andOp_12.andOp_12_in1
	// Insensitive connections
	assign andOp_12_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_12_in1 = state_0_is_active;
	// controller for andOp_121.andOp_121_in0
	// controller for andOp_121.andOp_121_in1
	// Insensitive connections
	assign andOp_121_in0 = notOp_120_out;
	assign andOp_121_in1 = 1'd1;
	// controller for andOp_123.andOp_123_in0
	// controller for andOp_123.andOp_123_in1
	// Insensitive connections
	assign andOp_123_in0 = notOp_122_out;
	assign andOp_123_in1 = 1'd1;
	// controller for andOp_125.andOp_125_in0
	// controller for andOp_125.andOp_125_in1
	// Insensitive connections
	assign andOp_125_in0 = notOp_124_out;
	assign andOp_125_in1 = 1'd1;
	// controller for andOp_127.andOp_127_in0
	// controller for andOp_127.andOp_127_in1
	// Insensitive connections
	assign andOp_127_in0 = notOp_126_out;
	assign andOp_127_in1 = 1'd1;
	// controller for andOp_129.andOp_129_in0
	// controller for andOp_129.andOp_129_in1
	// Insensitive connections
	assign andOp_129_in0 = notOp_128_out;
	assign andOp_129_in1 = andOp_127_out;
	// controller for andOp_139.andOp_139_in0
	// controller for andOp_139.andOp_139_in1
	// Insensitive connections
	assign andOp_139_in0 = bb_2_active_in_state_1_out_data;
	assign andOp_139_in1 = state_1_is_active;
	// controller for andOp_14.andOp_14_in0
	// controller for andOp_14.andOp_14_in1
	// Insensitive connections
	assign andOp_14_in0 = bb_2_active_in_state_1_out_data;
	assign andOp_14_in1 = state_1_is_active;
	// controller for andOp_140.andOp_140_in0
	// controller for andOp_140.andOp_140_in1
	// Insensitive connections
	assign andOp_140_in0 = bb_2_active_in_state_1_out_data;
	assign andOp_140_in1 = state_1_is_active;
	// controller for andOp_143.andOp_143_in0
	// controller for andOp_143.andOp_143_in1
	// Insensitive connections
	assign andOp_143_in0 = bb_2_active_in_state_2_out_data;
	assign andOp_143_in1 = state_2_is_active;
	// controller for andOp_144.andOp_144_in0
	// controller for andOp_144.andOp_144_in1
	// Insensitive connections
	assign andOp_144_in0 = bb_2_active_in_state_2_out_data;
	assign andOp_144_in1 = state_2_is_active;
	// controller for andOp_158.andOp_158_in0
	// controller for andOp_158.andOp_158_in1
	// Insensitive connections
	assign andOp_158_in0 = bb_2_active_in_state_1_out_data;
	assign andOp_158_in1 = state_1_is_active;
	// controller for andOp_159.andOp_159_in0
	// controller for andOp_159.andOp_159_in1
	// Insensitive connections
	assign andOp_159_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_159_in1 = state_3_is_active;
	// controller for andOp_16.andOp_16_in0
	// controller for andOp_16.andOp_16_in1
	// Insensitive connections
	assign andOp_16_in0 = andOp_14_out;
	assign andOp_16_in1 = icmp_icmp3_out;
	// controller for andOp_160.andOp_160_in0
	// controller for andOp_160.andOp_160_in1
	// Insensitive connections
	assign andOp_160_in0 = bb_2_active_in_state_2_out_data;
	assign andOp_160_in1 = state_2_is_active;
	// controller for andOp_161.andOp_161_in0
	// controller for andOp_161.andOp_161_in1
	// Insensitive connections
	assign andOp_161_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_161_in1 = state_3_is_active;
	// controller for andOp_162.andOp_162_in0
	// controller for andOp_162.andOp_162_in1
	// Insensitive connections
	assign andOp_162_in0 = bb_2_active_in_state_1_out_data;
	assign andOp_162_in1 = state_1_is_active;
	// controller for andOp_163.andOp_163_in0
	// controller for andOp_163.andOp_163_in1
	// Insensitive connections
	assign andOp_163_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_163_in1 = state_3_is_active;
	// controller for andOp_164.andOp_164_in0
	// controller for andOp_164.andOp_164_in1
	// Insensitive connections
	assign andOp_164_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_164_in1 = state_3_is_active;
	// controller for andOp_18.andOp_18_in0
	// controller for andOp_18.andOp_18_in1
	// Insensitive connections
	assign andOp_18_in0 = andOp_14_out;
	assign andOp_18_in1 = notOp_17_out;
	// controller for andOp_19.andOp_19_in0
	// controller for andOp_19.andOp_19_in1
	// Insensitive connections
	assign andOp_19_in0 = bb_2_active_in_state_1_out_data;
	assign andOp_19_in1 = state_1_is_active;
	// controller for andOp_21.andOp_21_in0
	// controller for andOp_21.andOp_21_in1
	// Insensitive connections
	assign andOp_21_in0 = andOp_19_out;
	assign andOp_21_in1 = icmp_icmp3_out;
	// controller for andOp_23.andOp_23_in0
	// controller for andOp_23.andOp_23_in1
	// Insensitive connections
	assign andOp_23_in0 = andOp_19_out;
	assign andOp_23_in1 = notOp_22_out;
	// controller for andOp_24.andOp_24_in0
	// controller for andOp_24.andOp_24_in1
	// Insensitive connections
	assign andOp_24_in0 = bb_2_active_in_state_1_out_data;
	assign andOp_24_in1 = state_1_is_active;
	// controller for andOp_26.andOp_26_in0
	// controller for andOp_26.andOp_26_in1
	// Insensitive connections
	assign andOp_26_in0 = andOp_24_out;
	assign andOp_26_in1 = icmp_icmp3_out;
	// controller for andOp_28.andOp_28_in0
	// controller for andOp_28.andOp_28_in1
	// Insensitive connections
	assign andOp_28_in0 = andOp_24_out;
	assign andOp_28_in1 = notOp_27_out;
	// controller for andOp_29.andOp_29_in0
	// controller for andOp_29.andOp_29_in1
	// Insensitive connections
	assign andOp_29_in0 = bb_2_active_in_state_1_out_data;
	assign andOp_29_in1 = state_1_is_active;
	// controller for andOp_31.andOp_31_in0
	// controller for andOp_31.andOp_31_in1
	// Insensitive connections
	assign andOp_31_in0 = andOp_29_out;
	assign andOp_31_in1 = icmp_icmp3_out;
	// controller for andOp_33.andOp_33_in0
	// controller for andOp_33.andOp_33_in1
	// Insensitive connections
	assign andOp_33_in0 = andOp_29_out;
	assign andOp_33_in1 = notOp_32_out;
	// controller for andOp_34.andOp_34_in0
	// controller for andOp_34.andOp_34_in1
	// Insensitive connections
	assign andOp_34_in0 = bb_2_active_in_state_1_out_data;
	assign andOp_34_in1 = state_1_is_active;
	// controller for andOp_36.andOp_36_in0
	// controller for andOp_36.andOp_36_in1
	// Insensitive connections
	assign andOp_36_in0 = andOp_34_out;
	assign andOp_36_in1 = icmp_icmp3_out;
	// controller for andOp_38.andOp_38_in0
	// controller for andOp_38.andOp_38_in1
	// Insensitive connections
	assign andOp_38_in0 = andOp_34_out;
	assign andOp_38_in1 = notOp_37_out;
	// controller for andOp_39.andOp_39_in0
	// controller for andOp_39.andOp_39_in1
	// Insensitive connections
	assign andOp_39_in0 = bb_2_active_in_state_1_out_data;
	assign andOp_39_in1 = state_1_is_active;
	// controller for andOp_41.andOp_41_in0
	// controller for andOp_41.andOp_41_in1
	// Insensitive connections
	assign andOp_41_in0 = andOp_39_out;
	assign andOp_41_in1 = icmp_icmp3_out;
	// controller for andOp_43.andOp_43_in0
	// controller for andOp_43.andOp_43_in1
	// Insensitive connections
	assign andOp_43_in0 = andOp_39_out;
	assign andOp_43_in1 = notOp_42_out;
	// controller for andOp_60.andOp_60_in0
	// controller for andOp_60.andOp_60_in1
	// Insensitive connections
	assign andOp_60_in0 = bb_2_active_in_state_1_out_data;
	assign andOp_60_in1 = state_1_is_active;
	// controller for andOp_63.andOp_63_in0
	// controller for andOp_63.andOp_63_in1
	// Insensitive connections
	assign andOp_63_in0 = bb_2_active_in_state_1_out_data;
	assign andOp_63_in1 = state_1_is_active;
	// controller for andOp_64.andOp_64_in0
	// controller for andOp_64.andOp_64_in1
	// Insensitive connections
	assign andOp_64_in0 = bb_2_active_in_state_1_out_data;
	assign andOp_64_in1 = state_1_is_active;
	// controller for andOp_65.andOp_65_in0
	// controller for andOp_65.andOp_65_in1
	// Insensitive connections
	assign andOp_65_in0 = bb_2_active_in_state_1_out_data;
	assign andOp_65_in1 = state_1_is_active;
	// controller for andOp_66.andOp_66_in0
	// controller for andOp_66.andOp_66_in1
	// Insensitive connections
	assign andOp_66_in0 = bb_2_active_in_state_2_out_data;
	assign andOp_66_in1 = state_2_is_active;
	// controller for andOp_67.andOp_67_in0
	// controller for andOp_67.andOp_67_in1
	// Insensitive connections
	assign andOp_67_in0 = bb_2_active_in_state_2_out_data;
	assign andOp_67_in1 = state_2_is_active;
	// controller for andOp_68.andOp_68_in0
	// controller for andOp_68.andOp_68_in1
	// Insensitive connections
	assign andOp_68_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_68_in1 = state_3_is_active;
	// controller for andOp_69.andOp_69_in0
	// controller for andOp_69.andOp_69_in1
	// Insensitive connections
	assign andOp_69_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_69_in1 = state_3_is_active;
	// controller for andOp_70.andOp_70_in0
	// controller for andOp_70.andOp_70_in1
	// Insensitive connections
	assign andOp_70_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_70_in1 = state_3_is_active;
	// controller for andOp_71.andOp_71_in0
	// controller for andOp_71.andOp_71_in1
	// Insensitive connections
	assign andOp_71_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_71_in1 = state_3_is_active;
	// controller for andOp_72.andOp_72_in0
	// controller for andOp_72.andOp_72_in1
	// Insensitive connections
	assign andOp_72_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_72_in1 = state_3_is_active;
	// controller for andOp_73.andOp_73_in0
	// controller for andOp_73.andOp_73_in1
	// Insensitive connections
	assign andOp_73_in0 = bb_1_active_in_state_7_out_data;
	assign andOp_73_in1 = state_7_is_active;
	// controller for andOp_75.andOp_75_in0
	// controller for andOp_75.andOp_75_in1
	// Insensitive connections
	assign andOp_75_in0 = 1'd1;
	assign andOp_75_in1 = notOp_74_out;
	// controller for andOp_77.andOp_77_in0
	// controller for andOp_77.andOp_77_in1
	// Insensitive connections
	assign andOp_77_in0 = andOp_75_out;
	assign andOp_77_in1 = notOp_76_out;
	// controller for andOp_79.andOp_79_in0
	// controller for andOp_79.andOp_79_in1
	// Insensitive connections
	assign andOp_79_in0 = andOp_77_out;
	assign andOp_79_in1 = notOp_78_out;
	// controller for andOp_81.andOp_81_in0
	// controller for andOp_81.andOp_81_in1
	// Insensitive connections
	assign andOp_81_in0 = andOp_79_out;
	assign andOp_81_in1 = notOp_80_out;
	// controller for andOp_83.andOp_83_in0
	// controller for andOp_83.andOp_83_in1
	// Insensitive connections
	assign andOp_83_in0 = andOp_81_out;
	assign andOp_83_in1 = notOp_82_out;
	// controller for andOp_84.andOp_84_in0
	// controller for andOp_84.andOp_84_in1
	// Insensitive connections
	assign andOp_84_in0 = in_pipeline_0_out_data;
	assign andOp_84_in1 = andOp_83_out;
	// controller for andOp_85.andOp_85_in0
	// controller for andOp_85.andOp_85_in1
	// Insensitive connections
	assign andOp_85_in0 = andOp_84_out;
	assign andOp_85_in1 = out_of_pipe_1_7;
	// controller for andOp_86.andOp_86_in0
	// controller for andOp_86.andOp_86_in1
	// Insensitive connections
	assign andOp_86_in0 = andOp_84_out;
	assign andOp_86_in1 = out_of_pipe_1_7;
	// controller for andOp_88.andOp_88_in0
	// controller for andOp_88.andOp_88_in1
	// Insensitive connections
	assign andOp_88_in0 = 1'd1;
	assign andOp_88_in1 = notOp_87_out;
	// controller for andOp_90.andOp_90_in0
	// controller for andOp_90.andOp_90_in1
	// Insensitive connections
	assign andOp_90_in0 = andOp_88_out;
	assign andOp_90_in1 = notOp_89_out;
	// controller for andOp_92.andOp_92_in0
	// controller for andOp_92.andOp_92_in1
	// Insensitive connections
	assign andOp_92_in0 = andOp_90_out;
	assign andOp_92_in1 = notOp_91_out;
	// controller for andOp_94.andOp_94_in0
	// controller for andOp_94.andOp_94_in1
	// Insensitive connections
	assign andOp_94_in0 = andOp_92_out;
	assign andOp_94_in1 = notOp_93_out;
	// controller for andOp_96.andOp_96_in0
	// controller for andOp_96.andOp_96_in1
	// Insensitive connections
	assign andOp_96_in0 = andOp_94_out;
	assign andOp_96_in1 = notOp_95_out;
	// controller for andOp_97.andOp_97_in0
	// controller for andOp_97.andOp_97_in1
	// Insensitive connections
	assign andOp_97_in0 = in_pipeline_0_out_data;
	assign andOp_97_in1 = andOp_96_out;
	// controller for andOp_98.andOp_98_in0
	// controller for andOp_98.andOp_98_in1
	// Insensitive connections
	assign andOp_98_in0 = andOp_97_out;
	assign andOp_98_in1 = out_of_pipe_bb_1_7;
	// controller for arg_0.arg_0_raddr_0_reg
	always @(*) begin
		if (andOp_65_out) begin 
			arg_0_raddr_0_reg = phi_phi1_out;
		end else begin
			arg_0_raddr_0_reg = 0;
		end
	end
	// controller for arg_1.arg_1_waddr_0_reg
	always @(*) begin
		if (andOp_68_out) begin 
			arg_1_waddr_0_reg = data_in_3_9_out_data;
		end else begin
			arg_1_waddr_0_reg = 0;
		end
	end
	// controller for arg_1.arg_1_wdata_0_reg
	always @(*) begin
		if (andOp_69_out) begin 
			arg_1_wdata_0_reg = add_add10_out;
		end else begin
			arg_1_wdata_0_reg = 0;
		end
	end
	// controller for arg_1.arg_1_wen_0_reg
	always @(*) begin
		if (andOp_70_out) begin 
			arg_1_wen_0_reg = -(1'd1);
		end else begin
			arg_1_wen_0_reg = 0;
		end
	end
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_44_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_52_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_7.bb_1_active_in_state_7_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_7_in_data = eq_51_out;
		end else begin
			bb_1_active_in_state_7_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_7.bb_1_predecessor_in_state_7_in_data
	always @(*) begin
		if (eq_59_out) begin 
			bb_1_predecessor_in_state_7_in_data = state_7_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_7_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_1.bb_2_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_1_in_data = eq_45_out;
		end else begin
			bb_2_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_2.bb_2_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_2_in_data = eq_46_out;
		end else begin
			bb_2_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_3.bb_2_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_3_in_data = eq_47_out;
		end else begin
			bb_2_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_4.bb_2_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_4_in_data = eq_48_out;
		end else begin
			bb_2_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_5.bb_2_active_in_state_5_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_5_in_data = eq_49_out;
		end else begin
			bb_2_active_in_state_5_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_6.bb_2_active_in_state_6_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_6_in_data = eq_50_out;
		end else begin
			bb_2_active_in_state_6_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_1.bb_2_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_53_out) begin 
			bb_2_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_2.bb_2_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_54_out) begin 
			bb_2_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_3.bb_2_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_55_out) begin 
			bb_2_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_4.bb_2_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_56_out) begin 
			bb_2_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_5.bb_2_predecessor_in_state_5_in_data
	always @(*) begin
		if (eq_57_out) begin 
			bb_2_predecessor_in_state_5_in_data = state_5_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_5_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_6.bb_2_predecessor_in_state_6_in_data
	always @(*) begin
		if (eq_58_out) begin 
			bb_2_predecessor_in_state_6_in_data = state_6_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_6_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_12_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_13_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_2_happened_in_state_1.br_2_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_14_out) begin 
			br_2_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_15_out) begin 
			br_2_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_2_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_2_happened_in_state_2.br_2_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_19_out) begin 
			br_2_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_20_out) begin 
			br_2_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_2_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_2_happened_in_state_3.br_2_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_24_out) begin 
			br_2_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_25_out) begin 
			br_2_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_2_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_2_happened_in_state_4.br_2_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_29_out) begin 
			br_2_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_30_out) begin 
			br_2_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_2_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_2_happened_in_state_5.br_2_happened_in_state_5_in_data
	always @(*) begin
		if (andOp_34_out) begin 
			br_2_happened_in_state_5_in_data = 1'd1;
		end else if (notOp_35_out) begin 
			br_2_happened_in_state_5_in_data = 1'd0;
		end else begin
			br_2_happened_in_state_5_in_data = 0;
		end
	end
	// controller for br_2_happened_in_state_6.br_2_happened_in_state_6_in_data
	always @(*) begin
		if (andOp_39_out) begin 
			br_2_happened_in_state_6_in_data = 1'd1;
		end else if (notOp_40_out) begin 
			br_2_happened_in_state_6_in_data = 1'd0;
		end else begin
			br_2_happened_in_state_6_in_data = 0;
		end
	end
	// controller for concat_61.concat_61_in0
	// controller for concat_61.concat_61_in1
	// Insensitive connections
	assign concat_61_in0 = data_in_1_4_out_data;
	assign concat_61_in1 = 32'd0;
	// controller for concat_62.concat_62_in0
	// controller for concat_62.concat_62_in1
	// Insensitive connections
	assign concat_62_in0 = 32'd2;
	assign concat_62_in1 = 32'd0;
	// controller for data_in_0_1.data_in_0_1_in_data
	always @(*) begin
		if (eq_136_out) begin 
			data_in_0_1_in_data = data_store_0_0;
		end else begin
			data_in_0_1_in_data = 0;
		end
	end
	// controller for data_in_1_4.data_in_1_4_in_data
	always @(*) begin
		if (eq_137_out) begin 
			data_in_1_4_in_data = data_store_0_0;
		end else if (eq_138_out) begin 
			data_in_1_4_in_data = data_store_1_3;
		end else begin
			data_in_1_4_in_data = 0;
		end
	end
	// controller for data_in_2_6.data_in_2_6_in_data
	always @(*) begin
		if (eq_141_out) begin 
			data_in_2_6_in_data = data_store_1_2;
		end else if (eq_142_out) begin 
			data_in_2_6_in_data = data_store_2_5;
		end else begin
			data_in_2_6_in_data = 0;
		end
	end
	// controller for data_in_3_10.data_in_3_10_in_data
	always @(*) begin
		if (eq_145_out) begin 
			data_in_3_10_in_data = data_store_2_7;
		end else if (eq_146_out) begin 
			data_in_3_10_in_data = 32'd0;
		end else begin
			data_in_3_10_in_data = 0;
		end
	end
	// controller for data_in_3_11.data_in_3_11_in_data
	always @(*) begin
		if (eq_145_out) begin 
			data_in_3_11_in_data = data_store_2_8;
		end else if (eq_146_out) begin 
			data_in_3_11_in_data = 32'd0;
		end else begin
			data_in_3_11_in_data = 0;
		end
	end
	// controller for data_in_3_9.data_in_3_9_in_data
	always @(*) begin
		if (eq_145_out) begin 
			data_in_3_9_in_data = data_store_2_5;
		end else if (eq_146_out) begin 
			data_in_3_9_in_data = 32'd0;
		end else begin
			data_in_3_9_in_data = 0;
		end
	end
	// controller for eq_103.eq_103_in0
	// controller for eq_103.eq_103_in1
	// Insensitive connections
	assign eq_103_in0 = counter__99;
	assign eq_103_in1 = 32'd1;
	// controller for eq_136.eq_136_in0
	// controller for eq_136.eq_136_in1
	// Insensitive connections
	assign eq_136_in0 = 32'd0;
	assign eq_136_in1 = state_0_last_state;
	// controller for eq_137.eq_137_in0
	// controller for eq_137.eq_137_in1
	// Insensitive connections
	assign eq_137_in0 = 32'd0;
	assign eq_137_in1 = state_1_last_state;
	// controller for eq_138.eq_138_in0
	// controller for eq_138.eq_138_in1
	// Insensitive connections
	assign eq_138_in0 = 32'd1;
	assign eq_138_in1 = state_1_last_state;
	// controller for eq_141.eq_141_in0
	// controller for eq_141.eq_141_in1
	// Insensitive connections
	assign eq_141_in0 = 32'd1;
	assign eq_141_in1 = state_2_last_state;
	// controller for eq_142.eq_142_in0
	// controller for eq_142.eq_142_in1
	// Insensitive connections
	assign eq_142_in0 = 32'd2;
	assign eq_142_in1 = state_2_last_state;
	// controller for eq_145.eq_145_in0
	// controller for eq_145.eq_145_in1
	// Insensitive connections
	assign eq_145_in0 = 32'd2;
	assign eq_145_in1 = state_3_last_state;
	// controller for eq_146.eq_146_in0
	// controller for eq_146.eq_146_in1
	// Insensitive connections
	assign eq_146_in0 = 32'd3;
	assign eq_146_in1 = state_3_last_state;
	// controller for eq_147.eq_147_in0
	// controller for eq_147.eq_147_in1
	// Insensitive connections
	assign eq_147_in0 = 32'd3;
	assign eq_147_in1 = state_4_last_state;
	// controller for eq_148.eq_148_in0
	// controller for eq_148.eq_148_in1
	// Insensitive connections
	assign eq_148_in0 = 32'd4;
	assign eq_148_in1 = state_4_last_state;
	// controller for eq_149.eq_149_in0
	// controller for eq_149.eq_149_in1
	// Insensitive connections
	assign eq_149_in0 = 32'd4;
	assign eq_149_in1 = state_5_last_state;
	// controller for eq_150.eq_150_in0
	// controller for eq_150.eq_150_in1
	// Insensitive connections
	assign eq_150_in0 = 32'd5;
	assign eq_150_in1 = state_5_last_state;
	// controller for eq_151.eq_151_in0
	// controller for eq_151.eq_151_in1
	// Insensitive connections
	assign eq_151_in0 = 32'd5;
	assign eq_151_in1 = state_6_last_state;
	// controller for eq_152.eq_152_in0
	// controller for eq_152.eq_152_in1
	// Insensitive connections
	assign eq_152_in0 = 32'd6;
	assign eq_152_in1 = state_6_last_state;
	// controller for eq_153.eq_153_in0
	// controller for eq_153.eq_153_in1
	// Insensitive connections
	assign eq_153_in0 = 32'd1;
	assign eq_153_in1 = state_7_last_state;
	// controller for eq_154.eq_154_in0
	// controller for eq_154.eq_154_in1
	// Insensitive connections
	assign eq_154_in0 = 32'd6;
	assign eq_154_in1 = state_7_last_state;
	// controller for eq_155.eq_155_in0
	// controller for eq_155.eq_155_in1
	// Insensitive connections
	assign eq_155_in0 = 32'd7;
	assign eq_155_in1 = state_7_last_state;
	// controller for eq_44.eq_44_in0
	// controller for eq_44.eq_44_in1
	// Insensitive connections
	assign eq_44_in0 = 32'd0;
	assign eq_44_in1 = state_0_entry_BB_reg;
	// controller for eq_45.eq_45_in0
	// controller for eq_45.eq_45_in1
	// Insensitive connections
	assign eq_45_in0 = 32'd2;
	assign eq_45_in1 = state_1_entry_BB_reg;
	// controller for eq_46.eq_46_in0
	// controller for eq_46.eq_46_in1
	// Insensitive connections
	assign eq_46_in0 = 32'd2;
	assign eq_46_in1 = state_2_entry_BB_reg;
	// controller for eq_47.eq_47_in0
	// controller for eq_47.eq_47_in1
	// Insensitive connections
	assign eq_47_in0 = 32'd2;
	assign eq_47_in1 = state_3_entry_BB_reg;
	// controller for eq_48.eq_48_in0
	// controller for eq_48.eq_48_in1
	// Insensitive connections
	assign eq_48_in0 = 32'd2;
	assign eq_48_in1 = state_4_entry_BB_reg;
	// controller for eq_49.eq_49_in0
	// controller for eq_49.eq_49_in1
	// Insensitive connections
	assign eq_49_in0 = 32'd2;
	assign eq_49_in1 = state_5_entry_BB_reg;
	// controller for eq_50.eq_50_in0
	// controller for eq_50.eq_50_in1
	// Insensitive connections
	assign eq_50_in0 = 32'd2;
	assign eq_50_in1 = state_6_entry_BB_reg;
	// controller for eq_51.eq_51_in0
	// controller for eq_51.eq_51_in1
	// Insensitive connections
	assign eq_51_in0 = 32'd1;
	assign eq_51_in1 = state_7_entry_BB_reg;
	// controller for eq_52.eq_52_in0
	// controller for eq_52.eq_52_in1
	// Insensitive connections
	assign eq_52_in0 = 32'd0;
	assign eq_52_in1 = state_0_entry_BB_reg;
	// controller for eq_53.eq_53_in0
	// controller for eq_53.eq_53_in1
	// Insensitive connections
	assign eq_53_in0 = 32'd2;
	assign eq_53_in1 = state_1_entry_BB_reg;
	// controller for eq_54.eq_54_in0
	// controller for eq_54.eq_54_in1
	// Insensitive connections
	assign eq_54_in0 = 32'd2;
	assign eq_54_in1 = state_2_entry_BB_reg;
	// controller for eq_55.eq_55_in0
	// controller for eq_55.eq_55_in1
	// Insensitive connections
	assign eq_55_in0 = 32'd2;
	assign eq_55_in1 = state_3_entry_BB_reg;
	// controller for eq_56.eq_56_in0
	// controller for eq_56.eq_56_in1
	// Insensitive connections
	assign eq_56_in0 = 32'd2;
	assign eq_56_in1 = state_4_entry_BB_reg;
	// controller for eq_57.eq_57_in0
	// controller for eq_57.eq_57_in1
	// Insensitive connections
	assign eq_57_in0 = 32'd2;
	assign eq_57_in1 = state_5_entry_BB_reg;
	// controller for eq_58.eq_58_in0
	// controller for eq_58.eq_58_in1
	// Insensitive connections
	assign eq_58_in0 = 32'd2;
	assign eq_58_in1 = state_6_entry_BB_reg;
	// controller for eq_59.eq_59_in0
	// controller for eq_59.eq_59_in1
	// Insensitive connections
	assign eq_59_in0 = 32'd1;
	assign eq_59_in1 = state_7_entry_BB_reg;
	// controller for icmp_icmp3.icmp_icmp3_in0
	// controller for icmp_icmp3.icmp_icmp3_in1
	// Insensitive connections
	assign icmp_icmp3_in0 = add_add2_out;
	assign icmp_icmp3_in1 = 32'd5;
	// controller for in_pipeline_0.in_pipeline_0_in_data
	always @(*) begin
		if (1'd1) begin 
			in_pipeline_0_in_data = orOp_135_out;
		end else begin
			in_pipeline_0_in_data = 0;
		end
	end
	// controller for mul_mul6.mul_mul6_in0
	// controller for mul_mul6.mul_mul6_in1
	// Insensitive connections
	assign mul_mul6_in0 = arg_0_rdata_0;
	assign mul_mul6_in1 = 32'd3;
	// controller for mul_mul9.mul_mul9_in0
	// controller for mul_mul9.mul_mul9_in1
	// Insensitive connections
	assign mul_mul9_in0 = data_in_3_11_out_data;
	assign mul_mul9_in1 = 32'd7;
	// controller for notOp_101.notOp_101_in0
	// Insensitive connections
	assign notOp_101_in0 = state_1_is_active;
	// controller for notOp_112.notOp_112_in0
	// Insensitive connections
	assign notOp_112_in0 = andOp_105_out;
	// controller for notOp_114.notOp_114_in0
	// Insensitive connections
	assign notOp_114_in0 = andOp_12_out;
	// controller for notOp_116.notOp_116_in0
	// Insensitive connections
	assign notOp_116_in0 = andOp_106_out;
	// controller for notOp_118.notOp_118_in0
	// Insensitive connections
	assign notOp_118_in0 = andOp_107_out;
	// controller for notOp_120.notOp_120_in0
	// Insensitive connections
	assign notOp_120_in0 = andOp_108_out;
	// controller for notOp_122.notOp_122_in0
	// Insensitive connections
	assign notOp_122_in0 = andOp_109_out;
	// controller for notOp_124.notOp_124_in0
	// Insensitive connections
	assign notOp_124_in0 = andOp_110_out;
	// controller for notOp_126.notOp_126_in0
	// Insensitive connections
	assign notOp_126_in0 = andOp_111_out;
	// controller for notOp_128.notOp_128_in0
	// Insensitive connections
	assign notOp_128_in0 = andOp_86_out;
	// controller for notOp_13.notOp_13_in0
	// Insensitive connections
	assign notOp_13_in0 = andOp_12_out;
	// controller for notOp_15.notOp_15_in0
	// Insensitive connections
	assign notOp_15_in0 = andOp_14_out;
	// controller for notOp_156.notOp_156_in0
	// Insensitive connections
	assign notOp_156_in0 = state_1_is_active;
	// controller for notOp_157.notOp_157_in0
	// Insensitive connections
	assign notOp_157_in0 = state_1_is_active;
	// controller for notOp_17.notOp_17_in0
	// Insensitive connections
	assign notOp_17_in0 = icmp_icmp3_out;
	// controller for notOp_20.notOp_20_in0
	// Insensitive connections
	assign notOp_20_in0 = andOp_19_out;
	// controller for notOp_22.notOp_22_in0
	// Insensitive connections
	assign notOp_22_in0 = icmp_icmp3_out;
	// controller for notOp_25.notOp_25_in0
	// Insensitive connections
	assign notOp_25_in0 = andOp_24_out;
	// controller for notOp_27.notOp_27_in0
	// Insensitive connections
	assign notOp_27_in0 = icmp_icmp3_out;
	// controller for notOp_30.notOp_30_in0
	// Insensitive connections
	assign notOp_30_in0 = andOp_29_out;
	// controller for notOp_32.notOp_32_in0
	// Insensitive connections
	assign notOp_32_in0 = icmp_icmp3_out;
	// controller for notOp_35.notOp_35_in0
	// Insensitive connections
	assign notOp_35_in0 = andOp_34_out;
	// controller for notOp_37.notOp_37_in0
	// Insensitive connections
	assign notOp_37_in0 = icmp_icmp3_out;
	// controller for notOp_40.notOp_40_in0
	// Insensitive connections
	assign notOp_40_in0 = andOp_39_out;
	// controller for notOp_42.notOp_42_in0
	// Insensitive connections
	assign notOp_42_in0 = icmp_icmp3_out;
	// controller for notOp_74.notOp_74_in0
	// Insensitive connections
	assign notOp_74_in0 = state_1_is_active;
	// controller for notOp_76.notOp_76_in0
	// Insensitive connections
	assign notOp_76_in0 = state_2_is_active;
	// controller for notOp_78.notOp_78_in0
	// Insensitive connections
	assign notOp_78_in0 = state_3_is_active;
	// controller for notOp_80.notOp_80_in0
	// Insensitive connections
	assign notOp_80_in0 = state_4_is_active;
	// controller for notOp_82.notOp_82_in0
	// Insensitive connections
	assign notOp_82_in0 = state_5_is_active;
	// controller for notOp_87.notOp_87_in0
	// Insensitive connections
	assign notOp_87_in0 = state_1_is_active;
	// controller for notOp_89.notOp_89_in0
	// Insensitive connections
	assign notOp_89_in0 = state_2_is_active;
	// controller for notOp_91.notOp_91_in0
	// Insensitive connections
	assign notOp_91_in0 = state_3_is_active;
	// controller for notOp_93.notOp_93_in0
	// Insensitive connections
	assign notOp_93_in0 = state_4_is_active;
	// controller for notOp_95.notOp_95_in0
	// Insensitive connections
	assign notOp_95_in0 = state_5_is_active;
	// controller for orOp_130.orOp_130_in0
	// controller for orOp_130.orOp_130_in1
	// Insensitive connections
	assign orOp_130_in0 = state_1_is_active;
	assign orOp_130_in1 = 1'd0;
	// controller for orOp_131.orOp_131_in0
	// controller for orOp_131.orOp_131_in1
	// Insensitive connections
	assign orOp_131_in0 = state_2_is_active;
	assign orOp_131_in1 = orOp_130_out;
	// controller for orOp_132.orOp_132_in0
	// controller for orOp_132.orOp_132_in1
	// Insensitive connections
	assign orOp_132_in0 = state_3_is_active;
	assign orOp_132_in1 = orOp_131_out;
	// controller for orOp_133.orOp_133_in0
	// controller for orOp_133.orOp_133_in1
	// Insensitive connections
	assign orOp_133_in0 = state_4_is_active;
	assign orOp_133_in1 = orOp_132_out;
	// controller for orOp_134.orOp_134_in0
	// controller for orOp_134.orOp_134_in1
	// Insensitive connections
	assign orOp_134_in0 = state_5_is_active;
	assign orOp_134_in1 = orOp_133_out;
	// controller for orOp_135.orOp_135_in0
	// controller for orOp_135.orOp_135_in1
	// Insensitive connections
	assign orOp_135_in0 = state_6_is_active;
	assign orOp_135_in1 = orOp_134_out;
	// controller for phi_phi1.phi_phi1_in
	// controller for phi_phi1.phi_phi1_last_block
	// controller for phi_phi1.phi_phi1_s
	// Insensitive connections
	assign phi_phi1_in = concat_61_out;
	assign phi_phi1_last_block = bb_2_predecessor_in_state_1_out_data;
	assign phi_phi1_s = concat_62_out;
	// controller for ret13.valid_reg
	always @(*) begin
		if (andOp_73_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			counter__99 <= 0;
		end else begin
			if (andOp_102_out) begin
				counter__99 <= add_100_out;
			end
			if (state_1_is_active) begin
				counter__99 <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_0 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_0 <= data_in_0_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_2 <= 0;
		end else begin
			if (andOp_139_out) begin
				data_store_1_2 <= phi_phi1_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_3 <= 0;
		end else begin
			if (andOp_140_out) begin
				data_store_1_3 <= add_add2_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_5 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_5 <= data_in_2_6_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_7 <= 0;
		end else begin
			if (andOp_143_out) begin
				data_store_2_7 <= mul_mul6_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_8 <= 0;
		end else begin
			if (andOp_144_out) begin
				data_store_2_8 <= arg_0_rdata_0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			delayed_signal__104 <= 0;
		end else begin
			if (state_1_is_active) begin
				delayed_signal__104 <= andOp_16_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_111_out) begin
				global_state <= 32'd7;
			end
			if (andOp_12_out) begin
				global_state <= 32'd200000;
			end
			if (andOp_85_out) begin
				global_state <= 32'd7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			out_of_pipe_1_7 <= 0;
		end else begin
			if (andOp_18_out) begin
				out_of_pipe_1_7 <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			out_of_pipe_bb_1_7 <= 0;
		end else begin
			if (andOp_18_out) begin
				out_of_pipe_bb_1_7 <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (1'd1) begin
				state_0_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_12_out) begin
				state_1_entry_BB_reg <= 32'd2;
			end
			if (andOp_16_out) begin
				state_1_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_105_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_115_out) begin
				state_1_is_active <= 1'd0;
			end
			if (andOp_12_out) begin
				state_1_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_12_out) begin
				state_1_last_BB_reg <= 32'd0;
			end
			if (andOp_16_out) begin
				state_1_last_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_12_out) begin
				state_1_last_state <= 32'd0;
			end
			if (andOp_16_out) begin
				state_1_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_106_out) begin
				state_2_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_106_out) begin
				state_2_is_active <= 1'd1;
			end
			if (andOp_117_out) begin
				state_2_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_106_out) begin
				state_2_last_BB_reg <= bb_2_predecessor_in_state_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_106_out) begin
				state_2_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_107_out) begin
				state_3_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_107_out) begin
				state_3_is_active <= 1'd1;
			end
			if (andOp_119_out) begin
				state_3_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_107_out) begin
				state_3_last_BB_reg <= bb_2_predecessor_in_state_2_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_state <= 0;
		end else begin
			if (andOp_107_out) begin
				state_3_last_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_108_out) begin
				state_4_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_108_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_121_out) begin
				state_4_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_108_out) begin
				state_4_last_BB_reg <= bb_2_predecessor_in_state_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_state <= 0;
		end else begin
			if (andOp_108_out) begin
				state_4_last_state <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_entry_BB_reg <= 0;
		end else begin
			if (andOp_109_out) begin
				state_5_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_is_active <= 0;
		end else begin
			if (andOp_109_out) begin
				state_5_is_active <= 1'd1;
			end
			if (andOp_123_out) begin
				state_5_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_last_BB_reg <= 0;
		end else begin
			if (andOp_109_out) begin
				state_5_last_BB_reg <= bb_2_predecessor_in_state_4_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_last_state <= 0;
		end else begin
			if (andOp_109_out) begin
				state_5_last_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_entry_BB_reg <= 0;
		end else begin
			if (andOp_110_out) begin
				state_6_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_is_active <= 0;
		end else begin
			if (andOp_110_out) begin
				state_6_is_active <= 1'd1;
			end
			if (andOp_125_out) begin
				state_6_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_last_BB_reg <= 0;
		end else begin
			if (andOp_110_out) begin
				state_6_last_BB_reg <= bb_2_predecessor_in_state_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_last_state <= 0;
		end else begin
			if (andOp_110_out) begin
				state_6_last_state <= 32'd5;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_entry_BB_reg <= 0;
		end else begin
			if (andOp_111_out) begin
				state_7_entry_BB_reg <= 32'd1;
			end
			if (andOp_98_out) begin
				state_7_entry_BB_reg <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_is_active <= 0;
		end else begin
			if (andOp_111_out) begin
				state_7_is_active <= 1'd1;
			end
			if (andOp_129_out) begin
				state_7_is_active <= 1'd0;
			end
			if (andOp_86_out) begin
				state_7_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_last_BB_reg <= 0;
		end else begin
			if (andOp_111_out) begin
				state_7_last_BB_reg <= bb_1_predecessor_in_state_7_out_data;
			end
			if (andOp_18_out) begin
				state_7_last_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_last_state <= 0;
		end else begin
			if (andOp_111_out) begin
				state_7_last_state <= 32'd7;
			end
			if (andOp_18_out) begin
				state_7_last_state <= 32'd1;
			end
		end
	end

endmodule

