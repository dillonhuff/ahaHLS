module channel_reduce_4(input [0:0] clk, input [0:0] rst, output [31:0] in_in_data, output [0:0] in_read_valid, output [0:0] in_rst, output [0:0] in_write_valid, input [31:0] in_out_data, input [0:0] in_read_ready, input [0:0] in_write_ready, output [0:0] valid, output [31:0] out_in_data, output [0:0] out_read_valid, output [0:0] out_rst, output [0:0] out_write_valid, input [31:0] out_out_data, input [0:0] out_read_ready, input [0:0] out_write_ready);

	reg [31:0] in_in_data_reg;
	reg [0:0] in_read_valid_reg;
	reg [0:0] in_rst_reg;
	reg [0:0] in_write_valid_reg;
	reg [0:0] valid_reg;
	reg [31:0] out_in_data_reg;
	reg [0:0] out_read_valid_reg;
	reg [0:0] out_rst_reg;
	reg [0:0] out_write_valid_reg;

	assign in_in_data = in_in_data_reg;
	assign in_read_valid = in_read_valid_reg;
	assign in_rst = in_rst_reg;
	assign in_write_valid = in_write_valid_reg;
	assign valid = valid_reg;
	assign out_in_data = out_in_data_reg;
	assign out_read_valid = out_read_valid_reg;
	assign out_rst = out_rst_reg;
	assign out_write_valid = out_write_valid_reg;

	// Start debug wires and ports

	initial begin
	end





	// End debug wires and ports

	// Start Functional Units
	br_dummy br_unit();

	add alloca_0();

	add bitcast_1();

	add call_2();

	reg [31:0] raddr_ram_0_reg;
	reg [31:0] waddr_ram_0_reg;
	reg [31:0] wdata_ram_0_reg;
	reg [0:0] wen_ram_0_reg;
	wire [31:0] rdata_ram_0;
	register #(.WIDTH(32)) ram_0(.clk(clk), .raddr(raddr_ram_0_reg), .rdata(rdata_ram_0), .rst(rst), .waddr(waddr_ram_0_reg), .wdata(wdata_ram_0_reg), .wen(wen_ram_0_reg));

	add call_21();

	reg [63:0] phi_in_phi_7;
	reg [31:0] phi_last_block_phi_7;
	reg [63:0] phi_s_phi_7;
	wire [31:0] phi_out_phi_7;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_7(.in(phi_in_phi_7), .last_block(phi_last_block_phi_7), .out(phi_out_phi_7), .s(phi_s_phi_7));

	reg [31:0] add_in0_add_14;
	reg [31:0] add_in1_add_14;
	wire [31:0] add_out_add_14;
	add #(.WIDTH(32)) add_add_14(.in0(add_in0_add_14), .in1(add_in1_add_14), .out(add_out_add_14));

	reg [31:0] add_in0_add_16;
	reg [31:0] add_in1_add_16;
	wire [31:0] add_out_add_16;
	add #(.WIDTH(32)) add_add_16(.in0(add_in0_add_16), .in1(add_in1_add_16), .out(add_out_add_16));

	reg [31:0] cmp_in0_icmp_17;
	reg [31:0] cmp_in1_icmp_17;
	wire [0:0] cmp_out_icmp_17;
	eq #(.WIDTH(32)) icmp_17(.in0(cmp_in0_icmp_17), .in1(cmp_in1_icmp_17), .out(cmp_out_icmp_17));

	reg [31:0] data_in_1_1_in_data;
	wire [31:0] data_in_1_1_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_1(.in_data(data_in_1_1_in_data), .out_data(data_in_1_1_out_data));

	reg [31:0] data_in_1_3_in_data;
	wire [31:0] data_in_1_3_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_3(.in_data(data_in_1_3_in_data), .out_data(data_in_1_3_out_data));

	reg [31:0] data_in_1_5_in_data;
	wire [31:0] data_in_1_5_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_5(.in_data(data_in_1_5_in_data), .out_data(data_in_1_5_out_data));

	reg [0:0] data_in_1_7_in_data;
	wire [0:0] data_in_1_7_out_data;
	hls_wire #(.WIDTH(1)) data_in_1_7(.in_data(data_in_1_7_in_data), .out_data(data_in_1_7_out_data));

	reg [31:0] data_in_2_9_in_data;
	wire [31:0] data_in_2_9_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_9(.in_data(data_in_2_9_in_data), .out_data(data_in_2_9_out_data));

	reg [31:0] data_in_2_11_in_data;
	wire [31:0] data_in_2_11_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_11(.in_data(data_in_2_11_in_data), .out_data(data_in_2_11_out_data));

	reg [31:0] data_in_2_13_in_data;
	wire [31:0] data_in_2_13_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_13(.in_data(data_in_2_13_in_data), .out_data(data_in_2_13_out_data));

	reg [0:0] data_in_2_15_in_data;
	wire [0:0] data_in_2_15_out_data;
	hls_wire #(.WIDTH(1)) data_in_2_15(.in_data(data_in_2_15_in_data), .out_data(data_in_2_15_out_data));

	reg [31:0] data_in_3_17_in_data;
	wire [31:0] data_in_3_17_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_17(.in_data(data_in_3_17_in_data), .out_data(data_in_3_17_out_data));

	reg [31:0] data_in_3_19_in_data;
	wire [31:0] data_in_3_19_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_19(.in_data(data_in_3_19_in_data), .out_data(data_in_3_19_out_data));

	reg [31:0] data_in_3_21_in_data;
	wire [31:0] data_in_3_21_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_21(.in_data(data_in_3_21_in_data), .out_data(data_in_3_21_out_data));

	reg [0:0] data_in_3_23_in_data;
	wire [0:0] data_in_3_23_out_data;
	hls_wire #(.WIDTH(1)) data_in_3_23(.in_data(data_in_3_23_in_data), .out_data(data_in_3_23_out_data));

	reg [31:0] data_in_4_25_in_data;
	wire [31:0] data_in_4_25_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_25(.in_data(data_in_4_25_in_data), .out_data(data_in_4_25_out_data));

	reg [31:0] data_in_4_27_in_data;
	wire [31:0] data_in_4_27_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_27(.in_data(data_in_4_27_in_data), .out_data(data_in_4_27_out_data));

	reg [31:0] data_in_4_29_in_data;
	wire [31:0] data_in_4_29_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_29(.in_data(data_in_4_29_in_data), .out_data(data_in_4_29_out_data));

	reg [0:0] data_in_4_31_in_data;
	wire [0:0] data_in_4_31_out_data;
	hls_wire #(.WIDTH(1)) data_in_4_31(.in_data(data_in_4_31_in_data), .out_data(data_in_4_31_out_data));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] bb_0_active_in_state_1_in_data;
	wire [0:0] bb_0_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_1(.in_data(bb_0_active_in_state_1_in_data), .out_data(bb_0_active_in_state_1_out_data));

	reg [31:0] bb_0_predecessor_in_state_1_in_data;
	wire [31:0] bb_0_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_1(.in_data(bb_0_predecessor_in_state_1_in_data), .out_data(bb_0_predecessor_in_state_1_out_data));

	reg [0:0] bb_3_active_in_state_1_in_data;
	wire [0:0] bb_3_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_1(.in_data(bb_3_active_in_state_1_in_data), .out_data(bb_3_active_in_state_1_out_data));

	reg [31:0] bb_3_predecessor_in_state_1_in_data;
	wire [31:0] bb_3_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_1(.in_data(bb_3_predecessor_in_state_1_in_data), .out_data(bb_3_predecessor_in_state_1_out_data));

	reg [0:0] bb_8_active_in_state_1_in_data;
	wire [0:0] bb_8_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active_in_state_1(.in_data(bb_8_active_in_state_1_in_data), .out_data(bb_8_active_in_state_1_out_data));

	reg [31:0] bb_8_predecessor_in_state_1_in_data;
	wire [31:0] bb_8_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor_in_state_1(.in_data(bb_8_predecessor_in_state_1_in_data), .out_data(bb_8_predecessor_in_state_1_out_data));

	reg [0:0] bb_9_active_in_state_1_in_data;
	wire [0:0] bb_9_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_9_active_in_state_1(.in_data(bb_9_active_in_state_1_in_data), .out_data(bb_9_active_in_state_1_out_data));

	reg [31:0] bb_9_predecessor_in_state_1_in_data;
	wire [31:0] bb_9_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_9_predecessor_in_state_1(.in_data(bb_9_predecessor_in_state_1_in_data), .out_data(bb_9_predecessor_in_state_1_out_data));

	reg [0:0] bb_10_active_in_state_2_in_data;
	wire [0:0] bb_10_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_2(.in_data(bb_10_active_in_state_2_in_data), .out_data(bb_10_active_in_state_2_out_data));

	reg [31:0] bb_10_predecessor_in_state_2_in_data;
	wire [31:0] bb_10_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_2(.in_data(bb_10_predecessor_in_state_2_in_data), .out_data(bb_10_predecessor_in_state_2_out_data));

	reg [0:0] bb_4_active_in_state_3_in_data;
	wire [0:0] bb_4_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_3(.in_data(bb_4_active_in_state_3_in_data), .out_data(bb_4_active_in_state_3_out_data));

	reg [31:0] bb_4_predecessor_in_state_3_in_data;
	wire [31:0] bb_4_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_3(.in_data(bb_4_predecessor_in_state_3_in_data), .out_data(bb_4_predecessor_in_state_3_out_data));

	reg [0:0] bb_10_active_in_state_3_in_data;
	wire [0:0] bb_10_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_3(.in_data(bb_10_active_in_state_3_in_data), .out_data(bb_10_active_in_state_3_out_data));

	reg [31:0] bb_10_predecessor_in_state_3_in_data;
	wire [31:0] bb_10_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_3(.in_data(bb_10_predecessor_in_state_3_in_data), .out_data(bb_10_predecessor_in_state_3_out_data));

	reg [0:0] bb_7_active_in_state_4_in_data;
	wire [0:0] bb_7_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_7_active_in_state_4(.in_data(bb_7_active_in_state_4_in_data), .out_data(bb_7_active_in_state_4_out_data));

	reg [31:0] bb_7_predecessor_in_state_4_in_data;
	wire [31:0] bb_7_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_7_predecessor_in_state_4(.in_data(bb_7_predecessor_in_state_4_in_data), .out_data(bb_7_predecessor_in_state_4_out_data));

	reg [0:0] bb_6_active_in_state_4_in_data;
	wire [0:0] bb_6_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_6_active_in_state_4(.in_data(bb_6_active_in_state_4_in_data), .out_data(bb_6_active_in_state_4_out_data));

	reg [31:0] bb_6_predecessor_in_state_4_in_data;
	wire [31:0] bb_6_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_6_predecessor_in_state_4(.in_data(bb_6_predecessor_in_state_4_in_data), .out_data(bb_6_predecessor_in_state_4_out_data));

	reg [0:0] bb_5_active_in_state_4_in_data;
	wire [0:0] bb_5_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_5_active_in_state_4(.in_data(bb_5_active_in_state_4_in_data), .out_data(bb_5_active_in_state_4_out_data));

	reg [31:0] bb_5_predecessor_in_state_4_in_data;
	wire [31:0] bb_5_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_5_predecessor_in_state_4(.in_data(bb_5_predecessor_in_state_4_in_data), .out_data(bb_5_predecessor_in_state_4_out_data));

	reg [0:0] bb_4_active_in_state_4_in_data;
	wire [0:0] bb_4_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_4(.in_data(bb_4_active_in_state_4_in_data), .out_data(bb_4_active_in_state_4_out_data));

	reg [31:0] bb_4_predecessor_in_state_4_in_data;
	wire [31:0] bb_4_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_4(.in_data(bb_4_predecessor_in_state_4_in_data), .out_data(bb_4_predecessor_in_state_4_out_data));

	reg [0:0] bb_2_active_in_state_4_in_data;
	wire [0:0] bb_2_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_4(.in_data(bb_2_active_in_state_4_in_data), .out_data(bb_2_active_in_state_4_out_data));

	reg [31:0] bb_2_predecessor_in_state_4_in_data;
	wire [31:0] bb_2_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_4(.in_data(bb_2_predecessor_in_state_4_in_data), .out_data(bb_2_predecessor_in_state_4_out_data));

	reg [0:0] bb_1_active_in_state_4_in_data;
	wire [0:0] bb_1_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_4(.in_data(bb_1_active_in_state_4_in_data), .out_data(bb_1_active_in_state_4_out_data));

	reg [31:0] bb_1_predecessor_in_state_4_in_data;
	wire [31:0] bb_1_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_4(.in_data(bb_1_predecessor_in_state_4_in_data), .out_data(bb_1_predecessor_in_state_4_out_data));

	reg [0:0] andOp_32_in0;
	reg [0:0] andOp_32_in1;
	wire [0:0] andOp_32_out;
	andOp #(.WIDTH(1)) andOp_32(.in0(andOp_32_in0), .in1(andOp_32_in1), .out(andOp_32_out));

	reg [0:0] andOp_33_in0;
	reg [0:0] andOp_33_in1;
	wire [0:0] andOp_33_out;
	andOp #(.WIDTH(1)) andOp_33(.in0(andOp_33_in0), .in1(andOp_33_in1), .out(andOp_33_out));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] notOp_34_in0;
	wire [0:0] notOp_34_out;
	notOp #(.WIDTH(1)) notOp_34(.in(notOp_34_in0), .out(notOp_34_out));

	reg [0:0] andOp_35_in0;
	reg [0:0] andOp_35_in1;
	wire [0:0] andOp_35_out;
	andOp #(.WIDTH(1)) andOp_35(.in0(andOp_35_in0), .in1(andOp_35_in1), .out(andOp_35_out));

	reg [0:0] andOp_36_in0;
	reg [0:0] andOp_36_in1;
	wire [0:0] andOp_36_out;
	andOp #(.WIDTH(1)) andOp_36(.in0(andOp_36_in0), .in1(andOp_36_in1), .out(andOp_36_out));

	reg [0:0] br_0_happened_in_state_1_in_data;
	wire [0:0] br_0_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_1(.in_data(br_0_happened_in_state_1_in_data), .out_data(br_0_happened_in_state_1_out_data));

	reg [0:0] notOp_37_in0;
	wire [0:0] notOp_37_out;
	notOp #(.WIDTH(1)) notOp_37(.in(notOp_37_in0), .out(notOp_37_out));

	reg [0:0] andOp_38_in0;
	reg [0:0] andOp_38_in1;
	wire [0:0] andOp_38_out;
	andOp #(.WIDTH(1)) andOp_38(.in0(andOp_38_in0), .in1(andOp_38_in1), .out(andOp_38_out));

	reg [0:0] andOp_39_in0;
	reg [0:0] andOp_39_in1;
	wire [0:0] andOp_39_out;
	andOp #(.WIDTH(1)) andOp_39(.in0(andOp_39_in0), .in1(andOp_39_in1), .out(andOp_39_out));

	reg [0:0] br_3_happened_in_state_1_in_data;
	wire [0:0] br_3_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_1(.in_data(br_3_happened_in_state_1_in_data), .out_data(br_3_happened_in_state_1_out_data));

	reg [0:0] notOp_40_in0;
	wire [0:0] notOp_40_out;
	notOp #(.WIDTH(1)) notOp_40(.in(notOp_40_in0), .out(notOp_40_out));

	reg [0:0] andOp_41_in0;
	reg [0:0] andOp_41_in1;
	wire [0:0] andOp_41_out;
	andOp #(.WIDTH(1)) andOp_41(.in0(andOp_41_in0), .in1(andOp_41_in1), .out(andOp_41_out));

	reg [0:0] andOp_42_in0;
	reg [0:0] andOp_42_in1;
	wire [0:0] andOp_42_out;
	andOp #(.WIDTH(1)) andOp_42(.in0(andOp_42_in0), .in1(andOp_42_in1), .out(andOp_42_out));

	reg [0:0] br_8_happened_in_state_1_in_data;
	wire [0:0] br_8_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_8_happened_in_state_1(.in_data(br_8_happened_in_state_1_in_data), .out_data(br_8_happened_in_state_1_out_data));

	reg [0:0] notOp_43_in0;
	wire [0:0] notOp_43_out;
	notOp #(.WIDTH(1)) notOp_43(.in(notOp_43_in0), .out(notOp_43_out));

	reg [0:0] andOp_44_in0;
	reg [0:0] andOp_44_in1;
	wire [0:0] andOp_44_out;
	andOp #(.WIDTH(1)) andOp_44(.in0(andOp_44_in0), .in1(andOp_44_in1), .out(andOp_44_out));

	reg [0:0] andOp_45_in0;
	reg [0:0] andOp_45_in1;
	wire [0:0] andOp_45_out;
	andOp #(.WIDTH(1)) andOp_45(.in0(andOp_45_in0), .in1(andOp_45_in1), .out(andOp_45_out));

	reg [0:0] br_9_happened_in_state_1_in_data;
	wire [0:0] br_9_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_9_happened_in_state_1(.in_data(br_9_happened_in_state_1_in_data), .out_data(br_9_happened_in_state_1_out_data));

	reg [0:0] notOp_46_in0;
	wire [0:0] notOp_46_out;
	notOp #(.WIDTH(1)) notOp_46(.in(notOp_46_in0), .out(notOp_46_out));

	reg [0:0] andOp_47_in0;
	reg [0:0] andOp_47_in1;
	wire [0:0] andOp_47_out;
	andOp #(.WIDTH(1)) andOp_47(.in0(andOp_47_in0), .in1(andOp_47_in1), .out(andOp_47_out));

	reg [0:0] notOp_48_in0;
	wire [0:0] notOp_48_out;
	notOp #(.WIDTH(1)) notOp_48(.in(notOp_48_in0), .out(notOp_48_out));

	reg [0:0] andOp_49_in0;
	reg [0:0] andOp_49_in1;
	wire [0:0] andOp_49_out;
	andOp #(.WIDTH(1)) andOp_49(.in0(andOp_49_in0), .in1(andOp_49_in1), .out(andOp_49_out));

	reg [0:0] andOp_50_in0;
	reg [0:0] andOp_50_in1;
	wire [0:0] andOp_50_out;
	andOp #(.WIDTH(1)) andOp_50(.in0(andOp_50_in0), .in1(andOp_50_in1), .out(andOp_50_out));

	reg [0:0] andOp_51_in0;
	reg [0:0] andOp_51_in1;
	wire [0:0] andOp_51_out;
	andOp #(.WIDTH(1)) andOp_51(.in0(andOp_51_in0), .in1(andOp_51_in1), .out(andOp_51_out));

	reg [0:0] br_10_happened_in_state_2_in_data;
	wire [0:0] br_10_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_2(.in_data(br_10_happened_in_state_2_in_data), .out_data(br_10_happened_in_state_2_out_data));

	reg [0:0] notOp_52_in0;
	wire [0:0] notOp_52_out;
	notOp #(.WIDTH(1)) notOp_52(.in(notOp_52_in0), .out(notOp_52_out));

	reg [0:0] andOp_53_in0;
	reg [0:0] andOp_53_in1;
	wire [0:0] andOp_53_out;
	andOp #(.WIDTH(1)) andOp_53(.in0(andOp_53_in0), .in1(andOp_53_in1), .out(andOp_53_out));

	reg [0:0] andOp_54_in0;
	reg [0:0] andOp_54_in1;
	wire [0:0] andOp_54_out;
	andOp #(.WIDTH(1)) andOp_54(.in0(andOp_54_in0), .in1(andOp_54_in1), .out(andOp_54_out));

	reg [0:0] br_4_happened_in_state_3_in_data;
	wire [0:0] br_4_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_3(.in_data(br_4_happened_in_state_3_in_data), .out_data(br_4_happened_in_state_3_out_data));

	reg [0:0] notOp_55_in0;
	wire [0:0] notOp_55_out;
	notOp #(.WIDTH(1)) notOp_55(.in(notOp_55_in0), .out(notOp_55_out));

	reg [0:0] andOp_56_in0;
	reg [0:0] andOp_56_in1;
	wire [0:0] andOp_56_out;
	andOp #(.WIDTH(1)) andOp_56(.in0(andOp_56_in0), .in1(andOp_56_in1), .out(andOp_56_out));

	reg [0:0] notOp_57_in0;
	wire [0:0] notOp_57_out;
	notOp #(.WIDTH(1)) notOp_57(.in(notOp_57_in0), .out(notOp_57_out));

	reg [0:0] andOp_58_in0;
	reg [0:0] andOp_58_in1;
	wire [0:0] andOp_58_out;
	andOp #(.WIDTH(1)) andOp_58(.in0(andOp_58_in0), .in1(andOp_58_in1), .out(andOp_58_out));

	reg [0:0] andOp_59_in0;
	reg [0:0] andOp_59_in1;
	wire [0:0] andOp_59_out;
	andOp #(.WIDTH(1)) andOp_59(.in0(andOp_59_in0), .in1(andOp_59_in1), .out(andOp_59_out));

	reg [0:0] andOp_60_in0;
	reg [0:0] andOp_60_in1;
	wire [0:0] andOp_60_out;
	andOp #(.WIDTH(1)) andOp_60(.in0(andOp_60_in0), .in1(andOp_60_in1), .out(andOp_60_out));

	reg [0:0] br_10_happened_in_state_3_in_data;
	wire [0:0] br_10_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_3(.in_data(br_10_happened_in_state_3_in_data), .out_data(br_10_happened_in_state_3_out_data));

	reg [0:0] notOp_61_in0;
	wire [0:0] notOp_61_out;
	notOp #(.WIDTH(1)) notOp_61(.in(notOp_61_in0), .out(notOp_61_out));

	reg [0:0] andOp_62_in0;
	reg [0:0] andOp_62_in1;
	wire [0:0] andOp_62_out;
	andOp #(.WIDTH(1)) andOp_62(.in0(andOp_62_in0), .in1(andOp_62_in1), .out(andOp_62_out));

	reg [0:0] andOp_63_in0;
	reg [0:0] andOp_63_in1;
	wire [0:0] andOp_63_out;
	andOp #(.WIDTH(1)) andOp_63(.in0(andOp_63_in0), .in1(andOp_63_in1), .out(andOp_63_out));

	reg [0:0] br_7_happened_in_state_4_in_data;
	wire [0:0] br_7_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_7_happened_in_state_4(.in_data(br_7_happened_in_state_4_in_data), .out_data(br_7_happened_in_state_4_out_data));

	reg [0:0] notOp_64_in0;
	wire [0:0] notOp_64_out;
	notOp #(.WIDTH(1)) notOp_64(.in(notOp_64_in0), .out(notOp_64_out));

	reg [0:0] andOp_65_in0;
	reg [0:0] andOp_65_in1;
	wire [0:0] andOp_65_out;
	andOp #(.WIDTH(1)) andOp_65(.in0(andOp_65_in0), .in1(andOp_65_in1), .out(andOp_65_out));

	reg [0:0] andOp_66_in0;
	reg [0:0] andOp_66_in1;
	wire [0:0] andOp_66_out;
	andOp #(.WIDTH(1)) andOp_66(.in0(andOp_66_in0), .in1(andOp_66_in1), .out(andOp_66_out));

	reg [0:0] br_6_happened_in_state_4_in_data;
	wire [0:0] br_6_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_6_happened_in_state_4(.in_data(br_6_happened_in_state_4_in_data), .out_data(br_6_happened_in_state_4_out_data));

	reg [0:0] notOp_67_in0;
	wire [0:0] notOp_67_out;
	notOp #(.WIDTH(1)) notOp_67(.in(notOp_67_in0), .out(notOp_67_out));

	reg [0:0] andOp_68_in0;
	reg [0:0] andOp_68_in1;
	wire [0:0] andOp_68_out;
	andOp #(.WIDTH(1)) andOp_68(.in0(andOp_68_in0), .in1(andOp_68_in1), .out(andOp_68_out));

	reg [0:0] notOp_69_in0;
	wire [0:0] notOp_69_out;
	notOp #(.WIDTH(1)) notOp_69(.in(notOp_69_in0), .out(notOp_69_out));

	reg [0:0] andOp_70_in0;
	reg [0:0] andOp_70_in1;
	wire [0:0] andOp_70_out;
	andOp #(.WIDTH(1)) andOp_70(.in0(andOp_70_in0), .in1(andOp_70_in1), .out(andOp_70_out));

	reg [0:0] andOp_71_in0;
	reg [0:0] andOp_71_in1;
	wire [0:0] andOp_71_out;
	andOp #(.WIDTH(1)) andOp_71(.in0(andOp_71_in0), .in1(andOp_71_in1), .out(andOp_71_out));

	reg [0:0] andOp_72_in0;
	reg [0:0] andOp_72_in1;
	wire [0:0] andOp_72_out;
	andOp #(.WIDTH(1)) andOp_72(.in0(andOp_72_in0), .in1(andOp_72_in1), .out(andOp_72_out));

	reg [0:0] br_5_happened_in_state_4_in_data;
	wire [0:0] br_5_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_5_happened_in_state_4(.in_data(br_5_happened_in_state_4_in_data), .out_data(br_5_happened_in_state_4_out_data));

	reg [0:0] notOp_73_in0;
	wire [0:0] notOp_73_out;
	notOp #(.WIDTH(1)) notOp_73(.in(notOp_73_in0), .out(notOp_73_out));

	reg [0:0] andOp_74_in0;
	reg [0:0] andOp_74_in1;
	wire [0:0] andOp_74_out;
	andOp #(.WIDTH(1)) andOp_74(.in0(andOp_74_in0), .in1(andOp_74_in1), .out(andOp_74_out));

	reg [0:0] andOp_75_in0;
	reg [0:0] andOp_75_in1;
	wire [0:0] andOp_75_out;
	andOp #(.WIDTH(1)) andOp_75(.in0(andOp_75_in0), .in1(andOp_75_in1), .out(andOp_75_out));

	reg [0:0] br_4_happened_in_state_4_in_data;
	wire [0:0] br_4_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_4(.in_data(br_4_happened_in_state_4_in_data), .out_data(br_4_happened_in_state_4_out_data));

	reg [0:0] notOp_76_in0;
	wire [0:0] notOp_76_out;
	notOp #(.WIDTH(1)) notOp_76(.in(notOp_76_in0), .out(notOp_76_out));

	reg [0:0] andOp_77_in0;
	reg [0:0] andOp_77_in1;
	wire [0:0] andOp_77_out;
	andOp #(.WIDTH(1)) andOp_77(.in0(andOp_77_in0), .in1(andOp_77_in1), .out(andOp_77_out));

	reg [0:0] notOp_78_in0;
	wire [0:0] notOp_78_out;
	notOp #(.WIDTH(1)) notOp_78(.in(notOp_78_in0), .out(notOp_78_out));

	reg [0:0] andOp_79_in0;
	reg [0:0] andOp_79_in1;
	wire [0:0] andOp_79_out;
	andOp #(.WIDTH(1)) andOp_79(.in0(andOp_79_in0), .in1(andOp_79_in1), .out(andOp_79_out));

	reg [0:0] andOp_80_in0;
	reg [0:0] andOp_80_in1;
	wire [0:0] andOp_80_out;
	andOp #(.WIDTH(1)) andOp_80(.in0(andOp_80_in0), .in1(andOp_80_in1), .out(andOp_80_out));

	reg [0:0] andOp_81_in0;
	reg [0:0] andOp_81_in1;
	wire [0:0] andOp_81_out;
	andOp #(.WIDTH(1)) andOp_81(.in0(andOp_81_in0), .in1(andOp_81_in1), .out(andOp_81_out));

	reg [0:0] br_1_happened_in_state_4_in_data;
	wire [0:0] br_1_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened_in_state_4(.in_data(br_1_happened_in_state_4_in_data), .out_data(br_1_happened_in_state_4_out_data));

	reg [0:0] notOp_82_in0;
	wire [0:0] notOp_82_out;
	notOp #(.WIDTH(1)) notOp_82(.in(notOp_82_in0), .out(notOp_82_out));

	reg [31:0] eq_83_in0;
	reg [31:0] eq_83_in1;
	wire [0:0] eq_83_out;
	eq #(.WIDTH(32)) eq_83(.in0(eq_83_in0), .in1(eq_83_in1), .out(eq_83_out));

	reg [31:0] eq_84_in0;
	reg [31:0] eq_84_in1;
	wire [0:0] eq_84_out;
	eq #(.WIDTH(32)) eq_84(.in0(eq_84_in0), .in1(eq_84_in1), .out(eq_84_out));

	reg [31:0] eq_85_in0;
	reg [31:0] eq_85_in1;
	wire [0:0] eq_85_out;
	eq #(.WIDTH(32)) eq_85(.in0(eq_85_in0), .in1(eq_85_in1), .out(eq_85_out));

	reg [0:0] orOp_86_in0;
	reg [0:0] orOp_86_in1;
	wire [0:0] orOp_86_out;
	orOp #(.WIDTH(1)) orOp_86(.in0(orOp_86_in0), .in1(orOp_86_in1), .out(orOp_86_out));

	reg [31:0] eq_87_in0;
	reg [31:0] eq_87_in1;
	wire [0:0] eq_87_out;
	eq #(.WIDTH(32)) eq_87(.in0(eq_87_in0), .in1(eq_87_in1), .out(eq_87_out));

	reg [0:0] orOp_88_in0;
	reg [0:0] orOp_88_in1;
	wire [0:0] orOp_88_out;
	orOp #(.WIDTH(1)) orOp_88(.in0(orOp_88_in0), .in1(orOp_88_in1), .out(orOp_88_out));

	reg [31:0] eq_89_in0;
	reg [31:0] eq_89_in1;
	wire [0:0] eq_89_out;
	eq #(.WIDTH(32)) eq_89(.in0(eq_89_in0), .in1(eq_89_in1), .out(eq_89_out));

	reg [0:0] orOp_90_in0;
	reg [0:0] orOp_90_in1;
	wire [0:0] orOp_90_out;
	orOp #(.WIDTH(1)) orOp_90(.in0(orOp_90_in0), .in1(orOp_90_in1), .out(orOp_90_out));

	reg [31:0] eq_91_in0;
	reg [31:0] eq_91_in1;
	wire [0:0] eq_91_out;
	eq #(.WIDTH(32)) eq_91(.in0(eq_91_in0), .in1(eq_91_in1), .out(eq_91_out));

	reg [31:0] eq_92_in0;
	reg [31:0] eq_92_in1;
	wire [0:0] eq_92_out;
	eq #(.WIDTH(32)) eq_92(.in0(eq_92_in0), .in1(eq_92_in1), .out(eq_92_out));

	reg [0:0] orOp_93_in0;
	reg [0:0] orOp_93_in1;
	wire [0:0] orOp_93_out;
	orOp #(.WIDTH(1)) orOp_93(.in0(orOp_93_in0), .in1(orOp_93_in1), .out(orOp_93_out));

	reg [31:0] eq_94_in0;
	reg [31:0] eq_94_in1;
	wire [0:0] eq_94_out;
	eq #(.WIDTH(32)) eq_94(.in0(eq_94_in0), .in1(eq_94_in1), .out(eq_94_out));

	reg [31:0] eq_95_in0;
	reg [31:0] eq_95_in1;
	wire [0:0] eq_95_out;
	eq #(.WIDTH(32)) eq_95(.in0(eq_95_in0), .in1(eq_95_in1), .out(eq_95_out));

	reg [0:0] orOp_96_in0;
	reg [0:0] orOp_96_in1;
	wire [0:0] orOp_96_out;
	orOp #(.WIDTH(1)) orOp_96(.in0(orOp_96_in0), .in1(orOp_96_in1), .out(orOp_96_out));

	reg [31:0] eq_97_in0;
	reg [31:0] eq_97_in1;
	wire [0:0] eq_97_out;
	eq #(.WIDTH(32)) eq_97(.in0(eq_97_in0), .in1(eq_97_in1), .out(eq_97_out));

	reg [0:0] orOp_98_in0;
	reg [0:0] orOp_98_in1;
	wire [0:0] orOp_98_out;
	orOp #(.WIDTH(1)) orOp_98(.in0(orOp_98_in0), .in1(orOp_98_in1), .out(orOp_98_out));

	reg [31:0] eq_99_in0;
	reg [31:0] eq_99_in1;
	wire [0:0] eq_99_out;
	eq #(.WIDTH(32)) eq_99(.in0(eq_99_in0), .in1(eq_99_in1), .out(eq_99_out));

	reg [0:0] orOp_100_in0;
	reg [0:0] orOp_100_in1;
	wire [0:0] orOp_100_out;
	orOp #(.WIDTH(1)) orOp_100(.in0(orOp_100_in0), .in1(orOp_100_in1), .out(orOp_100_out));

	reg [31:0] eq_101_in0;
	reg [31:0] eq_101_in1;
	wire [0:0] eq_101_out;
	eq #(.WIDTH(32)) eq_101(.in0(eq_101_in0), .in1(eq_101_in1), .out(eq_101_out));

	reg [31:0] eq_102_in0;
	reg [31:0] eq_102_in1;
	wire [0:0] eq_102_out;
	eq #(.WIDTH(32)) eq_102(.in0(eq_102_in0), .in1(eq_102_in1), .out(eq_102_out));

	reg [0:0] orOp_103_in0;
	reg [0:0] orOp_103_in1;
	wire [0:0] orOp_103_out;
	orOp #(.WIDTH(1)) orOp_103(.in0(orOp_103_in0), .in1(orOp_103_in1), .out(orOp_103_out));

	reg [31:0] eq_104_in0;
	reg [31:0] eq_104_in1;
	wire [0:0] eq_104_out;
	eq #(.WIDTH(32)) eq_104(.in0(eq_104_in0), .in1(eq_104_in1), .out(eq_104_out));

	reg [0:0] orOp_105_in0;
	reg [0:0] orOp_105_in1;
	wire [0:0] orOp_105_out;
	orOp #(.WIDTH(1)) orOp_105(.in0(orOp_105_in0), .in1(orOp_105_in1), .out(orOp_105_out));

	reg [31:0] eq_106_in0;
	reg [31:0] eq_106_in1;
	wire [0:0] eq_106_out;
	eq #(.WIDTH(32)) eq_106(.in0(eq_106_in0), .in1(eq_106_in1), .out(eq_106_out));

	reg [31:0] eq_107_in0;
	reg [31:0] eq_107_in1;
	wire [0:0] eq_107_out;
	eq #(.WIDTH(32)) eq_107(.in0(eq_107_in0), .in1(eq_107_in1), .out(eq_107_out));

	reg [31:0] eq_108_in0;
	reg [31:0] eq_108_in1;
	wire [0:0] eq_108_out;
	eq #(.WIDTH(32)) eq_108(.in0(eq_108_in0), .in1(eq_108_in1), .out(eq_108_out));

	reg [0:0] notOp_109_in0;
	wire [0:0] notOp_109_out;
	notOp #(.WIDTH(1)) notOp_109(.in(notOp_109_in0), .out(notOp_109_out));

	reg [0:0] andOp_110_in0;
	reg [0:0] andOp_110_in1;
	wire [0:0] andOp_110_out;
	andOp #(.WIDTH(1)) andOp_110(.in0(andOp_110_in0), .in1(andOp_110_in1), .out(andOp_110_out));

	reg [31:0] eq_111_in0;
	reg [31:0] eq_111_in1;
	wire [0:0] eq_111_out;
	eq #(.WIDTH(32)) eq_111(.in0(eq_111_in0), .in1(eq_111_in1), .out(eq_111_out));

	reg [0:0] notOp_112_in0;
	wire [0:0] notOp_112_out;
	notOp #(.WIDTH(1)) notOp_112(.in(notOp_112_in0), .out(notOp_112_out));

	reg [0:0] andOp_113_in0;
	reg [0:0] andOp_113_in1;
	wire [0:0] andOp_113_out;
	andOp #(.WIDTH(1)) andOp_113(.in0(andOp_113_in0), .in1(andOp_113_in1), .out(andOp_113_out));

	reg [31:0] eq_114_in0;
	reg [31:0] eq_114_in1;
	wire [0:0] eq_114_out;
	eq #(.WIDTH(32)) eq_114(.in0(eq_114_in0), .in1(eq_114_in1), .out(eq_114_out));

	reg [0:0] notOp_115_in0;
	wire [0:0] notOp_115_out;
	notOp #(.WIDTH(1)) notOp_115(.in(notOp_115_in0), .out(notOp_115_out));

	reg [0:0] andOp_116_in0;
	reg [0:0] andOp_116_in1;
	wire [0:0] andOp_116_out;
	andOp #(.WIDTH(1)) andOp_116(.in0(andOp_116_in0), .in1(andOp_116_in1), .out(andOp_116_out));

	reg [31:0] eq_117_in0;
	reg [31:0] eq_117_in1;
	wire [0:0] eq_117_out;
	eq #(.WIDTH(32)) eq_117(.in0(eq_117_in0), .in1(eq_117_in1), .out(eq_117_out));

	reg [31:0] eq_118_in0;
	reg [31:0] eq_118_in1;
	wire [0:0] eq_118_out;
	eq #(.WIDTH(32)) eq_118(.in0(eq_118_in0), .in1(eq_118_in1), .out(eq_118_out));

	reg [0:0] notOp_119_in0;
	wire [0:0] notOp_119_out;
	notOp #(.WIDTH(1)) notOp_119(.in(notOp_119_in0), .out(notOp_119_out));

	reg [0:0] andOp_120_in0;
	reg [0:0] andOp_120_in1;
	wire [0:0] andOp_120_out;
	andOp #(.WIDTH(1)) andOp_120(.in0(andOp_120_in0), .in1(andOp_120_in1), .out(andOp_120_out));

	reg [31:0] eq_121_in0;
	reg [31:0] eq_121_in1;
	wire [0:0] eq_121_out;
	eq #(.WIDTH(32)) eq_121(.in0(eq_121_in0), .in1(eq_121_in1), .out(eq_121_out));

	reg [31:0] eq_122_in0;
	reg [31:0] eq_122_in1;
	wire [0:0] eq_122_out;
	eq #(.WIDTH(32)) eq_122(.in0(eq_122_in0), .in1(eq_122_in1), .out(eq_122_out));

	reg [0:0] notOp_123_in0;
	wire [0:0] notOp_123_out;
	notOp #(.WIDTH(1)) notOp_123(.in(notOp_123_in0), .out(notOp_123_out));

	reg [0:0] andOp_124_in0;
	reg [0:0] andOp_124_in1;
	wire [0:0] andOp_124_out;
	andOp #(.WIDTH(1)) andOp_124(.in0(andOp_124_in0), .in1(andOp_124_in1), .out(andOp_124_out));

	reg [31:0] eq_125_in0;
	reg [31:0] eq_125_in1;
	wire [0:0] eq_125_out;
	eq #(.WIDTH(32)) eq_125(.in0(eq_125_in0), .in1(eq_125_in1), .out(eq_125_out));

	reg [0:0] notOp_126_in0;
	wire [0:0] notOp_126_out;
	notOp #(.WIDTH(1)) notOp_126(.in(notOp_126_in0), .out(notOp_126_out));

	reg [0:0] andOp_127_in0;
	reg [0:0] andOp_127_in1;
	wire [0:0] andOp_127_out;
	andOp #(.WIDTH(1)) andOp_127(.in0(andOp_127_in0), .in1(andOp_127_in1), .out(andOp_127_out));

	reg [31:0] eq_128_in0;
	reg [31:0] eq_128_in1;
	wire [0:0] eq_128_out;
	eq #(.WIDTH(32)) eq_128(.in0(eq_128_in0), .in1(eq_128_in1), .out(eq_128_out));

	reg [0:0] notOp_129_in0;
	wire [0:0] notOp_129_out;
	notOp #(.WIDTH(1)) notOp_129(.in(notOp_129_in0), .out(notOp_129_out));

	reg [0:0] andOp_130_in0;
	reg [0:0] andOp_130_in1;
	wire [0:0] andOp_130_out;
	andOp #(.WIDTH(1)) andOp_130(.in0(andOp_130_in0), .in1(andOp_130_in1), .out(andOp_130_out));

	reg [31:0] eq_131_in0;
	reg [31:0] eq_131_in1;
	wire [0:0] eq_131_out;
	eq #(.WIDTH(32)) eq_131(.in0(eq_131_in0), .in1(eq_131_in1), .out(eq_131_out));

	reg [31:0] eq_132_in0;
	reg [31:0] eq_132_in1;
	wire [0:0] eq_132_out;
	eq #(.WIDTH(32)) eq_132(.in0(eq_132_in0), .in1(eq_132_in1), .out(eq_132_out));

	reg [0:0] notOp_133_in0;
	wire [0:0] notOp_133_out;
	notOp #(.WIDTH(1)) notOp_133(.in(notOp_133_in0), .out(notOp_133_out));

	reg [0:0] andOp_134_in0;
	reg [0:0] andOp_134_in1;
	wire [0:0] andOp_134_out;
	andOp #(.WIDTH(1)) andOp_134(.in0(andOp_134_in0), .in1(andOp_134_in1), .out(andOp_134_out));

	reg [31:0] eq_135_in0;
	reg [31:0] eq_135_in1;
	wire [0:0] eq_135_out;
	eq #(.WIDTH(32)) eq_135(.in0(eq_135_in0), .in1(eq_135_in1), .out(eq_135_out));

	reg [0:0] notOp_136_in0;
	wire [0:0] notOp_136_out;
	notOp #(.WIDTH(1)) notOp_136(.in(notOp_136_in0), .out(notOp_136_out));

	reg [0:0] andOp_137_in0;
	reg [0:0] andOp_137_in1;
	wire [0:0] andOp_137_out;
	andOp #(.WIDTH(1)) andOp_137(.in0(andOp_137_in0), .in1(andOp_137_in1), .out(andOp_137_out));

	reg [0:0] andOp_138_in0;
	reg [0:0] andOp_138_in1;
	wire [0:0] andOp_138_out;
	andOp #(.WIDTH(1)) andOp_138(.in0(andOp_138_in0), .in1(andOp_138_in1), .out(andOp_138_out));

	reg [0:0] andOp_139_in0;
	reg [0:0] andOp_139_in1;
	wire [0:0] andOp_139_out;
	andOp #(.WIDTH(1)) andOp_139(.in0(andOp_139_in0), .in1(andOp_139_in1), .out(andOp_139_out));

	reg [0:0] andOp_140_in0;
	reg [0:0] andOp_140_in1;
	wire [0:0] andOp_140_out;
	andOp #(.WIDTH(1)) andOp_140(.in0(andOp_140_in0), .in1(andOp_140_in1), .out(andOp_140_out));

	reg [0:0] andOp_141_in0;
	reg [0:0] andOp_141_in1;
	wire [0:0] andOp_141_out;
	andOp #(.WIDTH(1)) andOp_141(.in0(andOp_141_in0), .in1(andOp_141_in1), .out(andOp_141_out));

	reg [0:0] andOp_142_in0;
	reg [0:0] andOp_142_in1;
	wire [0:0] andOp_142_out;
	andOp #(.WIDTH(1)) andOp_142(.in0(andOp_142_in0), .in1(andOp_142_in1), .out(andOp_142_out));

	reg [0:0] andOp_143_in0;
	reg [0:0] andOp_143_in1;
	wire [0:0] andOp_143_out;
	andOp #(.WIDTH(1)) andOp_143(.in0(andOp_143_in0), .in1(andOp_143_in1), .out(andOp_143_out));

	reg [0:0] andOp_144_in0;
	reg [0:0] andOp_144_in1;
	wire [0:0] andOp_144_out;
	andOp #(.WIDTH(1)) andOp_144(.in0(andOp_144_in0), .in1(andOp_144_in1), .out(andOp_144_out));

	reg [0:0] andOp_145_in0;
	reg [0:0] andOp_145_in1;
	wire [0:0] andOp_145_out;
	andOp #(.WIDTH(1)) andOp_145(.in0(andOp_145_in0), .in1(andOp_145_in1), .out(andOp_145_out));

	reg [0:0] andOp_146_in0;
	reg [0:0] andOp_146_in1;
	wire [0:0] andOp_146_out;
	andOp #(.WIDTH(1)) andOp_146(.in0(andOp_146_in0), .in1(andOp_146_in1), .out(andOp_146_out));

	reg [0:0] andOp_147_in0;
	reg [0:0] andOp_147_in1;
	wire [0:0] andOp_147_out;
	andOp #(.WIDTH(1)) andOp_147(.in0(andOp_147_in0), .in1(andOp_147_in1), .out(andOp_147_out));

	reg [0:0] andOp_148_in0;
	reg [0:0] andOp_148_in1;
	wire [0:0] andOp_148_out;
	andOp #(.WIDTH(1)) andOp_148(.in0(andOp_148_in0), .in1(andOp_148_in1), .out(andOp_148_out));

	reg [31:0] concat_149_in0;
	reg [31:0] concat_149_in1;
	wire [63:0] concat_149_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_149(.in0(concat_149_in0), .in1(concat_149_in1), .out(concat_149_out));

	reg [31:0] concat_150_in0;
	reg [31:0] concat_150_in1;
	wire [63:0] concat_150_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_150(.in0(concat_150_in0), .in1(concat_150_in1), .out(concat_150_out));

	reg [0:0] andOp_151_in0;
	reg [0:0] andOp_151_in1;
	wire [0:0] andOp_151_out;
	andOp #(.WIDTH(1)) andOp_151(.in0(andOp_151_in0), .in1(andOp_151_in1), .out(andOp_151_out));

	reg [31:0] tmp_output_152_in_data;
	wire [31:0] tmp_output_152_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_152(.in_data(tmp_output_152_in_data), .out_data(tmp_output_152_out_data));

	reg [31:0] eq_153_in0;
	reg [31:0] eq_153_in1;
	wire [0:0] eq_153_out;
	eq #(.WIDTH(32)) eq_153(.in0(eq_153_in0), .in1(eq_153_in1), .out(eq_153_out));

	reg [0:0] andOp_154_in0;
	reg [0:0] andOp_154_in1;
	wire [0:0] andOp_154_out;
	andOp #(.WIDTH(1)) andOp_154(.in0(andOp_154_in0), .in1(andOp_154_in1), .out(andOp_154_out));

	reg [0:0] andOp_155_in0;
	reg [0:0] andOp_155_in1;
	wire [0:0] andOp_155_out;
	andOp #(.WIDTH(1)) andOp_155(.in0(andOp_155_in0), .in1(andOp_155_in1), .out(andOp_155_out));

	reg [0:0] andOp_156_in0;
	reg [0:0] andOp_156_in1;
	wire [0:0] andOp_156_out;
	andOp #(.WIDTH(1)) andOp_156(.in0(andOp_156_in0), .in1(andOp_156_in1), .out(andOp_156_out));

	reg [0:0] andOp_157_in0;
	reg [0:0] andOp_157_in1;
	wire [0:0] andOp_157_out;
	andOp #(.WIDTH(1)) andOp_157(.in0(andOp_157_in0), .in1(andOp_157_in1), .out(andOp_157_out));

	reg [0:0] andOp_158_in0;
	reg [0:0] andOp_158_in1;
	wire [0:0] andOp_158_out;
	andOp #(.WIDTH(1)) andOp_158(.in0(andOp_158_in0), .in1(andOp_158_in1), .out(andOp_158_out));

	reg [0:0] andOp_159_in0;
	reg [0:0] andOp_159_in1;
	wire [0:0] andOp_159_out;
	andOp #(.WIDTH(1)) andOp_159(.in0(andOp_159_in0), .in1(andOp_159_in1), .out(andOp_159_out));

	reg [0:0] andOp_160_in0;
	reg [0:0] andOp_160_in1;
	wire [0:0] andOp_160_out;
	andOp #(.WIDTH(1)) andOp_160(.in0(andOp_160_in0), .in1(andOp_160_in1), .out(andOp_160_out));

	reg [0:0] andOp_161_in0;
	reg [0:0] andOp_161_in1;
	wire [0:0] andOp_161_out;
	andOp #(.WIDTH(1)) andOp_161(.in0(andOp_161_in0), .in1(andOp_161_in1), .out(andOp_161_out));

	reg [0:0] andOp_162_in0;
	reg [0:0] andOp_162_in1;
	wire [0:0] andOp_162_out;
	andOp #(.WIDTH(1)) andOp_162(.in0(andOp_162_in0), .in1(andOp_162_in1), .out(andOp_162_out));

	reg [0:0] andOp_163_in0;
	reg [0:0] andOp_163_in1;
	wire [0:0] andOp_163_out;
	andOp #(.WIDTH(1)) andOp_163(.in0(andOp_163_in0), .in1(andOp_163_in1), .out(andOp_163_out));

	reg [0:0] andOp_164_in0;
	reg [0:0] andOp_164_in1;
	wire [0:0] andOp_164_out;
	andOp #(.WIDTH(1)) andOp_164(.in0(andOp_164_in0), .in1(andOp_164_in1), .out(andOp_164_out));

	reg [0:0] notOp_165_in0;
	wire [0:0] notOp_165_out;
	notOp #(.WIDTH(1)) notOp_165(.in(notOp_165_in0), .out(notOp_165_out));

	reg [0:0] andOp_166_in0;
	reg [0:0] andOp_166_in1;
	wire [0:0] andOp_166_out;
	andOp #(.WIDTH(1)) andOp_166(.in0(andOp_166_in0), .in1(andOp_166_in1), .out(andOp_166_out));

	reg [0:0] notOp_167_in0;
	wire [0:0] notOp_167_out;
	notOp #(.WIDTH(1)) notOp_167(.in(notOp_167_in0), .out(notOp_167_out));

	reg [0:0] andOp_168_in0;
	reg [0:0] andOp_168_in1;
	wire [0:0] andOp_168_out;
	andOp #(.WIDTH(1)) andOp_168(.in0(andOp_168_in0), .in1(andOp_168_in1), .out(andOp_168_out));

	reg [0:0] notOp_169_in0;
	wire [0:0] notOp_169_out;
	notOp #(.WIDTH(1)) notOp_169(.in(notOp_169_in0), .out(notOp_169_out));

	reg [0:0] andOp_170_in0;
	reg [0:0] andOp_170_in1;
	wire [0:0] andOp_170_out;
	andOp #(.WIDTH(1)) andOp_170(.in0(andOp_170_in0), .in1(andOp_170_in1), .out(andOp_170_out));

	reg [0:0] notOp_171_in0;
	wire [0:0] notOp_171_out;
	notOp #(.WIDTH(1)) notOp_171(.in(notOp_171_in0), .out(notOp_171_out));

	reg [0:0] andOp_172_in0;
	reg [0:0] andOp_172_in1;
	wire [0:0] andOp_172_out;
	andOp #(.WIDTH(1)) andOp_172(.in0(andOp_172_in0), .in1(andOp_172_in1), .out(andOp_172_out));

	reg [0:0] notOp_173_in0;
	wire [0:0] notOp_173_out;
	notOp #(.WIDTH(1)) notOp_173(.in(notOp_173_in0), .out(notOp_173_out));

	reg [0:0] andOp_174_in0;
	reg [0:0] andOp_174_in1;
	wire [0:0] andOp_174_out;
	andOp #(.WIDTH(1)) andOp_174(.in0(andOp_174_in0), .in1(andOp_174_in1), .out(andOp_174_out));

	reg [0:0] notOp_175_in0;
	wire [0:0] notOp_175_out;
	notOp #(.WIDTH(1)) notOp_175(.in(notOp_175_in0), .out(notOp_175_out));

	reg [0:0] andOp_176_in0;
	reg [0:0] andOp_176_in1;
	wire [0:0] andOp_176_out;
	andOp #(.WIDTH(1)) andOp_176(.in0(andOp_176_in0), .in1(andOp_176_in1), .out(andOp_176_out));

	reg [0:0] notOp_177_in0;
	wire [0:0] notOp_177_out;
	notOp #(.WIDTH(1)) notOp_177(.in(notOp_177_in0), .out(notOp_177_out));

	reg [0:0] andOp_178_in0;
	reg [0:0] andOp_178_in1;
	wire [0:0] andOp_178_out;
	andOp #(.WIDTH(1)) andOp_178(.in0(andOp_178_in0), .in1(andOp_178_in1), .out(andOp_178_out));

	reg [0:0] notOp_179_in0;
	wire [0:0] notOp_179_out;
	notOp #(.WIDTH(1)) notOp_179(.in(notOp_179_in0), .out(notOp_179_out));

	reg [0:0] andOp_180_in0;
	reg [0:0] andOp_180_in1;
	wire [0:0] andOp_180_out;
	andOp #(.WIDTH(1)) andOp_180(.in0(andOp_180_in0), .in1(andOp_180_in1), .out(andOp_180_out));

	reg [31:0] eq_181_in0;
	reg [31:0] eq_181_in1;
	wire [0:0] eq_181_out;
	eq #(.WIDTH(32)) eq_181(.in0(eq_181_in0), .in1(eq_181_in1), .out(eq_181_out));

	reg [31:0] eq_182_in0;
	reg [31:0] eq_182_in1;
	wire [0:0] eq_182_out;
	eq #(.WIDTH(32)) eq_182(.in0(eq_182_in0), .in1(eq_182_in1), .out(eq_182_out));

	reg [31:0] eq_183_in0;
	reg [31:0] eq_183_in1;
	wire [0:0] eq_183_out;
	eq #(.WIDTH(32)) eq_183(.in0(eq_183_in0), .in1(eq_183_in1), .out(eq_183_out));

	reg [31:0] eq_184_in0;
	reg [31:0] eq_184_in1;
	wire [0:0] eq_184_out;
	eq #(.WIDTH(32)) eq_184(.in0(eq_184_in0), .in1(eq_184_in1), .out(eq_184_out));

	reg [0:0] andOp_185_in0;
	reg [0:0] andOp_185_in1;
	wire [0:0] andOp_185_out;
	andOp #(.WIDTH(1)) andOp_185(.in0(andOp_185_in0), .in1(andOp_185_in1), .out(andOp_185_out));

	reg [0:0] andOp_186_in0;
	reg [0:0] andOp_186_in1;
	wire [0:0] andOp_186_out;
	andOp #(.WIDTH(1)) andOp_186(.in0(andOp_186_in0), .in1(andOp_186_in1), .out(andOp_186_out));

	reg [31:0] eq_187_in0;
	reg [31:0] eq_187_in1;
	wire [0:0] eq_187_out;
	eq #(.WIDTH(32)) eq_187(.in0(eq_187_in0), .in1(eq_187_in1), .out(eq_187_out));

	reg [31:0] eq_188_in0;
	reg [31:0] eq_188_in1;
	wire [0:0] eq_188_out;
	eq #(.WIDTH(32)) eq_188(.in0(eq_188_in0), .in1(eq_188_in1), .out(eq_188_out));

	reg [31:0] eq_189_in0;
	reg [31:0] eq_189_in1;
	wire [0:0] eq_189_out;
	eq #(.WIDTH(32)) eq_189(.in0(eq_189_in0), .in1(eq_189_in1), .out(eq_189_out));

	reg [31:0] eq_190_in0;
	reg [31:0] eq_190_in1;
	wire [0:0] eq_190_out;
	eq #(.WIDTH(32)) eq_190(.in0(eq_190_in0), .in1(eq_190_in1), .out(eq_190_out));

	reg [0:0] andOp_191_in0;
	reg [0:0] andOp_191_in1;
	wire [0:0] andOp_191_out;
	andOp #(.WIDTH(1)) andOp_191(.in0(andOp_191_in0), .in1(andOp_191_in1), .out(andOp_191_out));

	reg [0:0] andOp_192_in0;
	reg [0:0] andOp_192_in1;
	wire [0:0] andOp_192_out;
	andOp #(.WIDTH(1)) andOp_192(.in0(andOp_192_in0), .in1(andOp_192_in1), .out(andOp_192_out));

	reg [0:0] andOp_193_in0;
	reg [0:0] andOp_193_in1;
	wire [0:0] andOp_193_out;
	andOp #(.WIDTH(1)) andOp_193(.in0(andOp_193_in0), .in1(andOp_193_in1), .out(andOp_193_out));

	reg [0:0] andOp_194_in0;
	reg [0:0] andOp_194_in1;
	wire [0:0] andOp_194_out;
	andOp #(.WIDTH(1)) andOp_194(.in0(andOp_194_in0), .in1(andOp_194_in1), .out(andOp_194_out));

	reg [0:0] andOp_195_in0;
	reg [0:0] andOp_195_in1;
	wire [0:0] andOp_195_out;
	andOp #(.WIDTH(1)) andOp_195(.in0(andOp_195_in0), .in1(andOp_195_in1), .out(andOp_195_out));

	reg [0:0] andOp_196_in0;
	reg [0:0] andOp_196_in1;
	wire [0:0] andOp_196_out;
	andOp #(.WIDTH(1)) andOp_196(.in0(andOp_196_in0), .in1(andOp_196_in1), .out(andOp_196_out));

	reg [31:0] eq_197_in0;
	reg [31:0] eq_197_in1;
	wire [0:0] eq_197_out;
	eq #(.WIDTH(32)) eq_197(.in0(eq_197_in0), .in1(eq_197_in1), .out(eq_197_out));

	reg [31:0] eq_198_in0;
	reg [31:0] eq_198_in1;
	wire [0:0] eq_198_out;
	eq #(.WIDTH(32)) eq_198(.in0(eq_198_in0), .in1(eq_198_in1), .out(eq_198_out));

	// End Functional Units

	reg [31:0] data_store_1_0;
	reg [31:0] data_store_1_2;
	reg [31:0] data_store_1_4;
	reg [0:0] data_store_1_6;
	reg [31:0] data_store_2_10;
	reg [31:0] data_store_2_12;
	reg [0:0] data_store_2_14;
	reg [31:0] data_store_2_8;
	reg [31:0] data_store_3_16;
	reg [31:0] data_store_3_18;
	reg [31:0] data_store_3_20;
	reg [0:0] data_store_3_22;
	reg [31:0] data_store_4_24;
	reg [31:0] data_store_4_26;
	reg [31:0] data_store_4_28;
	reg [0:0] data_store_4_30;
	reg [31:0] global_state;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_3_last_state;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;
	reg [31:0] state_4_last_state;

	// controller for add_add_14.add_in0_add_14
	// controller for add_add_14.add_in1_add_14
	// Insensitive connections
	always @(*) begin
		add_in0_add_14 = valid ? rdata_ram_0 : rdata_ram_0;
		add_in1_add_14 = valid ? tmp_output_152_out_data : tmp_output_152_out_data;
	end
	// controller for add_add_16.add_in0_add_16
	// controller for add_add_16.add_in1_add_16
	// Insensitive connections
	always @(*) begin
		add_in0_add_16 = valid ? data_in_3_19_out_data : data_in_3_19_out_data;
		add_in1_add_16 = valid ? 32'd1 : 32'd1;
	end
	// controller for andOp_110.andOp_110_in0
	// controller for andOp_110.andOp_110_in1
	// Insensitive connections
	always @(*) begin
		andOp_110_in0 = valid ? notOp_109_out : notOp_109_out;
		andOp_110_in1 = valid ? andOp_33_out : andOp_33_out;
	end
	// controller for andOp_113.andOp_113_in0
	// controller for andOp_113.andOp_113_in1
	// Insensitive connections
	always @(*) begin
		andOp_113_in0 = valid ? notOp_112_out : notOp_112_out;
		andOp_113_in1 = valid ? andOp_39_out : andOp_39_out;
	end
	// controller for andOp_116.andOp_116_in0
	// controller for andOp_116.andOp_116_in1
	// Insensitive connections
	always @(*) begin
		andOp_116_in0 = valid ? notOp_115_out : notOp_115_out;
		andOp_116_in1 = valid ? andOp_42_out : andOp_42_out;
	end
	// controller for andOp_120.andOp_120_in0
	// controller for andOp_120.andOp_120_in1
	// Insensitive connections
	always @(*) begin
		andOp_120_in0 = valid ? notOp_119_out : notOp_119_out;
		andOp_120_in1 = valid ? andOp_51_out : andOp_51_out;
	end
	// controller for andOp_124.andOp_124_in0
	// controller for andOp_124.andOp_124_in1
	// Insensitive connections
	always @(*) begin
		andOp_124_in0 = valid ? notOp_123_out : notOp_123_out;
		andOp_124_in1 = valid ? andOp_68_out : andOp_68_out;
	end
	// controller for andOp_127.andOp_127_in0
	// controller for andOp_127.andOp_127_in1
	// Insensitive connections
	always @(*) begin
		andOp_127_in0 = valid ? notOp_126_out : notOp_126_out;
		andOp_127_in1 = valid ? andOp_72_out : andOp_72_out;
	end
	// controller for andOp_130.andOp_130_in0
	// controller for andOp_130.andOp_130_in1
	// Insensitive connections
	always @(*) begin
		andOp_130_in0 = valid ? notOp_129_out : notOp_129_out;
		andOp_130_in1 = valid ? andOp_81_out : andOp_81_out;
	end
	// controller for andOp_134.andOp_134_in0
	// controller for andOp_134.andOp_134_in1
	// Insensitive connections
	always @(*) begin
		andOp_134_in0 = valid ? notOp_133_out : notOp_133_out;
		andOp_134_in1 = valid ? andOp_63_out : andOp_63_out;
	end
	// controller for andOp_137.andOp_137_in0
	// controller for andOp_137.andOp_137_in1
	// Insensitive connections
	always @(*) begin
		andOp_137_in0 = valid ? notOp_136_out : notOp_136_out;
		andOp_137_in1 = valid ? andOp_56_out : andOp_56_out;
	end
	// controller for andOp_138.andOp_138_in0
	// controller for andOp_138.andOp_138_in1
	// Insensitive connections
	always @(*) begin
		andOp_138_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_138_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_139.andOp_139_in0
	// controller for andOp_139.andOp_139_in1
	// Insensitive connections
	always @(*) begin
		andOp_139_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_139_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_140.andOp_140_in0
	// controller for andOp_140.andOp_140_in1
	// Insensitive connections
	always @(*) begin
		andOp_140_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_140_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_141.andOp_141_in0
	// controller for andOp_141.andOp_141_in1
	// Insensitive connections
	always @(*) begin
		andOp_141_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_141_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_142.andOp_142_in0
	// controller for andOp_142.andOp_142_in1
	// Insensitive connections
	always @(*) begin
		andOp_142_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_142_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_143.andOp_143_in0
	// controller for andOp_143.andOp_143_in1
	// Insensitive connections
	always @(*) begin
		andOp_143_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_143_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_144.andOp_144_in0
	// controller for andOp_144.andOp_144_in1
	// Insensitive connections
	always @(*) begin
		andOp_144_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_144_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_145.andOp_145_in0
	// controller for andOp_145.andOp_145_in1
	// Insensitive connections
	always @(*) begin
		andOp_145_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
		andOp_145_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_146.andOp_146_in0
	// controller for andOp_146.andOp_146_in1
	// Insensitive connections
	always @(*) begin
		andOp_146_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_146_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_147.andOp_147_in0
	// controller for andOp_147.andOp_147_in1
	// Insensitive connections
	always @(*) begin
		andOp_147_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_147_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_148.andOp_148_in0
	// controller for andOp_148.andOp_148_in1
	// Insensitive connections
	always @(*) begin
		andOp_148_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_148_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_151.andOp_151_in0
	// controller for andOp_151.andOp_151_in1
	// Insensitive connections
	always @(*) begin
		andOp_151_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_151_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_154.andOp_154_in0
	// controller for andOp_154.andOp_154_in1
	// Insensitive connections
	always @(*) begin
		andOp_154_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_154_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_155.andOp_155_in0
	// controller for andOp_155.andOp_155_in1
	// Insensitive connections
	always @(*) begin
		andOp_155_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_155_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_156.andOp_156_in0
	// controller for andOp_156.andOp_156_in1
	// Insensitive connections
	always @(*) begin
		andOp_156_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_156_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_157.andOp_157_in0
	// controller for andOp_157.andOp_157_in1
	// Insensitive connections
	always @(*) begin
		andOp_157_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_157_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_158.andOp_158_in0
	// controller for andOp_158.andOp_158_in1
	// Insensitive connections
	always @(*) begin
		andOp_158_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_158_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_159.andOp_159_in0
	// controller for andOp_159.andOp_159_in1
	// Insensitive connections
	always @(*) begin
		andOp_159_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_159_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_160.andOp_160_in0
	// controller for andOp_160.andOp_160_in1
	// Insensitive connections
	always @(*) begin
		andOp_160_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
		andOp_160_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_161.andOp_161_in0
	// controller for andOp_161.andOp_161_in1
	// Insensitive connections
	always @(*) begin
		andOp_161_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_161_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_162.andOp_162_in0
	// controller for andOp_162.andOp_162_in1
	// Insensitive connections
	always @(*) begin
		andOp_162_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_162_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_163.andOp_163_in0
	// controller for andOp_163.andOp_163_in1
	// Insensitive connections
	always @(*) begin
		andOp_163_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_163_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_164.andOp_164_in0
	// controller for andOp_164.andOp_164_in1
	// Insensitive connections
	always @(*) begin
		andOp_164_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_164_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_166.andOp_166_in0
	// controller for andOp_166.andOp_166_in1
	// Insensitive connections
	always @(*) begin
		andOp_166_in0 = valid ? notOp_165_out : notOp_165_out;
		andOp_166_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_168.andOp_168_in0
	// controller for andOp_168.andOp_168_in1
	// Insensitive connections
	always @(*) begin
		andOp_168_in0 = valid ? notOp_167_out : notOp_167_out;
		andOp_168_in1 = valid ? andOp_166_out : andOp_166_out;
	end
	// controller for andOp_170.andOp_170_in0
	// controller for andOp_170.andOp_170_in1
	// Insensitive connections
	always @(*) begin
		andOp_170_in0 = valid ? notOp_169_out : notOp_169_out;
		andOp_170_in1 = valid ? andOp_168_out : andOp_168_out;
	end
	// controller for andOp_172.andOp_172_in0
	// controller for andOp_172.andOp_172_in1
	// Insensitive connections
	always @(*) begin
		andOp_172_in0 = valid ? notOp_171_out : notOp_171_out;
		andOp_172_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_174.andOp_174_in0
	// controller for andOp_174.andOp_174_in1
	// Insensitive connections
	always @(*) begin
		andOp_174_in0 = valid ? notOp_173_out : notOp_173_out;
		andOp_174_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_176.andOp_176_in0
	// controller for andOp_176.andOp_176_in1
	// Insensitive connections
	always @(*) begin
		andOp_176_in0 = valid ? notOp_175_out : notOp_175_out;
		andOp_176_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_178.andOp_178_in0
	// controller for andOp_178.andOp_178_in1
	// Insensitive connections
	always @(*) begin
		andOp_178_in0 = valid ? notOp_177_out : notOp_177_out;
		andOp_178_in1 = valid ? andOp_176_out : andOp_176_out;
	end
	// controller for andOp_180.andOp_180_in0
	// controller for andOp_180.andOp_180_in1
	// Insensitive connections
	always @(*) begin
		andOp_180_in0 = valid ? notOp_179_out : notOp_179_out;
		andOp_180_in1 = valid ? andOp_178_out : andOp_178_out;
	end
	// controller for andOp_185.andOp_185_in0
	// controller for andOp_185.andOp_185_in1
	// Insensitive connections
	always @(*) begin
		andOp_185_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_185_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_186.andOp_186_in0
	// controller for andOp_186.andOp_186_in1
	// Insensitive connections
	always @(*) begin
		andOp_186_in0 = valid ? andOp_185_out : andOp_185_out;
		andOp_186_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_191.andOp_191_in0
	// controller for andOp_191.andOp_191_in1
	// Insensitive connections
	always @(*) begin
		andOp_191_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_191_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_192.andOp_192_in0
	// controller for andOp_192.andOp_192_in1
	// Insensitive connections
	always @(*) begin
		andOp_192_in0 = valid ? andOp_191_out : andOp_191_out;
		andOp_192_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_193.andOp_193_in0
	// controller for andOp_193.andOp_193_in1
	// Insensitive connections
	always @(*) begin
		andOp_193_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_193_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_194.andOp_194_in0
	// controller for andOp_194.andOp_194_in1
	// Insensitive connections
	always @(*) begin
		andOp_194_in0 = valid ? andOp_193_out : andOp_193_out;
		andOp_194_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_195.andOp_195_in0
	// controller for andOp_195.andOp_195_in1
	// Insensitive connections
	always @(*) begin
		andOp_195_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_195_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_196.andOp_196_in0
	// controller for andOp_196.andOp_196_in1
	// Insensitive connections
	always @(*) begin
		andOp_196_in0 = valid ? andOp_195_out : andOp_195_out;
		andOp_196_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_32.andOp_32_in0
	// controller for andOp_32.andOp_32_in1
	// Insensitive connections
	always @(*) begin
		andOp_32_in0 = valid ? bb_0_active_in_state_1_out_data : bb_0_active_in_state_1_out_data;
		andOp_32_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_33.andOp_33_in0
	// controller for andOp_33.andOp_33_in1
	// Insensitive connections
	always @(*) begin
		andOp_33_in0 = valid ? andOp_32_out : andOp_32_out;
		andOp_33_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_35.andOp_35_in0
	// controller for andOp_35.andOp_35_in1
	// Insensitive connections
	always @(*) begin
		andOp_35_in0 = valid ? bb_0_active_in_state_1_out_data : bb_0_active_in_state_1_out_data;
		andOp_35_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_36.andOp_36_in0
	// controller for andOp_36.andOp_36_in1
	// Insensitive connections
	always @(*) begin
		andOp_36_in0 = valid ? andOp_35_out : andOp_35_out;
		andOp_36_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_38.andOp_38_in0
	// controller for andOp_38.andOp_38_in1
	// Insensitive connections
	always @(*) begin
		andOp_38_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_38_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_39.andOp_39_in0
	// controller for andOp_39.andOp_39_in1
	// Insensitive connections
	always @(*) begin
		andOp_39_in0 = valid ? andOp_38_out : andOp_38_out;
		andOp_39_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_41.andOp_41_in0
	// controller for andOp_41.andOp_41_in1
	// Insensitive connections
	always @(*) begin
		andOp_41_in0 = valid ? bb_8_active_in_state_1_out_data : bb_8_active_in_state_1_out_data;
		andOp_41_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_42.andOp_42_in0
	// controller for andOp_42.andOp_42_in1
	// Insensitive connections
	always @(*) begin
		andOp_42_in0 = valid ? andOp_41_out : andOp_41_out;
		andOp_42_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_44.andOp_44_in0
	// controller for andOp_44.andOp_44_in1
	// Insensitive connections
	always @(*) begin
		andOp_44_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
		andOp_44_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_45.andOp_45_in0
	// controller for andOp_45.andOp_45_in1
	// Insensitive connections
	always @(*) begin
		andOp_45_in0 = valid ? andOp_44_out : andOp_44_out;
		andOp_45_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_47.andOp_47_in0
	// controller for andOp_47.andOp_47_in1
	// Insensitive connections
	always @(*) begin
		andOp_47_in0 = valid ? andOp_45_out : andOp_45_out;
		andOp_47_in1 = valid ? in_read_ready : in_read_ready;
	end
	// controller for andOp_49.andOp_49_in0
	// controller for andOp_49.andOp_49_in1
	// Insensitive connections
	always @(*) begin
		andOp_49_in0 = valid ? andOp_45_out : andOp_45_out;
		andOp_49_in1 = valid ? notOp_48_out : notOp_48_out;
	end
	// controller for andOp_50.andOp_50_in0
	// controller for andOp_50.andOp_50_in1
	// Insensitive connections
	always @(*) begin
		andOp_50_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_50_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_51.andOp_51_in0
	// controller for andOp_51.andOp_51_in1
	// Insensitive connections
	always @(*) begin
		andOp_51_in0 = valid ? andOp_50_out : andOp_50_out;
		andOp_51_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_53.andOp_53_in0
	// controller for andOp_53.andOp_53_in1
	// Insensitive connections
	always @(*) begin
		andOp_53_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_53_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_54.andOp_54_in0
	// controller for andOp_54.andOp_54_in1
	// Insensitive connections
	always @(*) begin
		andOp_54_in0 = valid ? andOp_53_out : andOp_53_out;
		andOp_54_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_56.andOp_56_in0
	// controller for andOp_56.andOp_56_in1
	// Insensitive connections
	always @(*) begin
		andOp_56_in0 = valid ? andOp_54_out : andOp_54_out;
		andOp_56_in1 = valid ? data_in_4_31_out_data : data_in_4_31_out_data;
	end
	// controller for andOp_58.andOp_58_in0
	// controller for andOp_58.andOp_58_in1
	// Insensitive connections
	always @(*) begin
		andOp_58_in0 = valid ? andOp_54_out : andOp_54_out;
		andOp_58_in1 = valid ? notOp_57_out : notOp_57_out;
	end
	// controller for andOp_59.andOp_59_in0
	// controller for andOp_59.andOp_59_in1
	// Insensitive connections
	always @(*) begin
		andOp_59_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_59_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_60.andOp_60_in0
	// controller for andOp_60.andOp_60_in1
	// Insensitive connections
	always @(*) begin
		andOp_60_in0 = valid ? andOp_59_out : andOp_59_out;
		andOp_60_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_62.andOp_62_in0
	// controller for andOp_62.andOp_62_in1
	// Insensitive connections
	always @(*) begin
		andOp_62_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_62_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_63.andOp_63_in0
	// controller for andOp_63.andOp_63_in1
	// Insensitive connections
	always @(*) begin
		andOp_63_in0 = valid ? andOp_62_out : andOp_62_out;
		andOp_63_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_65.andOp_65_in0
	// controller for andOp_65.andOp_65_in1
	// Insensitive connections
	always @(*) begin
		andOp_65_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
		andOp_65_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_66.andOp_66_in0
	// controller for andOp_66.andOp_66_in1
	// Insensitive connections
	always @(*) begin
		andOp_66_in0 = valid ? andOp_65_out : andOp_65_out;
		andOp_66_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_68.andOp_68_in0
	// controller for andOp_68.andOp_68_in1
	// Insensitive connections
	always @(*) begin
		andOp_68_in0 = valid ? andOp_66_out : andOp_66_out;
		andOp_68_in1 = valid ? out_write_ready : out_write_ready;
	end
	// controller for andOp_70.andOp_70_in0
	// controller for andOp_70.andOp_70_in1
	// Insensitive connections
	always @(*) begin
		andOp_70_in0 = valid ? andOp_66_out : andOp_66_out;
		andOp_70_in1 = valid ? notOp_69_out : notOp_69_out;
	end
	// controller for andOp_71.andOp_71_in0
	// controller for andOp_71.andOp_71_in1
	// Insensitive connections
	always @(*) begin
		andOp_71_in0 = valid ? bb_5_active_in_state_4_out_data : bb_5_active_in_state_4_out_data;
		andOp_71_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_72.andOp_72_in0
	// controller for andOp_72.andOp_72_in1
	// Insensitive connections
	always @(*) begin
		andOp_72_in0 = valid ? andOp_71_out : andOp_71_out;
		andOp_72_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_74.andOp_74_in0
	// controller for andOp_74.andOp_74_in1
	// Insensitive connections
	always @(*) begin
		andOp_74_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_74_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_75.andOp_75_in0
	// controller for andOp_75.andOp_75_in1
	// Insensitive connections
	always @(*) begin
		andOp_75_in0 = valid ? andOp_74_out : andOp_74_out;
		andOp_75_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_77.andOp_77_in0
	// controller for andOp_77.andOp_77_in1
	// Insensitive connections
	always @(*) begin
		andOp_77_in0 = valid ? andOp_75_out : andOp_75_out;
		andOp_77_in1 = valid ? data_in_4_31_out_data : data_in_4_31_out_data;
	end
	// controller for andOp_79.andOp_79_in0
	// controller for andOp_79.andOp_79_in1
	// Insensitive connections
	always @(*) begin
		andOp_79_in0 = valid ? andOp_75_out : andOp_75_out;
		andOp_79_in1 = valid ? notOp_78_out : notOp_78_out;
	end
	// controller for andOp_80.andOp_80_in0
	// controller for andOp_80.andOp_80_in1
	// Insensitive connections
	always @(*) begin
		andOp_80_in0 = valid ? bb_1_active_in_state_4_out_data : bb_1_active_in_state_4_out_data;
		andOp_80_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_81.andOp_81_in0
	// controller for andOp_81.andOp_81_in1
	// Insensitive connections
	always @(*) begin
		andOp_81_in0 = valid ? andOp_80_out : andOp_80_out;
		andOp_81_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_83_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_active_in_state_1.bb_0_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_1_in_data = eq_84_out;
		end else begin
			bb_0_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_106_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_1.bb_0_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_107_out) begin 
			bb_0_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_2.bb_10_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_2_in_data = eq_91_out;
		end else begin
			bb_10_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_3.bb_10_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_3_in_data = eq_94_out;
		end else begin
			bb_10_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_2.bb_10_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_117_out) begin 
			bb_10_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_3.bb_10_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_121_out) begin 
			bb_10_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_4.bb_1_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_4_in_data = orOp_105_out;
		end else begin
			bb_1_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_4.bb_1_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_137_out) begin 
			bb_1_predecessor_in_state_4_in_data = 32'd4;
		end else if (eq_135_out) begin 
			bb_1_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_4.bb_2_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_4_in_data = orOp_103_out;
		end else begin
			bb_2_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_4.bb_2_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_134_out) begin 
			bb_2_predecessor_in_state_4_in_data = 32'd7;
		end else if (eq_132_out) begin 
			bb_2_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_1.bb_3_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_1_in_data = orOp_86_out;
		end else begin
			bb_3_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_1.bb_3_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_110_out) begin 
			bb_3_predecessor_in_state_1_in_data = 32'd0;
		end else if (eq_108_out) begin 
			bb_3_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_3.bb_4_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_3_in_data = orOp_93_out;
		end else begin
			bb_4_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_4.bb_4_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_4_in_data = eq_101_out;
		end else begin
			bb_4_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_3.bb_4_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_120_out) begin 
			bb_4_predecessor_in_state_3_in_data = 32'd10;
		end else if (eq_118_out) begin 
			bb_4_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_4.bb_4_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_131_out) begin 
			bb_4_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_5_active_in_state_4.bb_5_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_5_active_in_state_4_in_data = orOp_100_out;
		end else begin
			bb_5_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_5_predecessor_in_state_4.bb_5_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_130_out) begin 
			bb_5_predecessor_in_state_4_in_data = 32'd1;
		end else if (eq_128_out) begin 
			bb_5_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_5_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_6_active_in_state_4.bb_6_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_6_active_in_state_4_in_data = orOp_98_out;
		end else begin
			bb_6_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_6_predecessor_in_state_4.bb_6_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_127_out) begin 
			bb_6_predecessor_in_state_4_in_data = 32'd5;
		end else if (eq_125_out) begin 
			bb_6_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_6_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_7_active_in_state_4.bb_7_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_7_active_in_state_4_in_data = orOp_96_out;
		end else begin
			bb_7_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_7_predecessor_in_state_4.bb_7_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_124_out) begin 
			bb_7_predecessor_in_state_4_in_data = 32'd6;
		end else if (eq_122_out) begin 
			bb_7_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_7_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_8_active_in_state_1.bb_8_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_state_1_in_data = orOp_88_out;
		end else begin
			bb_8_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_8_predecessor_in_state_1.bb_8_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_113_out) begin 
			bb_8_predecessor_in_state_1_in_data = 32'd3;
		end else if (eq_111_out) begin 
			bb_8_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_8_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_9_active_in_state_1.bb_9_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_9_active_in_state_1_in_data = orOp_90_out;
		end else begin
			bb_9_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_9_predecessor_in_state_1.bb_9_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_116_out) begin 
			bb_9_predecessor_in_state_1_in_data = 32'd8;
		end else if (eq_114_out) begin 
			bb_9_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_9_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_33_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_34_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_1.br_0_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_36_out) begin 
			br_0_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_37_out) begin 
			br_0_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_2.br_10_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_51_out) begin 
			br_10_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_52_out) begin 
			br_10_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_3.br_10_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_60_out) begin 
			br_10_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_61_out) begin 
			br_10_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_1_happened_in_state_4.br_1_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_81_out) begin 
			br_1_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_82_out) begin 
			br_1_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_1_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_1.br_3_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_39_out) begin 
			br_3_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_40_out) begin 
			br_3_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_3.br_4_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_54_out) begin 
			br_4_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_55_out) begin 
			br_4_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_4.br_4_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_75_out) begin 
			br_4_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_76_out) begin 
			br_4_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_5_happened_in_state_4.br_5_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_72_out) begin 
			br_5_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_73_out) begin 
			br_5_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_5_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_6_happened_in_state_4.br_6_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_66_out) begin 
			br_6_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_67_out) begin 
			br_6_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_6_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_7_happened_in_state_4.br_7_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_63_out) begin 
			br_7_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_64_out) begin 
			br_7_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_7_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_8_happened_in_state_1.br_8_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_42_out) begin 
			br_8_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_43_out) begin 
			br_8_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_8_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_9_happened_in_state_1.br_9_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_45_out) begin 
			br_9_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_46_out) begin 
			br_9_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_9_happened_in_state_1_in_data = 0;
		end
	end
	// controller for concat_149.concat_149_in0
	// controller for concat_149.concat_149_in1
	// Insensitive connections
	always @(*) begin
		concat_149_in0 = valid ? data_in_1_5_out_data : data_in_1_5_out_data;
		concat_149_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for concat_150.concat_150_in0
	// controller for concat_150.concat_150_in1
	// Insensitive connections
	always @(*) begin
		concat_150_in0 = valid ? 32'd4 : 32'd4;
		concat_150_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for data_in_1_1.data_in_1_1_in_data
	always @(*) begin
		if (eq_182_out) begin 
			data_in_1_1_in_data = 32'd0;
		end else if (eq_183_out) begin 
			data_in_1_1_in_data = data_store_1_0;
		end else if (eq_184_out) begin 
			data_in_1_1_in_data = data_store_4_24;
		end else begin
			data_in_1_1_in_data = 0;
		end
	end
	// controller for data_in_1_3.data_in_1_3_in_data
	always @(*) begin
		if (eq_182_out) begin 
			data_in_1_3_in_data = 32'd0;
		end else if (eq_183_out) begin 
			data_in_1_3_in_data = data_store_1_2;
		end else if (eq_184_out) begin 
			data_in_1_3_in_data = data_store_4_26;
		end else begin
			data_in_1_3_in_data = 0;
		end
	end
	// controller for data_in_1_5.data_in_1_5_in_data
	always @(*) begin
		if (eq_182_out) begin 
			data_in_1_5_in_data = 32'd0;
		end else if (eq_183_out) begin 
			data_in_1_5_in_data = data_store_1_4;
		end else if (eq_184_out) begin 
			data_in_1_5_in_data = data_store_4_28;
		end else begin
			data_in_1_5_in_data = 0;
		end
	end
	// controller for data_in_1_7.data_in_1_7_in_data
	always @(*) begin
		if (eq_182_out) begin 
			data_in_1_7_in_data = 1'd0;
		end else if (eq_183_out) begin 
			data_in_1_7_in_data = data_store_1_6;
		end else if (eq_184_out) begin 
			data_in_1_7_in_data = data_store_4_30;
		end else begin
			data_in_1_7_in_data = 0;
		end
	end
	// controller for data_in_2_11.data_in_2_11_in_data
	always @(*) begin
		if (eq_187_out) begin 
			data_in_2_11_in_data = data_store_1_2;
		end else if (eq_188_out) begin 
			data_in_2_11_in_data = data_store_2_10;
		end else begin
			data_in_2_11_in_data = 0;
		end
	end
	// controller for data_in_2_13.data_in_2_13_in_data
	always @(*) begin
		if (eq_187_out) begin 
			data_in_2_13_in_data = data_store_1_4;
		end else if (eq_188_out) begin 
			data_in_2_13_in_data = data_store_2_12;
		end else begin
			data_in_2_13_in_data = 0;
		end
	end
	// controller for data_in_2_15.data_in_2_15_in_data
	always @(*) begin
		if (eq_187_out) begin 
			data_in_2_15_in_data = data_store_1_6;
		end else if (eq_188_out) begin 
			data_in_2_15_in_data = data_store_2_14;
		end else begin
			data_in_2_15_in_data = 0;
		end
	end
	// controller for data_in_2_9.data_in_2_9_in_data
	always @(*) begin
		if (eq_187_out) begin 
			data_in_2_9_in_data = data_store_1_0;
		end else if (eq_188_out) begin 
			data_in_2_9_in_data = data_store_2_8;
		end else begin
			data_in_2_9_in_data = 0;
		end
	end
	// controller for data_in_3_17.data_in_3_17_in_data
	always @(*) begin
		if (eq_189_out) begin 
			data_in_3_17_in_data = data_store_2_8;
		end else if (eq_190_out) begin 
			data_in_3_17_in_data = data_store_3_16;
		end else begin
			data_in_3_17_in_data = 0;
		end
	end
	// controller for data_in_3_19.data_in_3_19_in_data
	always @(*) begin
		if (eq_189_out) begin 
			data_in_3_19_in_data = data_store_2_10;
		end else if (eq_190_out) begin 
			data_in_3_19_in_data = data_store_3_18;
		end else begin
			data_in_3_19_in_data = 0;
		end
	end
	// controller for data_in_3_21.data_in_3_21_in_data
	always @(*) begin
		if (eq_189_out) begin 
			data_in_3_21_in_data = data_store_2_12;
		end else if (eq_190_out) begin 
			data_in_3_21_in_data = data_store_3_20;
		end else begin
			data_in_3_21_in_data = 0;
		end
	end
	// controller for data_in_3_23.data_in_3_23_in_data
	always @(*) begin
		if (eq_189_out) begin 
			data_in_3_23_in_data = data_store_2_14;
		end else if (eq_190_out) begin 
			data_in_3_23_in_data = data_store_3_22;
		end else begin
			data_in_3_23_in_data = 0;
		end
	end
	// controller for data_in_4_25.data_in_4_25_in_data
	always @(*) begin
		if (eq_197_out) begin 
			data_in_4_25_in_data = data_store_3_16;
		end else if (eq_198_out) begin 
			data_in_4_25_in_data = data_store_4_24;
		end else begin
			data_in_4_25_in_data = 0;
		end
	end
	// controller for data_in_4_27.data_in_4_27_in_data
	always @(*) begin
		if (eq_197_out) begin 
			data_in_4_27_in_data = data_store_3_18;
		end else if (eq_198_out) begin 
			data_in_4_27_in_data = data_store_4_26;
		end else begin
			data_in_4_27_in_data = 0;
		end
	end
	// controller for data_in_4_29.data_in_4_29_in_data
	always @(*) begin
		if (eq_197_out) begin 
			data_in_4_29_in_data = data_store_3_20;
		end else if (eq_198_out) begin 
			data_in_4_29_in_data = data_store_4_28;
		end else begin
			data_in_4_29_in_data = 0;
		end
	end
	// controller for data_in_4_31.data_in_4_31_in_data
	always @(*) begin
		if (eq_197_out) begin 
			data_in_4_31_in_data = data_store_3_22;
		end else if (eq_198_out) begin 
			data_in_4_31_in_data = data_store_4_30;
		end else begin
			data_in_4_31_in_data = 0;
		end
	end
	// controller for eq_101.eq_101_in0
	// controller for eq_101.eq_101_in1
	// Insensitive connections
	always @(*) begin
		eq_101_in0 = valid ? 32'd4 : 32'd4;
		eq_101_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_102.eq_102_in0
	// controller for eq_102.eq_102_in1
	// Insensitive connections
	always @(*) begin
		eq_102_in0 = valid ? 32'd2 : 32'd2;
		eq_102_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_104.eq_104_in0
	// controller for eq_104.eq_104_in1
	// Insensitive connections
	always @(*) begin
		eq_104_in0 = valid ? 32'd1 : 32'd1;
		eq_104_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_106.eq_106_in0
	// controller for eq_106.eq_106_in1
	// Insensitive connections
	always @(*) begin
		eq_106_in0 = valid ? 32'd0 : 32'd0;
		eq_106_in1 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
	end
	// controller for eq_107.eq_107_in0
	// controller for eq_107.eq_107_in1
	// Insensitive connections
	always @(*) begin
		eq_107_in0 = valid ? 32'd0 : 32'd0;
		eq_107_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_108.eq_108_in0
	// controller for eq_108.eq_108_in1
	// Insensitive connections
	always @(*) begin
		eq_108_in0 = valid ? 32'd3 : 32'd3;
		eq_108_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_111.eq_111_in0
	// controller for eq_111.eq_111_in1
	// Insensitive connections
	always @(*) begin
		eq_111_in0 = valid ? 32'd8 : 32'd8;
		eq_111_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_114.eq_114_in0
	// controller for eq_114.eq_114_in1
	// Insensitive connections
	always @(*) begin
		eq_114_in0 = valid ? 32'd9 : 32'd9;
		eq_114_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_117.eq_117_in0
	// controller for eq_117.eq_117_in1
	// Insensitive connections
	always @(*) begin
		eq_117_in0 = valid ? 32'd10 : 32'd10;
		eq_117_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_118.eq_118_in0
	// controller for eq_118.eq_118_in1
	// Insensitive connections
	always @(*) begin
		eq_118_in0 = valid ? 32'd4 : 32'd4;
		eq_118_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_121.eq_121_in0
	// controller for eq_121.eq_121_in1
	// Insensitive connections
	always @(*) begin
		eq_121_in0 = valid ? 32'd10 : 32'd10;
		eq_121_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_122.eq_122_in0
	// controller for eq_122.eq_122_in1
	// Insensitive connections
	always @(*) begin
		eq_122_in0 = valid ? 32'd7 : 32'd7;
		eq_122_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_125.eq_125_in0
	// controller for eq_125.eq_125_in1
	// Insensitive connections
	always @(*) begin
		eq_125_in0 = valid ? 32'd6 : 32'd6;
		eq_125_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_128.eq_128_in0
	// controller for eq_128.eq_128_in1
	// Insensitive connections
	always @(*) begin
		eq_128_in0 = valid ? 32'd5 : 32'd5;
		eq_128_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_131.eq_131_in0
	// controller for eq_131.eq_131_in1
	// Insensitive connections
	always @(*) begin
		eq_131_in0 = valid ? 32'd4 : 32'd4;
		eq_131_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_132.eq_132_in0
	// controller for eq_132.eq_132_in1
	// Insensitive connections
	always @(*) begin
		eq_132_in0 = valid ? 32'd2 : 32'd2;
		eq_132_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_135.eq_135_in0
	// controller for eq_135.eq_135_in1
	// Insensitive connections
	always @(*) begin
		eq_135_in0 = valid ? 32'd1 : 32'd1;
		eq_135_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_153.eq_153_in0
	// controller for eq_153.eq_153_in1
	// Insensitive connections
	always @(*) begin
		eq_153_in0 = valid ? 32'd10 : 32'd10;
		eq_153_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_181.eq_181_in0
	// controller for eq_181.eq_181_in1
	// Insensitive connections
	always @(*) begin
		eq_181_in0 = valid ? 32'd0 : 32'd0;
		eq_181_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_182.eq_182_in0
	// controller for eq_182.eq_182_in1
	// Insensitive connections
	always @(*) begin
		eq_182_in0 = valid ? 32'd0 : 32'd0;
		eq_182_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_183.eq_183_in0
	// controller for eq_183.eq_183_in1
	// Insensitive connections
	always @(*) begin
		eq_183_in0 = valid ? 32'd1 : 32'd1;
		eq_183_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_184.eq_184_in0
	// controller for eq_184.eq_184_in1
	// Insensitive connections
	always @(*) begin
		eq_184_in0 = valid ? 32'd4 : 32'd4;
		eq_184_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_187.eq_187_in0
	// controller for eq_187.eq_187_in1
	// Insensitive connections
	always @(*) begin
		eq_187_in0 = valid ? 32'd1 : 32'd1;
		eq_187_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_188.eq_188_in0
	// controller for eq_188.eq_188_in1
	// Insensitive connections
	always @(*) begin
		eq_188_in0 = valid ? 32'd2 : 32'd2;
		eq_188_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_189.eq_189_in0
	// controller for eq_189.eq_189_in1
	// Insensitive connections
	always @(*) begin
		eq_189_in0 = valid ? 32'd2 : 32'd2;
		eq_189_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_190.eq_190_in0
	// controller for eq_190.eq_190_in1
	// Insensitive connections
	always @(*) begin
		eq_190_in0 = valid ? 32'd3 : 32'd3;
		eq_190_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_197.eq_197_in0
	// controller for eq_197.eq_197_in1
	// Insensitive connections
	always @(*) begin
		eq_197_in0 = valid ? 32'd3 : 32'd3;
		eq_197_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_198.eq_198_in0
	// controller for eq_198.eq_198_in1
	// Insensitive connections
	always @(*) begin
		eq_198_in0 = valid ? 32'd4 : 32'd4;
		eq_198_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_83.eq_83_in0
	// controller for eq_83.eq_83_in1
	// Insensitive connections
	always @(*) begin
		eq_83_in0 = valid ? 32'd0 : 32'd0;
		eq_83_in1 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
	end
	// controller for eq_84.eq_84_in0
	// controller for eq_84.eq_84_in1
	// Insensitive connections
	always @(*) begin
		eq_84_in0 = valid ? 32'd0 : 32'd0;
		eq_84_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_85.eq_85_in0
	// controller for eq_85.eq_85_in1
	// Insensitive connections
	always @(*) begin
		eq_85_in0 = valid ? 32'd3 : 32'd3;
		eq_85_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_87.eq_87_in0
	// controller for eq_87.eq_87_in1
	// Insensitive connections
	always @(*) begin
		eq_87_in0 = valid ? 32'd8 : 32'd8;
		eq_87_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_89.eq_89_in0
	// controller for eq_89.eq_89_in1
	// Insensitive connections
	always @(*) begin
		eq_89_in0 = valid ? 32'd9 : 32'd9;
		eq_89_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_91.eq_91_in0
	// controller for eq_91.eq_91_in1
	// Insensitive connections
	always @(*) begin
		eq_91_in0 = valid ? 32'd10 : 32'd10;
		eq_91_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_92.eq_92_in0
	// controller for eq_92.eq_92_in1
	// Insensitive connections
	always @(*) begin
		eq_92_in0 = valid ? 32'd4 : 32'd4;
		eq_92_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_94.eq_94_in0
	// controller for eq_94.eq_94_in1
	// Insensitive connections
	always @(*) begin
		eq_94_in0 = valid ? 32'd10 : 32'd10;
		eq_94_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_95.eq_95_in0
	// controller for eq_95.eq_95_in1
	// Insensitive connections
	always @(*) begin
		eq_95_in0 = valid ? 32'd7 : 32'd7;
		eq_95_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_97.eq_97_in0
	// controller for eq_97.eq_97_in1
	// Insensitive connections
	always @(*) begin
		eq_97_in0 = valid ? 32'd6 : 32'd6;
		eq_97_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_99.eq_99_in0
	// controller for eq_99.eq_99_in1
	// Insensitive connections
	always @(*) begin
		eq_99_in0 = valid ? 32'd5 : 32'd5;
		eq_99_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for icmp_17.cmp_in0_icmp_17
	// controller for icmp_17.cmp_in1_icmp_17
	// Insensitive connections
	always @(*) begin
		cmp_in0_icmp_17 = valid ? add_out_add_16 : add_out_add_16;
		cmp_in1_icmp_17 = valid ? 32'd4 : 32'd4;
	end
	// controller for in.in_read_valid_reg
	always @(*) begin
		if (andOp_146_out) begin 
			in_read_valid_reg = -(1'd1);
		end else begin
			in_read_valid_reg = 0;
		end
	end
	// controller for notOp_109.notOp_109_in0
	// Insensitive connections
	always @(*) begin
		notOp_109_in0 = valid ? eq_108_out : eq_108_out;
	end
	// controller for notOp_112.notOp_112_in0
	// Insensitive connections
	always @(*) begin
		notOp_112_in0 = valid ? eq_111_out : eq_111_out;
	end
	// controller for notOp_115.notOp_115_in0
	// Insensitive connections
	always @(*) begin
		notOp_115_in0 = valid ? eq_114_out : eq_114_out;
	end
	// controller for notOp_119.notOp_119_in0
	// Insensitive connections
	always @(*) begin
		notOp_119_in0 = valid ? eq_118_out : eq_118_out;
	end
	// controller for notOp_123.notOp_123_in0
	// Insensitive connections
	always @(*) begin
		notOp_123_in0 = valid ? eq_122_out : eq_122_out;
	end
	// controller for notOp_126.notOp_126_in0
	// Insensitive connections
	always @(*) begin
		notOp_126_in0 = valid ? eq_125_out : eq_125_out;
	end
	// controller for notOp_129.notOp_129_in0
	// Insensitive connections
	always @(*) begin
		notOp_129_in0 = valid ? eq_128_out : eq_128_out;
	end
	// controller for notOp_133.notOp_133_in0
	// Insensitive connections
	always @(*) begin
		notOp_133_in0 = valid ? eq_132_out : eq_132_out;
	end
	// controller for notOp_136.notOp_136_in0
	// Insensitive connections
	always @(*) begin
		notOp_136_in0 = valid ? eq_135_out : eq_135_out;
	end
	// controller for notOp_165.notOp_165_in0
	// Insensitive connections
	always @(*) begin
		notOp_165_in0 = valid ? andOp_161_out : andOp_161_out;
	end
	// controller for notOp_167.notOp_167_in0
	// Insensitive connections
	always @(*) begin
		notOp_167_in0 = valid ? andOp_49_out : andOp_49_out;
	end
	// controller for notOp_169.notOp_169_in0
	// Insensitive connections
	always @(*) begin
		notOp_169_in0 = valid ? andOp_58_out : andOp_58_out;
	end
	// controller for notOp_171.notOp_171_in0
	// Insensitive connections
	always @(*) begin
		notOp_171_in0 = valid ? andOp_47_out : andOp_47_out;
	end
	// controller for notOp_173.notOp_173_in0
	// Insensitive connections
	always @(*) begin
		notOp_173_in0 = valid ? andOp_162_out : andOp_162_out;
	end
	// controller for notOp_175.notOp_175_in0
	// Insensitive connections
	always @(*) begin
		notOp_175_in0 = valid ? andOp_163_out : andOp_163_out;
	end
	// controller for notOp_177.notOp_177_in0
	// Insensitive connections
	always @(*) begin
		notOp_177_in0 = valid ? andOp_164_out : andOp_164_out;
	end
	// controller for notOp_179.notOp_179_in0
	// Insensitive connections
	always @(*) begin
		notOp_179_in0 = valid ? andOp_70_out : andOp_70_out;
	end
	// controller for notOp_34.notOp_34_in0
	// Insensitive connections
	always @(*) begin
		notOp_34_in0 = valid ? andOp_33_out : andOp_33_out;
	end
	// controller for notOp_37.notOp_37_in0
	// Insensitive connections
	always @(*) begin
		notOp_37_in0 = valid ? andOp_36_out : andOp_36_out;
	end
	// controller for notOp_40.notOp_40_in0
	// Insensitive connections
	always @(*) begin
		notOp_40_in0 = valid ? andOp_39_out : andOp_39_out;
	end
	// controller for notOp_43.notOp_43_in0
	// Insensitive connections
	always @(*) begin
		notOp_43_in0 = valid ? andOp_42_out : andOp_42_out;
	end
	// controller for notOp_46.notOp_46_in0
	// Insensitive connections
	always @(*) begin
		notOp_46_in0 = valid ? andOp_45_out : andOp_45_out;
	end
	// controller for notOp_48.notOp_48_in0
	// Insensitive connections
	always @(*) begin
		notOp_48_in0 = valid ? in_read_ready : in_read_ready;
	end
	// controller for notOp_52.notOp_52_in0
	// Insensitive connections
	always @(*) begin
		notOp_52_in0 = valid ? andOp_51_out : andOp_51_out;
	end
	// controller for notOp_55.notOp_55_in0
	// Insensitive connections
	always @(*) begin
		notOp_55_in0 = valid ? andOp_54_out : andOp_54_out;
	end
	// controller for notOp_57.notOp_57_in0
	// Insensitive connections
	always @(*) begin
		notOp_57_in0 = valid ? data_in_4_31_out_data : data_in_4_31_out_data;
	end
	// controller for notOp_61.notOp_61_in0
	// Insensitive connections
	always @(*) begin
		notOp_61_in0 = valid ? andOp_60_out : andOp_60_out;
	end
	// controller for notOp_64.notOp_64_in0
	// Insensitive connections
	always @(*) begin
		notOp_64_in0 = valid ? andOp_63_out : andOp_63_out;
	end
	// controller for notOp_67.notOp_67_in0
	// Insensitive connections
	always @(*) begin
		notOp_67_in0 = valid ? andOp_66_out : andOp_66_out;
	end
	// controller for notOp_69.notOp_69_in0
	// Insensitive connections
	always @(*) begin
		notOp_69_in0 = valid ? out_write_ready : out_write_ready;
	end
	// controller for notOp_73.notOp_73_in0
	// Insensitive connections
	always @(*) begin
		notOp_73_in0 = valid ? andOp_72_out : andOp_72_out;
	end
	// controller for notOp_76.notOp_76_in0
	// Insensitive connections
	always @(*) begin
		notOp_76_in0 = valid ? andOp_75_out : andOp_75_out;
	end
	// controller for notOp_78.notOp_78_in0
	// Insensitive connections
	always @(*) begin
		notOp_78_in0 = valid ? data_in_4_31_out_data : data_in_4_31_out_data;
	end
	// controller for notOp_82.notOp_82_in0
	// Insensitive connections
	always @(*) begin
		notOp_82_in0 = valid ? andOp_81_out : andOp_81_out;
	end
	// controller for orOp_100.orOp_100_in0
	// controller for orOp_100.orOp_100_in1
	// Insensitive connections
	always @(*) begin
		orOp_100_in0 = valid ? eq_99_out : eq_99_out;
		orOp_100_in1 = valid ? andOp_81_out : andOp_81_out;
	end
	// controller for orOp_103.orOp_103_in0
	// controller for orOp_103.orOp_103_in1
	// Insensitive connections
	always @(*) begin
		orOp_103_in0 = valid ? eq_102_out : eq_102_out;
		orOp_103_in1 = valid ? andOp_63_out : andOp_63_out;
	end
	// controller for orOp_105.orOp_105_in0
	// controller for orOp_105.orOp_105_in1
	// Insensitive connections
	always @(*) begin
		orOp_105_in0 = valid ? eq_104_out : eq_104_out;
		orOp_105_in1 = valid ? andOp_56_out : andOp_56_out;
	end
	// controller for orOp_86.orOp_86_in0
	// controller for orOp_86.orOp_86_in1
	// Insensitive connections
	always @(*) begin
		orOp_86_in0 = valid ? eq_85_out : eq_85_out;
		orOp_86_in1 = valid ? andOp_33_out : andOp_33_out;
	end
	// controller for orOp_88.orOp_88_in0
	// controller for orOp_88.orOp_88_in1
	// Insensitive connections
	always @(*) begin
		orOp_88_in0 = valid ? eq_87_out : eq_87_out;
		orOp_88_in1 = valid ? andOp_39_out : andOp_39_out;
	end
	// controller for orOp_90.orOp_90_in0
	// controller for orOp_90.orOp_90_in1
	// Insensitive connections
	always @(*) begin
		orOp_90_in0 = valid ? eq_89_out : eq_89_out;
		orOp_90_in1 = valid ? andOp_42_out : andOp_42_out;
	end
	// controller for orOp_93.orOp_93_in0
	// controller for orOp_93.orOp_93_in1
	// Insensitive connections
	always @(*) begin
		orOp_93_in0 = valid ? eq_92_out : eq_92_out;
		orOp_93_in1 = valid ? andOp_51_out : andOp_51_out;
	end
	// controller for orOp_96.orOp_96_in0
	// controller for orOp_96.orOp_96_in1
	// Insensitive connections
	always @(*) begin
		orOp_96_in0 = valid ? eq_95_out : eq_95_out;
		orOp_96_in1 = valid ? andOp_68_out : andOp_68_out;
	end
	// controller for orOp_98.orOp_98_in0
	// controller for orOp_98.orOp_98_in1
	// Insensitive connections
	always @(*) begin
		orOp_98_in0 = valid ? eq_97_out : eq_97_out;
		orOp_98_in1 = valid ? andOp_72_out : andOp_72_out;
	end
	// controller for out.out_in_data_reg
	always @(*) begin
		if (andOp_158_out) begin 
			out_in_data_reg = rdata_ram_0;
		end else begin
			out_in_data_reg = 0;
		end
	end
	// controller for out.out_write_valid_reg
	always @(*) begin
		if (andOp_159_out) begin 
			out_write_valid_reg = -(1'd1);
		end else begin
			out_write_valid_reg = 0;
		end
	end
	// controller for phi_7.phi_in_phi_7
	// controller for phi_7.phi_last_block_phi_7
	// controller for phi_7.phi_s_phi_7
	// Insensitive connections
	always @(*) begin
		phi_in_phi_7 = valid ? concat_149_out : concat_149_out;
		phi_last_block_phi_7 = valid ? bb_3_predecessor_in_state_1_out_data : bb_3_predecessor_in_state_1_out_data;
		phi_s_phi_7 = valid ? concat_150_out : concat_150_out;
	end
	// controller for ram_0.raddr_ram_0_reg
	always @(*) begin
		if (andOp_142_out) begin 
			raddr_ram_0_reg = 32'd0;
		end else if (andOp_144_out) begin 
			raddr_ram_0_reg = 32'd0;
		end else begin
			raddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.waddr_ram_0_reg
	always @(*) begin
		if (andOp_141_out) begin 
			waddr_ram_0_reg = 32'd0;
		end else if (andOp_143_out) begin 
			waddr_ram_0_reg = 32'd0;
		end else begin
			waddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wdata_ram_0_reg
	always @(*) begin
		if (andOp_141_out) begin 
			wdata_ram_0_reg = 32'd0;
		end else if (andOp_143_out) begin 
			wdata_ram_0_reg = add_out_add_14;
		end else begin
			wdata_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wen_ram_0_reg
	always @(*) begin
		if (andOp_141_out) begin 
			wen_ram_0_reg = 1'd1;
		end else if (andOp_143_out) begin 
			wen_ram_0_reg = 1'd1;
		end else begin
			wen_ram_0_reg = 0;
		end
	end
	// controller for ret_22.valid_reg
	always @(*) begin
		if (andOp_157_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// controller for tmp_output_152.tmp_output_152_in_data
	always @(*) begin
		if (eq_153_out) begin 
			tmp_output_152_in_data = in_out_data;
		end else begin
			tmp_output_152_in_data = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			data_store_1_0 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_0 <= data_in_1_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_2 <= 0;
		end else begin
			if (andOp_186_out) begin
				data_store_1_2 <= phi_out_phi_7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_4 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_4 <= data_in_1_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_6 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_6 <= data_in_1_7_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_10 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_10 <= data_in_2_11_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_12 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_12 <= data_in_2_13_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_14 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_14 <= data_in_2_15_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_8 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_8 <= data_in_2_9_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_16 <= 0;
		end else begin
			if (andOp_192_out) begin
				data_store_3_16 <= in_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_18 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_18 <= data_in_3_19_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_20 <= 0;
		end else begin
			if (andOp_194_out) begin
				data_store_3_20 <= add_out_add_16;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_22 <= 0;
		end else begin
			if (andOp_196_out) begin
				data_store_3_22 <= cmp_out_icmp_17;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_24 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_24 <= data_in_4_25_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_26 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_26 <= data_in_4_27_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_28 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_28 <= data_in_4_29_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_30 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_30 <= data_in_4_31_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_161_out) begin
				global_state <= 32'd1;
			end
			if (andOp_162_out) begin
				global_state <= 32'd3;
			end
			if (andOp_163_out) begin
				global_state <= 32'd4;
			end
			if (andOp_164_out) begin
				global_state <= 32'd4;
			end
			if (andOp_47_out) begin
				global_state <= 32'd2;
			end
			if (andOp_49_out) begin
				global_state <= 32'd1;
			end
			if (andOp_58_out) begin
				global_state <= 32'd1;
			end
			if (andOp_70_out) begin
				global_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (1'd1) begin
				state_0_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_161_out) begin
				state_1_entry_BB_reg <= 32'd0;
			end
			if (andOp_49_out) begin
				state_1_entry_BB_reg <= 32'd9;
			end
			if (andOp_58_out) begin
				state_1_entry_BB_reg <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_161_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_170_out) begin
				state_1_is_active <= 1'd0;
			end
			if (andOp_49_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_58_out) begin
				state_1_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_161_out) begin
				state_1_last_BB_reg <= bb_0_predecessor_in_state_0_out_data;
			end
			if (andOp_49_out) begin
				state_1_last_BB_reg <= 32'd9;
			end
			if (andOp_58_out) begin
				state_1_last_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_161_out) begin
				state_1_last_state <= 32'd0;
			end
			if (andOp_49_out) begin
				state_1_last_state <= 32'd1;
			end
			if (andOp_58_out) begin
				state_1_last_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_47_out) begin
				state_2_entry_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_172_out) begin
				state_2_is_active <= 1'd0;
			end
			if (andOp_47_out) begin
				state_2_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_47_out) begin
				state_2_last_BB_reg <= 32'd9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_47_out) begin
				state_2_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_162_out) begin
				state_3_entry_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_162_out) begin
				state_3_is_active <= 1'd1;
			end
			if (andOp_174_out) begin
				state_3_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_162_out) begin
				state_3_last_BB_reg <= bb_10_predecessor_in_state_2_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_state <= 0;
		end else begin
			if (andOp_162_out) begin
				state_3_last_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_163_out) begin
				state_4_entry_BB_reg <= 32'd4;
			end
			if (andOp_164_out) begin
				state_4_entry_BB_reg <= 32'd2;
			end
			if (andOp_70_out) begin
				state_4_entry_BB_reg <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_163_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_164_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_180_out) begin
				state_4_is_active <= 1'd0;
			end
			if (andOp_70_out) begin
				state_4_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_163_out) begin
				state_4_last_BB_reg <= bb_4_predecessor_in_state_3_out_data;
			end
			if (andOp_164_out) begin
				state_4_last_BB_reg <= bb_2_predecessor_in_state_4_out_data;
			end
			if (andOp_70_out) begin
				state_4_last_BB_reg <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_state <= 0;
		end else begin
			if (andOp_163_out) begin
				state_4_last_state <= 32'd3;
			end
			if (andOp_164_out) begin
				state_4_last_state <= 32'd4;
			end
			if (andOp_70_out) begin
				state_4_last_state <= 32'd4;
			end
		end
	end

endmodule

