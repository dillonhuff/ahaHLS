module vadd_smul_fifo(input [0:0] clk, input [0:0] rst, output [0:0] valid, output [31:0] arg_0_in_data, input [31:0] arg_0_out_data, input [0:0] arg_0_read_ready, output [0:0] arg_0_read_valid, input [0:0] arg_0_write_ready, output [0:0] arg_0_write_valid, output [31:0] arg_1_in_data, input [31:0] arg_1_out_data, input [0:0] arg_1_read_ready, output [0:0] arg_1_read_valid, input [0:0] arg_1_write_ready, output [0:0] arg_1_write_valid, output [31:0] arg_2_in_data, input [31:0] arg_2_out_data, input [0:0] arg_2_read_ready, output [0:0] arg_2_read_valid, input [0:0] arg_2_write_ready, output [0:0] arg_2_write_valid);

	reg [0:0] valid_reg;
	reg [31:0] arg_0_in_data_reg;
	reg [0:0] arg_0_read_valid_reg;
	reg [0:0] arg_0_write_valid_reg;
	reg [31:0] arg_1_in_data_reg;
	reg [0:0] arg_1_read_valid_reg;
	reg [0:0] arg_1_write_valid_reg;
	reg [31:0] arg_2_in_data_reg;
	reg [0:0] arg_2_read_valid_reg;
	reg [0:0] arg_2_write_valid_reg;

	assign valid = valid_reg;
	assign arg_0_in_data = arg_0_in_data_reg;
	assign arg_0_read_valid = arg_0_read_valid_reg;
	assign arg_0_write_valid = arg_0_write_valid_reg;
	assign arg_1_in_data = arg_1_in_data_reg;
	assign arg_1_read_valid = arg_1_read_valid_reg;
	assign arg_1_write_valid = arg_1_write_valid_reg;
	assign arg_2_in_data = arg_2_in_data_reg;
	assign arg_2_read_valid = arg_2_read_valid_reg;
	assign arg_2_write_valid = arg_2_write_valid_reg;

	// Start debug wires and ports

	initial begin
	end






	// End debug wires and ports

	// Start Functional Units
	br_dummy br_unit();

	wire [31:0] icmp_icmp16_in0;
	wire [31:0] icmp_icmp16_in1;
	wire [0:0] icmp_icmp16_out;
	ne #(.WIDTH(32)) icmp_icmp16(.in0(icmp_icmp16_in0), .in1(icmp_icmp16_in1), .out(icmp_icmp16_out));

	wire [63:0] phi_phi28_in;
	wire [31:0] phi_phi28_last_block;
	wire [63:0] phi_phi28_s;
	wire [31:0] phi_phi28_out;
	phi #(.DEBUG_ID(1), .NB_PAIR(2), .WIDTH(32)) phi_phi28(.in(phi_phi28_in), .last_block(phi_phi28_last_block), .out(phi_phi28_out), .s(phi_phi28_s));

	reg [31:0] _____dlr_0___eq___alloca___dlr_builtin_fifo_32_in_data;
	reg [0:0] _____dlr_0___eq___alloca___dlr_builtin_fifo_32_read_valid;
	reg [0:0] _____dlr_0___eq___alloca___dlr_builtin_fifo_32_write_valid;
	wire [31:0] _____dlr_0___eq___alloca___dlr_builtin_fifo_32_out_data;
	wire [0:0] _____dlr_0___eq___alloca___dlr_builtin_fifo_32_read_ready;
	wire [0:0] _____dlr_0___eq___alloca___dlr_builtin_fifo_32_write_ready;
	fifo #(.DEPTH(16), .WIDTH(32)) _____dlr_0___eq___alloca___dlr_builtin_fifo_32(.clk(clk), .in_data(_____dlr_0___eq___alloca___dlr_builtin_fifo_32_in_data), .out_data(_____dlr_0___eq___alloca___dlr_builtin_fifo_32_out_data), .read_ready(_____dlr_0___eq___alloca___dlr_builtin_fifo_32_read_ready), .read_valid(_____dlr_0___eq___alloca___dlr_builtin_fifo_32_read_valid), .rst(rst), .write_ready(_____dlr_0___eq___alloca___dlr_builtin_fifo_32_write_ready), .write_valid(_____dlr_0___eq___alloca___dlr_builtin_fifo_32_write_valid));

	wire [63:0] phi_phi3_in;
	wire [31:0] phi_phi3_last_block;
	wire [63:0] phi_phi3_s;
	wire [31:0] phi_phi3_out;
	phi #(.DEBUG_ID(2), .NB_PAIR(2), .WIDTH(32)) phi_phi3(.in(phi_phi3_in), .last_block(phi_phi3_last_block), .out(phi_phi3_out), .s(phi_phi3_s));

	wire [31:0] icmp_icmp37_in0;
	wire [31:0] icmp_icmp37_in1;
	wire [0:0] icmp_icmp37_out;
	ne #(.WIDTH(32)) icmp_icmp37(.in0(icmp_icmp37_in0), .in1(icmp_icmp37_in1), .out(icmp_icmp37_out));

	wire [31:0] mul_mul39_in0;
	wire [31:0] mul_mul39_in1;
	wire [31:0] mul_mul39_out;
	mul #(.WIDTH(32)) mul_mul39(.in0(mul_mul39_in0), .in1(mul_mul39_in1), .out(mul_mul39_out));

	wire [31:0] add_add5_in0;
	wire [31:0] add_add5_in1;
	wire [31:0] add_add5_out;
	add #(.WIDTH(32)) add_add5(.in0(add_add5_in0), .in1(add_add5_in1), .out(add_add5_out));

	wire [31:0] add_add26_in0;
	wire [31:0] add_add26_in1;
	wire [31:0] add_add26_out;
	add #(.WIDTH(32)) add_add26(.in0(add_add26_in0), .in1(add_add26_in1), .out(add_add26_out));

	wire [31:0] add_add29_in0;
	wire [31:0] add_add29_in1;
	wire [31:0] add_add29_out;
	add #(.WIDTH(32)) add_add29(.in0(add_add29_in0), .in1(add_add29_in1), .out(add_add29_out));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] bb_15_active_in_state_1_in_data;
	wire [0:0] bb_15_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_15_active_in_state_1(.in_data(bb_15_active_in_state_1_in_data), .out_data(bb_15_active_in_state_1_out_data));

	reg [31:0] bb_15_predecessor_in_state_1_in_data;
	wire [31:0] bb_15_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_15_predecessor_in_state_1(.in_data(bb_15_predecessor_in_state_1_in_data), .out_data(bb_15_predecessor_in_state_1_out_data));

	reg [0:0] br_15_happened_in_state_1_in_data;
	wire [0:0] br_15_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_15_happened_in_state_1(.in_data(br_15_happened_in_state_1_in_data), .out_data(br_15_happened_in_state_1_out_data));

	reg [0:0] bb_4_active_in_state_1_in_data;
	wire [0:0] bb_4_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_1(.in_data(bb_4_active_in_state_1_in_data), .out_data(bb_4_active_in_state_1_out_data));

	reg [31:0] bb_4_predecessor_in_state_1_in_data;
	wire [31:0] bb_4_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_1(.in_data(bb_4_predecessor_in_state_1_in_data), .out_data(bb_4_predecessor_in_state_1_out_data));

	reg [0:0] br_4_happened_in_state_1_in_data;
	wire [0:0] br_4_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_1(.in_data(br_4_happened_in_state_1_in_data), .out_data(br_4_happened_in_state_1_out_data));

	reg [0:0] bb_16_active_in_state_1_in_data;
	wire [0:0] bb_16_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_16_active_in_state_1(.in_data(bb_16_active_in_state_1_in_data), .out_data(bb_16_active_in_state_1_out_data));

	reg [31:0] bb_16_predecessor_in_state_1_in_data;
	wire [31:0] bb_16_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_16_predecessor_in_state_1(.in_data(bb_16_predecessor_in_state_1_in_data), .out_data(bb_16_predecessor_in_state_1_out_data));

	reg [0:0] br_16_happened_in_state_1_in_data;
	wire [0:0] br_16_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_16_happened_in_state_1(.in_data(br_16_happened_in_state_1_in_data), .out_data(br_16_happened_in_state_1_out_data));

	reg [0:0] bb_17_active_in_state_2_in_data;
	wire [0:0] bb_17_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_17_active_in_state_2(.in_data(bb_17_active_in_state_2_in_data), .out_data(bb_17_active_in_state_2_out_data));

	reg [31:0] bb_17_predecessor_in_state_2_in_data;
	wire [31:0] bb_17_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_17_predecessor_in_state_2(.in_data(bb_17_predecessor_in_state_2_in_data), .out_data(bb_17_predecessor_in_state_2_out_data));

	reg [0:0] br_17_happened_in_state_2_in_data;
	wire [0:0] br_17_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_17_happened_in_state_2(.in_data(br_17_happened_in_state_2_in_data), .out_data(br_17_happened_in_state_2_out_data));

	reg [0:0] bb_17_active_in_state_3_in_data;
	wire [0:0] bb_17_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_17_active_in_state_3(.in_data(bb_17_active_in_state_3_in_data), .out_data(bb_17_active_in_state_3_out_data));

	reg [31:0] bb_17_predecessor_in_state_3_in_data;
	wire [31:0] bb_17_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_17_predecessor_in_state_3(.in_data(bb_17_predecessor_in_state_3_in_data), .out_data(bb_17_predecessor_in_state_3_out_data));

	reg [0:0] br_17_happened_in_state_3_in_data;
	wire [0:0] br_17_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_17_happened_in_state_3(.in_data(br_17_happened_in_state_3_in_data), .out_data(br_17_happened_in_state_3_out_data));

	reg [0:0] bb_18_active_in_state_3_in_data;
	wire [0:0] bb_18_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_18_active_in_state_3(.in_data(bb_18_active_in_state_3_in_data), .out_data(bb_18_active_in_state_3_out_data));

	reg [31:0] bb_18_predecessor_in_state_3_in_data;
	wire [31:0] bb_18_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_18_predecessor_in_state_3(.in_data(bb_18_predecessor_in_state_3_in_data), .out_data(bb_18_predecessor_in_state_3_out_data));

	reg [0:0] br_18_happened_in_state_3_in_data;
	wire [0:0] br_18_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_18_happened_in_state_3(.in_data(br_18_happened_in_state_3_in_data), .out_data(br_18_happened_in_state_3_out_data));

	reg [0:0] bb_19_active_in_state_3_in_data;
	wire [0:0] bb_19_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_19_active_in_state_3(.in_data(bb_19_active_in_state_3_in_data), .out_data(bb_19_active_in_state_3_out_data));

	reg [31:0] bb_19_predecessor_in_state_3_in_data;
	wire [31:0] bb_19_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_19_predecessor_in_state_3(.in_data(bb_19_predecessor_in_state_3_in_data), .out_data(bb_19_predecessor_in_state_3_out_data));

	reg [0:0] br_19_happened_in_state_3_in_data;
	wire [0:0] br_19_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_19_happened_in_state_3(.in_data(br_19_happened_in_state_3_in_data), .out_data(br_19_happened_in_state_3_out_data));

	reg [0:0] bb_5_active_in_state_3_in_data;
	wire [0:0] bb_5_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_5_active_in_state_3(.in_data(bb_5_active_in_state_3_in_data), .out_data(bb_5_active_in_state_3_out_data));

	reg [31:0] bb_5_predecessor_in_state_3_in_data;
	wire [31:0] bb_5_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_5_predecessor_in_state_3(.in_data(bb_5_predecessor_in_state_3_in_data), .out_data(bb_5_predecessor_in_state_3_out_data));

	reg [0:0] br_5_happened_in_state_3_in_data;
	wire [0:0] br_5_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_5_happened_in_state_3(.in_data(br_5_happened_in_state_3_in_data), .out_data(br_5_happened_in_state_3_out_data));

	reg [0:0] bb_20_active_in_state_4_in_data;
	wire [0:0] bb_20_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_20_active_in_state_4(.in_data(bb_20_active_in_state_4_in_data), .out_data(bb_20_active_in_state_4_out_data));

	reg [31:0] bb_20_predecessor_in_state_4_in_data;
	wire [31:0] bb_20_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_20_predecessor_in_state_4(.in_data(bb_20_predecessor_in_state_4_in_data), .out_data(bb_20_predecessor_in_state_4_out_data));

	reg [0:0] br_20_happened_in_state_4_in_data;
	wire [0:0] br_20_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_20_happened_in_state_4(.in_data(br_20_happened_in_state_4_in_data), .out_data(br_20_happened_in_state_4_out_data));

	reg [0:0] bb_22_active_in_state_5_in_data;
	wire [0:0] bb_22_active_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) bb_22_active_in_state_5(.in_data(bb_22_active_in_state_5_in_data), .out_data(bb_22_active_in_state_5_out_data));

	reg [31:0] bb_22_predecessor_in_state_5_in_data;
	wire [31:0] bb_22_predecessor_in_state_5_out_data;
	hls_wire #(.WIDTH(32)) bb_22_predecessor_in_state_5(.in_data(bb_22_predecessor_in_state_5_in_data), .out_data(bb_22_predecessor_in_state_5_out_data));

	reg [0:0] br_22_happened_in_state_5_in_data;
	wire [0:0] br_22_happened_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) br_22_happened_in_state_5(.in_data(br_22_happened_in_state_5_in_data), .out_data(br_22_happened_in_state_5_out_data));

	reg [0:0] bb_23_active_in_state_5_in_data;
	wire [0:0] bb_23_active_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) bb_23_active_in_state_5(.in_data(bb_23_active_in_state_5_in_data), .out_data(bb_23_active_in_state_5_out_data));

	reg [31:0] bb_23_predecessor_in_state_5_in_data;
	wire [31:0] bb_23_predecessor_in_state_5_out_data;
	hls_wire #(.WIDTH(32)) bb_23_predecessor_in_state_5(.in_data(bb_23_predecessor_in_state_5_in_data), .out_data(bb_23_predecessor_in_state_5_out_data));

	reg [0:0] br_23_happened_in_state_5_in_data;
	wire [0:0] br_23_happened_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) br_23_happened_in_state_5(.in_data(br_23_happened_in_state_5_in_data), .out_data(br_23_happened_in_state_5_out_data));

	reg [0:0] bb_7_active_in_state_5_in_data;
	wire [0:0] bb_7_active_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) bb_7_active_in_state_5(.in_data(bb_7_active_in_state_5_in_data), .out_data(bb_7_active_in_state_5_out_data));

	reg [31:0] bb_7_predecessor_in_state_5_in_data;
	wire [31:0] bb_7_predecessor_in_state_5_out_data;
	hls_wire #(.WIDTH(32)) bb_7_predecessor_in_state_5(.in_data(bb_7_predecessor_in_state_5_in_data), .out_data(bb_7_predecessor_in_state_5_out_data));

	reg [0:0] br_7_happened_in_state_5_in_data;
	wire [0:0] br_7_happened_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) br_7_happened_in_state_5(.in_data(br_7_happened_in_state_5_in_data), .out_data(br_7_happened_in_state_5_out_data));

	reg [0:0] bb_21_active_in_state_5_in_data;
	wire [0:0] bb_21_active_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) bb_21_active_in_state_5(.in_data(bb_21_active_in_state_5_in_data), .out_data(bb_21_active_in_state_5_out_data));

	reg [31:0] bb_21_predecessor_in_state_5_in_data;
	wire [31:0] bb_21_predecessor_in_state_5_out_data;
	hls_wire #(.WIDTH(32)) bb_21_predecessor_in_state_5(.in_data(bb_21_predecessor_in_state_5_in_data), .out_data(bb_21_predecessor_in_state_5_out_data));

	reg [0:0] br_21_happened_in_state_5_in_data;
	wire [0:0] br_21_happened_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) br_21_happened_in_state_5(.in_data(br_21_happened_in_state_5_in_data), .out_data(br_21_happened_in_state_5_out_data));

	reg [0:0] bb_20_active_in_state_5_in_data;
	wire [0:0] bb_20_active_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) bb_20_active_in_state_5(.in_data(bb_20_active_in_state_5_in_data), .out_data(bb_20_active_in_state_5_out_data));

	reg [31:0] bb_20_predecessor_in_state_5_in_data;
	wire [31:0] bb_20_predecessor_in_state_5_out_data;
	hls_wire #(.WIDTH(32)) bb_20_predecessor_in_state_5(.in_data(bb_20_predecessor_in_state_5_in_data), .out_data(bb_20_predecessor_in_state_5_out_data));

	reg [0:0] br_20_happened_in_state_5_in_data;
	wire [0:0] br_20_happened_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) br_20_happened_in_state_5(.in_data(br_20_happened_in_state_5_in_data), .out_data(br_20_happened_in_state_5_out_data));

	reg [0:0] bb_6_active_in_state_5_in_data;
	wire [0:0] bb_6_active_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) bb_6_active_in_state_5(.in_data(bb_6_active_in_state_5_in_data), .out_data(bb_6_active_in_state_5_out_data));

	reg [31:0] bb_6_predecessor_in_state_5_in_data;
	wire [31:0] bb_6_predecessor_in_state_5_out_data;
	hls_wire #(.WIDTH(32)) bb_6_predecessor_in_state_5(.in_data(bb_6_predecessor_in_state_5_in_data), .out_data(bb_6_predecessor_in_state_5_out_data));

	reg [0:0] br_6_happened_in_state_5_in_data;
	wire [0:0] br_6_happened_in_state_5_out_data;
	hls_wire #(.WIDTH(1)) br_6_happened_in_state_5(.in_data(br_6_happened_in_state_5_in_data), .out_data(br_6_happened_in_state_5_out_data));

	reg [0:0] bb_9_active_in_state_6_in_data;
	wire [0:0] bb_9_active_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) bb_9_active_in_state_6(.in_data(bb_9_active_in_state_6_in_data), .out_data(bb_9_active_in_state_6_out_data));

	reg [31:0] bb_9_predecessor_in_state_6_in_data;
	wire [31:0] bb_9_predecessor_in_state_6_out_data;
	hls_wire #(.WIDTH(32)) bb_9_predecessor_in_state_6(.in_data(bb_9_predecessor_in_state_6_in_data), .out_data(bb_9_predecessor_in_state_6_out_data));

	reg [0:0] br_9_happened_in_state_6_in_data;
	wire [0:0] br_9_happened_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) br_9_happened_in_state_6(.in_data(br_9_happened_in_state_6_in_data), .out_data(br_9_happened_in_state_6_out_data));

	reg [0:0] bb_1_active_in_state_6_in_data;
	wire [0:0] bb_1_active_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_6(.in_data(bb_1_active_in_state_6_in_data), .out_data(bb_1_active_in_state_6_out_data));

	reg [31:0] bb_1_predecessor_in_state_6_in_data;
	wire [31:0] bb_1_predecessor_in_state_6_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_6(.in_data(bb_1_predecessor_in_state_6_in_data), .out_data(bb_1_predecessor_in_state_6_out_data));

	reg [0:0] br_1_happened_in_state_6_in_data;
	wire [0:0] br_1_happened_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened_in_state_6(.in_data(br_1_happened_in_state_6_in_data), .out_data(br_1_happened_in_state_6_out_data));

	reg [0:0] bb_10_active_in_state_6_in_data;
	wire [0:0] bb_10_active_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_6(.in_data(bb_10_active_in_state_6_in_data), .out_data(bb_10_active_in_state_6_out_data));

	reg [31:0] bb_10_predecessor_in_state_6_in_data;
	wire [31:0] bb_10_predecessor_in_state_6_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_6(.in_data(bb_10_predecessor_in_state_6_in_data), .out_data(bb_10_predecessor_in_state_6_out_data));

	reg [0:0] br_10_happened_in_state_6_in_data;
	wire [0:0] br_10_happened_in_state_6_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_6(.in_data(br_10_happened_in_state_6_in_data), .out_data(br_10_happened_in_state_6_out_data));

	reg [0:0] bb_11_active_in_state_7_in_data;
	wire [0:0] bb_11_active_in_state_7_out_data;
	hls_wire #(.WIDTH(1)) bb_11_active_in_state_7(.in_data(bb_11_active_in_state_7_in_data), .out_data(bb_11_active_in_state_7_out_data));

	reg [31:0] bb_11_predecessor_in_state_7_in_data;
	wire [31:0] bb_11_predecessor_in_state_7_out_data;
	hls_wire #(.WIDTH(32)) bb_11_predecessor_in_state_7(.in_data(bb_11_predecessor_in_state_7_in_data), .out_data(bb_11_predecessor_in_state_7_out_data));

	reg [0:0] br_11_happened_in_state_7_in_data;
	wire [0:0] br_11_happened_in_state_7_out_data;
	hls_wire #(.WIDTH(1)) br_11_happened_in_state_7(.in_data(br_11_happened_in_state_7_in_data), .out_data(br_11_happened_in_state_7_out_data));

	reg [0:0] bb_13_active_in_state_8_in_data;
	wire [0:0] bb_13_active_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) bb_13_active_in_state_8(.in_data(bb_13_active_in_state_8_in_data), .out_data(bb_13_active_in_state_8_out_data));

	reg [31:0] bb_13_predecessor_in_state_8_in_data;
	wire [31:0] bb_13_predecessor_in_state_8_out_data;
	hls_wire #(.WIDTH(32)) bb_13_predecessor_in_state_8(.in_data(bb_13_predecessor_in_state_8_in_data), .out_data(bb_13_predecessor_in_state_8_out_data));

	reg [0:0] br_13_happened_in_state_8_in_data;
	wire [0:0] br_13_happened_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) br_13_happened_in_state_8(.in_data(br_13_happened_in_state_8_in_data), .out_data(br_13_happened_in_state_8_out_data));

	reg [0:0] bb_14_active_in_state_8_in_data;
	wire [0:0] bb_14_active_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) bb_14_active_in_state_8(.in_data(bb_14_active_in_state_8_in_data), .out_data(bb_14_active_in_state_8_out_data));

	reg [31:0] bb_14_predecessor_in_state_8_in_data;
	wire [31:0] bb_14_predecessor_in_state_8_out_data;
	hls_wire #(.WIDTH(32)) bb_14_predecessor_in_state_8(.in_data(bb_14_predecessor_in_state_8_in_data), .out_data(bb_14_predecessor_in_state_8_out_data));

	reg [0:0] br_14_happened_in_state_8_in_data;
	wire [0:0] br_14_happened_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) br_14_happened_in_state_8(.in_data(br_14_happened_in_state_8_in_data), .out_data(br_14_happened_in_state_8_out_data));

	reg [0:0] bb_2_active_in_state_8_in_data;
	wire [0:0] bb_2_active_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_8(.in_data(bb_2_active_in_state_8_in_data), .out_data(bb_2_active_in_state_8_out_data));

	reg [31:0] bb_2_predecessor_in_state_8_in_data;
	wire [31:0] bb_2_predecessor_in_state_8_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_8(.in_data(bb_2_predecessor_in_state_8_in_data), .out_data(bb_2_predecessor_in_state_8_out_data));

	reg [0:0] br_2_happened_in_state_8_in_data;
	wire [0:0] br_2_happened_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) br_2_happened_in_state_8(.in_data(br_2_happened_in_state_8_in_data), .out_data(br_2_happened_in_state_8_out_data));

	reg [0:0] bb_11_active_in_state_8_in_data;
	wire [0:0] bb_11_active_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) bb_11_active_in_state_8(.in_data(bb_11_active_in_state_8_in_data), .out_data(bb_11_active_in_state_8_out_data));

	reg [31:0] bb_11_predecessor_in_state_8_in_data;
	wire [31:0] bb_11_predecessor_in_state_8_out_data;
	hls_wire #(.WIDTH(32)) bb_11_predecessor_in_state_8(.in_data(bb_11_predecessor_in_state_8_in_data), .out_data(bb_11_predecessor_in_state_8_out_data));

	reg [0:0] br_11_happened_in_state_8_in_data;
	wire [0:0] br_11_happened_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) br_11_happened_in_state_8(.in_data(br_11_happened_in_state_8_in_data), .out_data(br_11_happened_in_state_8_out_data));

	reg [0:0] bb_3_active_in_state_8_in_data;
	wire [0:0] bb_3_active_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_8(.in_data(bb_3_active_in_state_8_in_data), .out_data(bb_3_active_in_state_8_out_data));

	reg [31:0] bb_3_predecessor_in_state_8_in_data;
	wire [31:0] bb_3_predecessor_in_state_8_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_8(.in_data(bb_3_predecessor_in_state_8_in_data), .out_data(bb_3_predecessor_in_state_8_out_data));

	reg [0:0] br_3_happened_in_state_8_in_data;
	wire [0:0] br_3_happened_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_8(.in_data(br_3_happened_in_state_8_in_data), .out_data(br_3_happened_in_state_8_out_data));

	reg [0:0] bb_12_active_in_state_8_in_data;
	wire [0:0] bb_12_active_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) bb_12_active_in_state_8(.in_data(bb_12_active_in_state_8_in_data), .out_data(bb_12_active_in_state_8_out_data));

	reg [31:0] bb_12_predecessor_in_state_8_in_data;
	wire [31:0] bb_12_predecessor_in_state_8_out_data;
	hls_wire #(.WIDTH(32)) bb_12_predecessor_in_state_8(.in_data(bb_12_predecessor_in_state_8_in_data), .out_data(bb_12_predecessor_in_state_8_out_data));

	reg [0:0] br_12_happened_in_state_8_in_data;
	wire [0:0] br_12_happened_in_state_8_out_data;
	hls_wire #(.WIDTH(1)) br_12_happened_in_state_8(.in_data(br_12_happened_in_state_8_in_data), .out_data(br_12_happened_in_state_8_out_data));

	reg [0:0] bb_8_active_in_state_9_in_data;
	wire [0:0] bb_8_active_in_state_9_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active_in_state_9(.in_data(bb_8_active_in_state_9_in_data), .out_data(bb_8_active_in_state_9_out_data));

	reg [31:0] bb_8_predecessor_in_state_9_in_data;
	wire [31:0] bb_8_predecessor_in_state_9_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor_in_state_9(.in_data(bb_8_predecessor_in_state_9_in_data), .out_data(bb_8_predecessor_in_state_9_out_data));

	reg [31:0] data_in_1_1_in_data;
	wire [31:0] data_in_1_1_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_1(.in_data(data_in_1_1_in_data), .out_data(data_in_1_1_out_data));

	reg [31:0] data_in_1_3_in_data;
	wire [31:0] data_in_1_3_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_3(.in_data(data_in_1_3_in_data), .out_data(data_in_1_3_out_data));

	reg [31:0] data_in_1_5_in_data;
	wire [31:0] data_in_1_5_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_5(.in_data(data_in_1_5_in_data), .out_data(data_in_1_5_out_data));

	reg [31:0] data_in_2_7_in_data;
	wire [31:0] data_in_2_7_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_7(.in_data(data_in_2_7_in_data), .out_data(data_in_2_7_out_data));

	reg [31:0] data_in_2_9_in_data;
	wire [31:0] data_in_2_9_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_9(.in_data(data_in_2_9_in_data), .out_data(data_in_2_9_out_data));

	reg [31:0] data_in_2_11_in_data;
	wire [31:0] data_in_2_11_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_11(.in_data(data_in_2_11_in_data), .out_data(data_in_2_11_out_data));

	reg [31:0] data_in_3_13_in_data;
	wire [31:0] data_in_3_13_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_13(.in_data(data_in_3_13_in_data), .out_data(data_in_3_13_out_data));

	reg [31:0] data_in_3_15_in_data;
	wire [31:0] data_in_3_15_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_15(.in_data(data_in_3_15_in_data), .out_data(data_in_3_15_out_data));

	reg [31:0] data_in_3_17_in_data;
	wire [31:0] data_in_3_17_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_17(.in_data(data_in_3_17_in_data), .out_data(data_in_3_17_out_data));

	reg [31:0] data_in_4_19_in_data;
	wire [31:0] data_in_4_19_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_19(.in_data(data_in_4_19_in_data), .out_data(data_in_4_19_out_data));

	reg [31:0] data_in_4_21_in_data;
	wire [31:0] data_in_4_21_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_21(.in_data(data_in_4_21_in_data), .out_data(data_in_4_21_out_data));

	reg [31:0] data_in_4_23_in_data;
	wire [31:0] data_in_4_23_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_23(.in_data(data_in_4_23_in_data), .out_data(data_in_4_23_out_data));

	reg [31:0] data_in_5_25_in_data;
	wire [31:0] data_in_5_25_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_25(.in_data(data_in_5_25_in_data), .out_data(data_in_5_25_out_data));

	reg [31:0] data_in_5_27_in_data;
	wire [31:0] data_in_5_27_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_27(.in_data(data_in_5_27_in_data), .out_data(data_in_5_27_out_data));

	reg [31:0] data_in_5_29_in_data;
	wire [31:0] data_in_5_29_out_data;
	hls_wire #(.WIDTH(32)) data_in_5_29(.in_data(data_in_5_29_in_data), .out_data(data_in_5_29_out_data));

	reg [31:0] data_in_6_31_in_data;
	wire [31:0] data_in_6_31_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_31(.in_data(data_in_6_31_in_data), .out_data(data_in_6_31_out_data));

	reg [31:0] data_in_6_33_in_data;
	wire [31:0] data_in_6_33_out_data;
	hls_wire #(.WIDTH(32)) data_in_6_33(.in_data(data_in_6_33_in_data), .out_data(data_in_6_33_out_data));

	reg [31:0] data_in_7_35_in_data;
	wire [31:0] data_in_7_35_out_data;
	hls_wire #(.WIDTH(32)) data_in_7_35(.in_data(data_in_7_35_in_data), .out_data(data_in_7_35_out_data));

	reg [31:0] data_in_7_37_in_data;
	wire [31:0] data_in_7_37_out_data;
	hls_wire #(.WIDTH(32)) data_in_7_37(.in_data(data_in_7_37_in_data), .out_data(data_in_7_37_out_data));

	reg [31:0] data_in_8_39_in_data;
	wire [31:0] data_in_8_39_out_data;
	hls_wire #(.WIDTH(32)) data_in_8_39(.in_data(data_in_8_39_in_data), .out_data(data_in_8_39_out_data));

	reg [31:0] data_in_8_41_in_data;
	wire [31:0] data_in_8_41_out_data;
	hls_wire #(.WIDTH(32)) data_in_8_41(.in_data(data_in_8_41_in_data), .out_data(data_in_8_41_out_data));

	wire [0:0] andOp_42_in0;
	wire [0:0] andOp_42_in1;
	wire [0:0] andOp_42_out;
	andOp #(.WIDTH(1)) andOp_42(.in0(andOp_42_in0), .in1(andOp_42_in1), .out(andOp_42_out));

	wire [0:0] notOp_43_in0;
	wire [0:0] notOp_43_out;
	notOp #(.WIDTH(1)) notOp_43(.in(notOp_43_in0), .out(notOp_43_out));

	wire [0:0] andOp_44_in0;
	wire [0:0] andOp_44_in1;
	wire [0:0] andOp_44_out;
	andOp #(.WIDTH(1)) andOp_44(.in0(andOp_44_in0), .in1(andOp_44_in1), .out(andOp_44_out));

	wire [0:0] notOp_45_in0;
	wire [0:0] notOp_45_out;
	notOp #(.WIDTH(1)) notOp_45(.in(notOp_45_in0), .out(notOp_45_out));

	wire [0:0] andOp_46_in0;
	wire [0:0] andOp_46_in1;
	wire [0:0] andOp_46_out;
	andOp #(.WIDTH(1)) andOp_46(.in0(andOp_46_in0), .in1(andOp_46_in1), .out(andOp_46_out));

	wire [0:0] notOp_47_in0;
	wire [0:0] notOp_47_out;
	notOp #(.WIDTH(1)) notOp_47(.in(notOp_47_in0), .out(notOp_47_out));

	wire [0:0] andOp_48_in0;
	wire [0:0] andOp_48_in1;
	wire [0:0] andOp_48_out;
	andOp #(.WIDTH(1)) andOp_48(.in0(andOp_48_in0), .in1(andOp_48_in1), .out(andOp_48_out));

	wire [0:0] notOp_49_in0;
	wire [0:0] notOp_49_out;
	notOp #(.WIDTH(1)) notOp_49(.in(notOp_49_in0), .out(notOp_49_out));

	wire [0:0] andOp_50_in0;
	wire [0:0] andOp_50_in1;
	wire [0:0] andOp_50_out;
	andOp #(.WIDTH(1)) andOp_50(.in0(andOp_50_in0), .in1(andOp_50_in1), .out(andOp_50_out));

	wire [0:0] notOp_51_in0;
	wire [0:0] notOp_51_out;
	notOp #(.WIDTH(1)) notOp_51(.in(notOp_51_in0), .out(notOp_51_out));

	wire [0:0] andOp_52_in0;
	wire [0:0] andOp_52_in1;
	wire [0:0] andOp_52_out;
	andOp #(.WIDTH(1)) andOp_52(.in0(andOp_52_in0), .in1(andOp_52_in1), .out(andOp_52_out));

	wire [0:0] andOp_53_in0;
	wire [0:0] andOp_53_in1;
	wire [0:0] andOp_53_out;
	andOp #(.WIDTH(1)) andOp_53(.in0(andOp_53_in0), .in1(andOp_53_in1), .out(andOp_53_out));

	wire [0:0] notOp_54_in0;
	wire [0:0] notOp_54_out;
	notOp #(.WIDTH(1)) notOp_54(.in(notOp_54_in0), .out(notOp_54_out));

	wire [0:0] andOp_55_in0;
	wire [0:0] andOp_55_in1;
	wire [0:0] andOp_55_out;
	andOp #(.WIDTH(1)) andOp_55(.in0(andOp_55_in0), .in1(andOp_55_in1), .out(andOp_55_out));

	wire [0:0] notOp_56_in0;
	wire [0:0] notOp_56_out;
	notOp #(.WIDTH(1)) notOp_56(.in(notOp_56_in0), .out(notOp_56_out));

	wire [0:0] andOp_57_in0;
	wire [0:0] andOp_57_in1;
	wire [0:0] andOp_57_out;
	andOp #(.WIDTH(1)) andOp_57(.in0(andOp_57_in0), .in1(andOp_57_in1), .out(andOp_57_out));

	wire [0:0] notOp_58_in0;
	wire [0:0] notOp_58_out;
	notOp #(.WIDTH(1)) notOp_58(.in(notOp_58_in0), .out(notOp_58_out));

	wire [0:0] andOp_59_in0;
	wire [0:0] andOp_59_in1;
	wire [0:0] andOp_59_out;
	andOp #(.WIDTH(1)) andOp_59(.in0(andOp_59_in0), .in1(andOp_59_in1), .out(andOp_59_out));

	wire [0:0] notOp_60_in0;
	wire [0:0] notOp_60_out;
	notOp #(.WIDTH(1)) notOp_60(.in(notOp_60_in0), .out(notOp_60_out));

	wire [0:0] andOp_61_in0;
	wire [0:0] andOp_61_in1;
	wire [0:0] andOp_61_out;
	andOp #(.WIDTH(1)) andOp_61(.in0(andOp_61_in0), .in1(andOp_61_in1), .out(andOp_61_out));

	wire [0:0] notOp_62_in0;
	wire [0:0] notOp_62_out;
	notOp #(.WIDTH(1)) notOp_62(.in(notOp_62_in0), .out(notOp_62_out));

	wire [0:0] andOp_63_in0;
	wire [0:0] andOp_63_in1;
	wire [0:0] andOp_63_out;
	andOp #(.WIDTH(1)) andOp_63(.in0(andOp_63_in0), .in1(andOp_63_in1), .out(andOp_63_out));

	wire [0:0] andOp_64_in0;
	wire [0:0] andOp_64_in1;
	wire [0:0] andOp_64_out;
	andOp #(.WIDTH(1)) andOp_64(.in0(andOp_64_in0), .in1(andOp_64_in1), .out(andOp_64_out));

	wire [0:0] notOp_65_in0;
	wire [0:0] notOp_65_out;
	notOp #(.WIDTH(1)) notOp_65(.in(notOp_65_in0), .out(notOp_65_out));

	wire [0:0] andOp_66_in0;
	wire [0:0] andOp_66_in1;
	wire [0:0] andOp_66_out;
	andOp #(.WIDTH(1)) andOp_66(.in0(andOp_66_in0), .in1(andOp_66_in1), .out(andOp_66_out));

	wire [0:0] notOp_67_in0;
	wire [0:0] notOp_67_out;
	notOp #(.WIDTH(1)) notOp_67(.in(notOp_67_in0), .out(notOp_67_out));

	wire [0:0] andOp_68_in0;
	wire [0:0] andOp_68_in1;
	wire [0:0] andOp_68_out;
	andOp #(.WIDTH(1)) andOp_68(.in0(andOp_68_in0), .in1(andOp_68_in1), .out(andOp_68_out));

	wire [0:0] notOp_69_in0;
	wire [0:0] notOp_69_out;
	notOp #(.WIDTH(1)) notOp_69(.in(notOp_69_in0), .out(notOp_69_out));

	wire [0:0] andOp_70_in0;
	wire [0:0] andOp_70_in1;
	wire [0:0] andOp_70_out;
	andOp #(.WIDTH(1)) andOp_70(.in0(andOp_70_in0), .in1(andOp_70_in1), .out(andOp_70_out));

	wire [0:0] notOp_71_in0;
	wire [0:0] notOp_71_out;
	notOp #(.WIDTH(1)) notOp_71(.in(notOp_71_in0), .out(notOp_71_out));

	wire [0:0] andOp_72_in0;
	wire [0:0] andOp_72_in1;
	wire [0:0] andOp_72_out;
	andOp #(.WIDTH(1)) andOp_72(.in0(andOp_72_in0), .in1(andOp_72_in1), .out(andOp_72_out));

	wire [0:0] andOp_73_in0;
	wire [0:0] andOp_73_in1;
	wire [0:0] andOp_73_out;
	andOp #(.WIDTH(1)) andOp_73(.in0(andOp_73_in0), .in1(andOp_73_in1), .out(andOp_73_out));

	wire [0:0] notOp_74_in0;
	wire [0:0] notOp_74_out;
	notOp #(.WIDTH(1)) notOp_74(.in(notOp_74_in0), .out(notOp_74_out));

	wire [0:0] andOp_75_in0;
	wire [0:0] andOp_75_in1;
	wire [0:0] andOp_75_out;
	andOp #(.WIDTH(1)) andOp_75(.in0(andOp_75_in0), .in1(andOp_75_in1), .out(andOp_75_out));

	wire [0:0] notOp_76_in0;
	wire [0:0] notOp_76_out;
	notOp #(.WIDTH(1)) notOp_76(.in(notOp_76_in0), .out(notOp_76_out));

	wire [0:0] andOp_77_in0;
	wire [0:0] andOp_77_in1;
	wire [0:0] andOp_77_out;
	andOp #(.WIDTH(1)) andOp_77(.in0(andOp_77_in0), .in1(andOp_77_in1), .out(andOp_77_out));

	wire [0:0] notOp_78_in0;
	wire [0:0] notOp_78_out;
	notOp #(.WIDTH(1)) notOp_78(.in(notOp_78_in0), .out(notOp_78_out));

	wire [0:0] andOp_79_in0;
	wire [0:0] andOp_79_in1;
	wire [0:0] andOp_79_out;
	andOp #(.WIDTH(1)) andOp_79(.in0(andOp_79_in0), .in1(andOp_79_in1), .out(andOp_79_out));

	wire [0:0] andOp_80_in0;
	wire [0:0] andOp_80_in1;
	wire [0:0] andOp_80_out;
	andOp #(.WIDTH(1)) andOp_80(.in0(andOp_80_in0), .in1(andOp_80_in1), .out(andOp_80_out));

	wire [0:0] notOp_81_in0;
	wire [0:0] notOp_81_out;
	notOp #(.WIDTH(1)) notOp_81(.in(notOp_81_in0), .out(notOp_81_out));

	wire [0:0] andOp_82_in0;
	wire [0:0] andOp_82_in1;
	wire [0:0] andOp_82_out;
	andOp #(.WIDTH(1)) andOp_82(.in0(andOp_82_in0), .in1(andOp_82_in1), .out(andOp_82_out));

	wire [0:0] notOp_83_in0;
	wire [0:0] notOp_83_out;
	notOp #(.WIDTH(1)) notOp_83(.in(notOp_83_in0), .out(notOp_83_out));

	wire [0:0] andOp_84_in0;
	wire [0:0] andOp_84_in1;
	wire [0:0] andOp_84_out;
	andOp #(.WIDTH(1)) andOp_84(.in0(andOp_84_in0), .in1(andOp_84_in1), .out(andOp_84_out));

	wire [0:0] notOp_85_in0;
	wire [0:0] notOp_85_out;
	notOp #(.WIDTH(1)) notOp_85(.in(notOp_85_in0), .out(notOp_85_out));

	wire [0:0] andOp_86_in0;
	wire [0:0] andOp_86_in1;
	wire [0:0] andOp_86_out;
	andOp #(.WIDTH(1)) andOp_86(.in0(andOp_86_in0), .in1(andOp_86_in1), .out(andOp_86_out));

	wire [0:0] notOp_87_in0;
	wire [0:0] notOp_87_out;
	notOp #(.WIDTH(1)) notOp_87(.in(notOp_87_in0), .out(notOp_87_out));

	wire [0:0] andOp_88_in0;
	wire [0:0] andOp_88_in1;
	wire [0:0] andOp_88_out;
	andOp #(.WIDTH(1)) andOp_88(.in0(andOp_88_in0), .in1(andOp_88_in1), .out(andOp_88_out));

	wire [0:0] notOp_89_in0;
	wire [0:0] notOp_89_out;
	notOp #(.WIDTH(1)) notOp_89(.in(notOp_89_in0), .out(notOp_89_out));

	wire [0:0] andOp_90_in0;
	wire [0:0] andOp_90_in1;
	wire [0:0] andOp_90_out;
	andOp #(.WIDTH(1)) andOp_90(.in0(andOp_90_in0), .in1(andOp_90_in1), .out(andOp_90_out));

	wire [0:0] notOp_91_in0;
	wire [0:0] notOp_91_out;
	notOp #(.WIDTH(1)) notOp_91(.in(notOp_91_in0), .out(notOp_91_out));

	wire [0:0] andOp_92_in0;
	wire [0:0] andOp_92_in1;
	wire [0:0] andOp_92_out;
	andOp #(.WIDTH(1)) andOp_92(.in0(andOp_92_in0), .in1(andOp_92_in1), .out(andOp_92_out));

	wire [0:0] notOp_93_in0;
	wire [0:0] notOp_93_out;
	notOp #(.WIDTH(1)) notOp_93(.in(notOp_93_in0), .out(notOp_93_out));

	wire [0:0] andOp_94_in0;
	wire [0:0] andOp_94_in1;
	wire [0:0] andOp_94_out;
	andOp #(.WIDTH(1)) andOp_94(.in0(andOp_94_in0), .in1(andOp_94_in1), .out(andOp_94_out));

	wire [0:0] andOp_95_in0;
	wire [0:0] andOp_95_in1;
	wire [0:0] andOp_95_out;
	andOp #(.WIDTH(1)) andOp_95(.in0(andOp_95_in0), .in1(andOp_95_in1), .out(andOp_95_out));

	wire [0:0] notOp_96_in0;
	wire [0:0] notOp_96_out;
	notOp #(.WIDTH(1)) notOp_96(.in(notOp_96_in0), .out(notOp_96_out));

	wire [0:0] andOp_97_in0;
	wire [0:0] andOp_97_in1;
	wire [0:0] andOp_97_out;
	andOp #(.WIDTH(1)) andOp_97(.in0(andOp_97_in0), .in1(andOp_97_in1), .out(andOp_97_out));

	wire [0:0] notOp_98_in0;
	wire [0:0] notOp_98_out;
	notOp #(.WIDTH(1)) notOp_98(.in(notOp_98_in0), .out(notOp_98_out));

	wire [0:0] andOp_99_in0;
	wire [0:0] andOp_99_in1;
	wire [0:0] andOp_99_out;
	andOp #(.WIDTH(1)) andOp_99(.in0(andOp_99_in0), .in1(andOp_99_in1), .out(andOp_99_out));

	wire [0:0] notOp_100_in0;
	wire [0:0] notOp_100_out;
	notOp #(.WIDTH(1)) notOp_100(.in(notOp_100_in0), .out(notOp_100_out));

	wire [0:0] andOp_101_in0;
	wire [0:0] andOp_101_in1;
	wire [0:0] andOp_101_out;
	andOp #(.WIDTH(1)) andOp_101(.in0(andOp_101_in0), .in1(andOp_101_in1), .out(andOp_101_out));

	wire [0:0] andOp_102_in0;
	wire [0:0] andOp_102_in1;
	wire [0:0] andOp_102_out;
	andOp #(.WIDTH(1)) andOp_102(.in0(andOp_102_in0), .in1(andOp_102_in1), .out(andOp_102_out));

	wire [0:0] notOp_103_in0;
	wire [0:0] notOp_103_out;
	notOp #(.WIDTH(1)) notOp_103(.in(notOp_103_in0), .out(notOp_103_out));

	wire [0:0] andOp_104_in0;
	wire [0:0] andOp_104_in1;
	wire [0:0] andOp_104_out;
	andOp #(.WIDTH(1)) andOp_104(.in0(andOp_104_in0), .in1(andOp_104_in1), .out(andOp_104_out));

	wire [0:0] notOp_105_in0;
	wire [0:0] notOp_105_out;
	notOp #(.WIDTH(1)) notOp_105(.in(notOp_105_in0), .out(notOp_105_out));

	wire [0:0] andOp_106_in0;
	wire [0:0] andOp_106_in1;
	wire [0:0] andOp_106_out;
	andOp #(.WIDTH(1)) andOp_106(.in0(andOp_106_in0), .in1(andOp_106_in1), .out(andOp_106_out));

	wire [0:0] notOp_107_in0;
	wire [0:0] notOp_107_out;
	notOp #(.WIDTH(1)) notOp_107(.in(notOp_107_in0), .out(notOp_107_out));

	wire [0:0] andOp_108_in0;
	wire [0:0] andOp_108_in1;
	wire [0:0] andOp_108_out;
	andOp #(.WIDTH(1)) andOp_108(.in0(andOp_108_in0), .in1(andOp_108_in1), .out(andOp_108_out));

	wire [0:0] notOp_109_in0;
	wire [0:0] notOp_109_out;
	notOp #(.WIDTH(1)) notOp_109(.in(notOp_109_in0), .out(notOp_109_out));

	wire [0:0] andOp_110_in0;
	wire [0:0] andOp_110_in1;
	wire [0:0] andOp_110_out;
	andOp #(.WIDTH(1)) andOp_110(.in0(andOp_110_in0), .in1(andOp_110_in1), .out(andOp_110_out));

	wire [0:0] notOp_111_in0;
	wire [0:0] notOp_111_out;
	notOp #(.WIDTH(1)) notOp_111(.in(notOp_111_in0), .out(notOp_111_out));

	wire [0:0] andOp_112_in0;
	wire [0:0] andOp_112_in1;
	wire [0:0] andOp_112_out;
	andOp #(.WIDTH(1)) andOp_112(.in0(andOp_112_in0), .in1(andOp_112_in1), .out(andOp_112_out));

	wire [0:0] andOp_113_in0;
	wire [0:0] andOp_113_in1;
	wire [0:0] andOp_113_out;
	andOp #(.WIDTH(1)) andOp_113(.in0(andOp_113_in0), .in1(andOp_113_in1), .out(andOp_113_out));

	wire [0:0] notOp_114_in0;
	wire [0:0] notOp_114_out;
	notOp #(.WIDTH(1)) notOp_114(.in(notOp_114_in0), .out(notOp_114_out));

	wire [31:0] eq_115_in0;
	wire [31:0] eq_115_in1;
	wire [0:0] eq_115_out;
	eq #(.WIDTH(32)) eq_115(.in0(eq_115_in0), .in1(eq_115_in1), .out(eq_115_out));

	wire [31:0] eq_116_in0;
	wire [31:0] eq_116_in1;
	wire [0:0] eq_116_out;
	eq #(.WIDTH(32)) eq_116(.in0(eq_116_in0), .in1(eq_116_in1), .out(eq_116_out));

	wire [0:0] orOp_117_in0;
	wire [0:0] orOp_117_in1;
	wire [0:0] orOp_117_out;
	orOp #(.WIDTH(1)) orOp_117(.in0(orOp_117_in0), .in1(orOp_117_in1), .out(orOp_117_out));

	wire [31:0] eq_118_in0;
	wire [31:0] eq_118_in1;
	wire [0:0] eq_118_out;
	eq #(.WIDTH(32)) eq_118(.in0(eq_118_in0), .in1(eq_118_in1), .out(eq_118_out));

	wire [31:0] eq_119_in0;
	wire [31:0] eq_119_in1;
	wire [0:0] eq_119_out;
	eq #(.WIDTH(32)) eq_119(.in0(eq_119_in0), .in1(eq_119_in1), .out(eq_119_out));

	wire [0:0] orOp_120_in0;
	wire [0:0] orOp_120_in1;
	wire [0:0] orOp_120_out;
	orOp #(.WIDTH(1)) orOp_120(.in0(orOp_120_in0), .in1(orOp_120_in1), .out(orOp_120_out));

	wire [31:0] eq_121_in0;
	wire [31:0] eq_121_in1;
	wire [0:0] eq_121_out;
	eq #(.WIDTH(32)) eq_121(.in0(eq_121_in0), .in1(eq_121_in1), .out(eq_121_out));

	wire [31:0] eq_122_in0;
	wire [31:0] eq_122_in1;
	wire [0:0] eq_122_out;
	eq #(.WIDTH(32)) eq_122(.in0(eq_122_in0), .in1(eq_122_in1), .out(eq_122_out));

	wire [31:0] eq_123_in0;
	wire [31:0] eq_123_in1;
	wire [0:0] eq_123_out;
	eq #(.WIDTH(32)) eq_123(.in0(eq_123_in0), .in1(eq_123_in1), .out(eq_123_out));

	wire [0:0] orOp_124_in0;
	wire [0:0] orOp_124_in1;
	wire [0:0] orOp_124_out;
	orOp #(.WIDTH(1)) orOp_124(.in0(orOp_124_in0), .in1(orOp_124_in1), .out(orOp_124_out));

	wire [31:0] eq_125_in0;
	wire [31:0] eq_125_in1;
	wire [0:0] eq_125_out;
	eq #(.WIDTH(32)) eq_125(.in0(eq_125_in0), .in1(eq_125_in1), .out(eq_125_out));

	wire [0:0] orOp_126_in0;
	wire [0:0] orOp_126_in1;
	wire [0:0] orOp_126_out;
	orOp #(.WIDTH(1)) orOp_126(.in0(orOp_126_in0), .in1(orOp_126_in1), .out(orOp_126_out));

	wire [31:0] eq_127_in0;
	wire [31:0] eq_127_in1;
	wire [0:0] eq_127_out;
	eq #(.WIDTH(32)) eq_127(.in0(eq_127_in0), .in1(eq_127_in1), .out(eq_127_out));

	wire [0:0] orOp_128_in0;
	wire [0:0] orOp_128_in1;
	wire [0:0] orOp_128_out;
	orOp #(.WIDTH(1)) orOp_128(.in0(orOp_128_in0), .in1(orOp_128_in1), .out(orOp_128_out));

	wire [31:0] eq_129_in0;
	wire [31:0] eq_129_in1;
	wire [0:0] eq_129_out;
	eq #(.WIDTH(32)) eq_129(.in0(eq_129_in0), .in1(eq_129_in1), .out(eq_129_out));

	wire [31:0] eq_130_in0;
	wire [31:0] eq_130_in1;
	wire [0:0] eq_130_out;
	eq #(.WIDTH(32)) eq_130(.in0(eq_130_in0), .in1(eq_130_in1), .out(eq_130_out));

	wire [0:0] orOp_131_in0;
	wire [0:0] orOp_131_in1;
	wire [0:0] orOp_131_out;
	orOp #(.WIDTH(1)) orOp_131(.in0(orOp_131_in0), .in1(orOp_131_in1), .out(orOp_131_out));

	wire [31:0] eq_132_in0;
	wire [31:0] eq_132_in1;
	wire [0:0] eq_132_out;
	eq #(.WIDTH(32)) eq_132(.in0(eq_132_in0), .in1(eq_132_in1), .out(eq_132_out));

	wire [0:0] orOp_133_in0;
	wire [0:0] orOp_133_in1;
	wire [0:0] orOp_133_out;
	orOp #(.WIDTH(1)) orOp_133(.in0(orOp_133_in0), .in1(orOp_133_in1), .out(orOp_133_out));

	wire [31:0] eq_134_in0;
	wire [31:0] eq_134_in1;
	wire [0:0] eq_134_out;
	eq #(.WIDTH(32)) eq_134(.in0(eq_134_in0), .in1(eq_134_in1), .out(eq_134_out));

	wire [0:0] orOp_135_in0;
	wire [0:0] orOp_135_in1;
	wire [0:0] orOp_135_out;
	orOp #(.WIDTH(1)) orOp_135(.in0(orOp_135_in0), .in1(orOp_135_in1), .out(orOp_135_out));

	wire [31:0] eq_136_in0;
	wire [31:0] eq_136_in1;
	wire [0:0] eq_136_out;
	eq #(.WIDTH(32)) eq_136(.in0(eq_136_in0), .in1(eq_136_in1), .out(eq_136_out));

	wire [0:0] orOp_137_in0;
	wire [0:0] orOp_137_in1;
	wire [0:0] orOp_137_out;
	orOp #(.WIDTH(1)) orOp_137(.in0(orOp_137_in0), .in1(orOp_137_in1), .out(orOp_137_out));

	wire [31:0] eq_138_in0;
	wire [31:0] eq_138_in1;
	wire [0:0] eq_138_out;
	eq #(.WIDTH(32)) eq_138(.in0(eq_138_in0), .in1(eq_138_in1), .out(eq_138_out));

	wire [31:0] eq_139_in0;
	wire [31:0] eq_139_in1;
	wire [0:0] eq_139_out;
	eq #(.WIDTH(32)) eq_139(.in0(eq_139_in0), .in1(eq_139_in1), .out(eq_139_out));

	wire [0:0] orOp_140_in0;
	wire [0:0] orOp_140_in1;
	wire [0:0] orOp_140_out;
	orOp #(.WIDTH(1)) orOp_140(.in0(orOp_140_in0), .in1(orOp_140_in1), .out(orOp_140_out));

	wire [31:0] eq_141_in0;
	wire [31:0] eq_141_in1;
	wire [0:0] eq_141_out;
	eq #(.WIDTH(32)) eq_141(.in0(eq_141_in0), .in1(eq_141_in1), .out(eq_141_out));

	wire [0:0] orOp_142_in0;
	wire [0:0] orOp_142_in1;
	wire [0:0] orOp_142_out;
	orOp #(.WIDTH(1)) orOp_142(.in0(orOp_142_in0), .in1(orOp_142_in1), .out(orOp_142_out));

	wire [31:0] eq_143_in0;
	wire [31:0] eq_143_in1;
	wire [0:0] eq_143_out;
	eq #(.WIDTH(32)) eq_143(.in0(eq_143_in0), .in1(eq_143_in1), .out(eq_143_out));

	wire [31:0] eq_144_in0;
	wire [31:0] eq_144_in1;
	wire [0:0] eq_144_out;
	eq #(.WIDTH(32)) eq_144(.in0(eq_144_in0), .in1(eq_144_in1), .out(eq_144_out));

	wire [0:0] orOp_145_in0;
	wire [0:0] orOp_145_in1;
	wire [0:0] orOp_145_out;
	orOp #(.WIDTH(1)) orOp_145(.in0(orOp_145_in0), .in1(orOp_145_in1), .out(orOp_145_out));

	wire [31:0] eq_146_in0;
	wire [31:0] eq_146_in1;
	wire [0:0] eq_146_out;
	eq #(.WIDTH(32)) eq_146(.in0(eq_146_in0), .in1(eq_146_in1), .out(eq_146_out));

	wire [31:0] eq_147_in0;
	wire [31:0] eq_147_in1;
	wire [0:0] eq_147_out;
	eq #(.WIDTH(32)) eq_147(.in0(eq_147_in0), .in1(eq_147_in1), .out(eq_147_out));

	wire [0:0] orOp_148_in0;
	wire [0:0] orOp_148_in1;
	wire [0:0] orOp_148_out;
	orOp #(.WIDTH(1)) orOp_148(.in0(orOp_148_in0), .in1(orOp_148_in1), .out(orOp_148_out));

	wire [31:0] eq_149_in0;
	wire [31:0] eq_149_in1;
	wire [0:0] eq_149_out;
	eq #(.WIDTH(32)) eq_149(.in0(eq_149_in0), .in1(eq_149_in1), .out(eq_149_out));

	wire [0:0] orOp_150_in0;
	wire [0:0] orOp_150_in1;
	wire [0:0] orOp_150_out;
	orOp #(.WIDTH(1)) orOp_150(.in0(orOp_150_in0), .in1(orOp_150_in1), .out(orOp_150_out));

	wire [31:0] eq_151_in0;
	wire [31:0] eq_151_in1;
	wire [0:0] eq_151_out;
	eq #(.WIDTH(32)) eq_151(.in0(eq_151_in0), .in1(eq_151_in1), .out(eq_151_out));

	wire [0:0] orOp_152_in0;
	wire [0:0] orOp_152_in1;
	wire [0:0] orOp_152_out;
	orOp #(.WIDTH(1)) orOp_152(.in0(orOp_152_in0), .in1(orOp_152_in1), .out(orOp_152_out));

	wire [31:0] eq_153_in0;
	wire [31:0] eq_153_in1;
	wire [0:0] eq_153_out;
	eq #(.WIDTH(32)) eq_153(.in0(eq_153_in0), .in1(eq_153_in1), .out(eq_153_out));

	wire [31:0] eq_154_in0;
	wire [31:0] eq_154_in1;
	wire [0:0] eq_154_out;
	eq #(.WIDTH(32)) eq_154(.in0(eq_154_in0), .in1(eq_154_in1), .out(eq_154_out));

	wire [0:0] orOp_155_in0;
	wire [0:0] orOp_155_in1;
	wire [0:0] orOp_155_out;
	orOp #(.WIDTH(1)) orOp_155(.in0(orOp_155_in0), .in1(orOp_155_in1), .out(orOp_155_out));

	wire [31:0] eq_156_in0;
	wire [31:0] eq_156_in1;
	wire [0:0] eq_156_out;
	eq #(.WIDTH(32)) eq_156(.in0(eq_156_in0), .in1(eq_156_in1), .out(eq_156_out));

	wire [0:0] orOp_157_in0;
	wire [0:0] orOp_157_in1;
	wire [0:0] orOp_157_out;
	orOp #(.WIDTH(1)) orOp_157(.in0(orOp_157_in0), .in1(orOp_157_in1), .out(orOp_157_out));

	wire [31:0] eq_158_in0;
	wire [31:0] eq_158_in1;
	wire [0:0] eq_158_out;
	eq #(.WIDTH(32)) eq_158(.in0(eq_158_in0), .in1(eq_158_in1), .out(eq_158_out));

	wire [31:0] eq_159_in0;
	wire [31:0] eq_159_in1;
	wire [0:0] eq_159_out;
	eq #(.WIDTH(32)) eq_159(.in0(eq_159_in0), .in1(eq_159_in1), .out(eq_159_out));

	wire [31:0] eq_160_in0;
	wire [31:0] eq_160_in1;
	wire [0:0] eq_160_out;
	eq #(.WIDTH(32)) eq_160(.in0(eq_160_in0), .in1(eq_160_in1), .out(eq_160_out));

	wire [0:0] notOp_161_in0;
	wire [0:0] notOp_161_out;
	notOp #(.WIDTH(1)) notOp_161(.in(notOp_161_in0), .out(notOp_161_out));

	wire [0:0] andOp_162_in0;
	wire [0:0] andOp_162_in1;
	wire [0:0] andOp_162_out;
	andOp #(.WIDTH(1)) andOp_162(.in0(andOp_162_in0), .in1(andOp_162_in1), .out(andOp_162_out));

	wire [31:0] eq_163_in0;
	wire [31:0] eq_163_in1;
	wire [0:0] eq_163_out;
	eq #(.WIDTH(32)) eq_163(.in0(eq_163_in0), .in1(eq_163_in1), .out(eq_163_out));

	wire [31:0] eq_164_in0;
	wire [31:0] eq_164_in1;
	wire [0:0] eq_164_out;
	eq #(.WIDTH(32)) eq_164(.in0(eq_164_in0), .in1(eq_164_in1), .out(eq_164_out));

	wire [0:0] notOp_165_in0;
	wire [0:0] notOp_165_out;
	notOp #(.WIDTH(1)) notOp_165(.in(notOp_165_in0), .out(notOp_165_out));

	wire [0:0] andOp_166_in0;
	wire [0:0] andOp_166_in1;
	wire [0:0] andOp_166_out;
	andOp #(.WIDTH(1)) andOp_166(.in0(andOp_166_in0), .in1(andOp_166_in1), .out(andOp_166_out));

	wire [31:0] eq_167_in0;
	wire [31:0] eq_167_in1;
	wire [0:0] eq_167_out;
	eq #(.WIDTH(32)) eq_167(.in0(eq_167_in0), .in1(eq_167_in1), .out(eq_167_out));

	wire [31:0] eq_168_in0;
	wire [31:0] eq_168_in1;
	wire [0:0] eq_168_out;
	eq #(.WIDTH(32)) eq_168(.in0(eq_168_in0), .in1(eq_168_in1), .out(eq_168_out));

	wire [31:0] eq_169_in0;
	wire [31:0] eq_169_in1;
	wire [0:0] eq_169_out;
	eq #(.WIDTH(32)) eq_169(.in0(eq_169_in0), .in1(eq_169_in1), .out(eq_169_out));

	wire [0:0] notOp_170_in0;
	wire [0:0] notOp_170_out;
	notOp #(.WIDTH(1)) notOp_170(.in(notOp_170_in0), .out(notOp_170_out));

	wire [0:0] andOp_171_in0;
	wire [0:0] andOp_171_in1;
	wire [0:0] andOp_171_out;
	andOp #(.WIDTH(1)) andOp_171(.in0(andOp_171_in0), .in1(andOp_171_in1), .out(andOp_171_out));

	wire [31:0] eq_172_in0;
	wire [31:0] eq_172_in1;
	wire [0:0] eq_172_out;
	eq #(.WIDTH(32)) eq_172(.in0(eq_172_in0), .in1(eq_172_in1), .out(eq_172_out));

	wire [0:0] notOp_173_in0;
	wire [0:0] notOp_173_out;
	notOp #(.WIDTH(1)) notOp_173(.in(notOp_173_in0), .out(notOp_173_out));

	wire [0:0] andOp_174_in0;
	wire [0:0] andOp_174_in1;
	wire [0:0] andOp_174_out;
	andOp #(.WIDTH(1)) andOp_174(.in0(andOp_174_in0), .in1(andOp_174_in1), .out(andOp_174_out));

	wire [31:0] eq_175_in0;
	wire [31:0] eq_175_in1;
	wire [0:0] eq_175_out;
	eq #(.WIDTH(32)) eq_175(.in0(eq_175_in0), .in1(eq_175_in1), .out(eq_175_out));

	wire [0:0] notOp_176_in0;
	wire [0:0] notOp_176_out;
	notOp #(.WIDTH(1)) notOp_176(.in(notOp_176_in0), .out(notOp_176_out));

	wire [0:0] andOp_177_in0;
	wire [0:0] andOp_177_in1;
	wire [0:0] andOp_177_out;
	andOp #(.WIDTH(1)) andOp_177(.in0(andOp_177_in0), .in1(andOp_177_in1), .out(andOp_177_out));

	wire [31:0] eq_178_in0;
	wire [31:0] eq_178_in1;
	wire [0:0] eq_178_out;
	eq #(.WIDTH(32)) eq_178(.in0(eq_178_in0), .in1(eq_178_in1), .out(eq_178_out));

	wire [31:0] eq_179_in0;
	wire [31:0] eq_179_in1;
	wire [0:0] eq_179_out;
	eq #(.WIDTH(32)) eq_179(.in0(eq_179_in0), .in1(eq_179_in1), .out(eq_179_out));

	wire [0:0] notOp_180_in0;
	wire [0:0] notOp_180_out;
	notOp #(.WIDTH(1)) notOp_180(.in(notOp_180_in0), .out(notOp_180_out));

	wire [0:0] andOp_181_in0;
	wire [0:0] andOp_181_in1;
	wire [0:0] andOp_181_out;
	andOp #(.WIDTH(1)) andOp_181(.in0(andOp_181_in0), .in1(andOp_181_in1), .out(andOp_181_out));

	wire [31:0] eq_182_in0;
	wire [31:0] eq_182_in1;
	wire [0:0] eq_182_out;
	eq #(.WIDTH(32)) eq_182(.in0(eq_182_in0), .in1(eq_182_in1), .out(eq_182_out));

	wire [0:0] notOp_183_in0;
	wire [0:0] notOp_183_out;
	notOp #(.WIDTH(1)) notOp_183(.in(notOp_183_in0), .out(notOp_183_out));

	wire [0:0] andOp_184_in0;
	wire [0:0] andOp_184_in1;
	wire [0:0] andOp_184_out;
	andOp #(.WIDTH(1)) andOp_184(.in0(andOp_184_in0), .in1(andOp_184_in1), .out(andOp_184_out));

	wire [31:0] eq_185_in0;
	wire [31:0] eq_185_in1;
	wire [0:0] eq_185_out;
	eq #(.WIDTH(32)) eq_185(.in0(eq_185_in0), .in1(eq_185_in1), .out(eq_185_out));

	wire [0:0] notOp_186_in0;
	wire [0:0] notOp_186_out;
	notOp #(.WIDTH(1)) notOp_186(.in(notOp_186_in0), .out(notOp_186_out));

	wire [0:0] andOp_187_in0;
	wire [0:0] andOp_187_in1;
	wire [0:0] andOp_187_out;
	andOp #(.WIDTH(1)) andOp_187(.in0(andOp_187_in0), .in1(andOp_187_in1), .out(andOp_187_out));

	wire [31:0] eq_188_in0;
	wire [31:0] eq_188_in1;
	wire [0:0] eq_188_out;
	eq #(.WIDTH(32)) eq_188(.in0(eq_188_in0), .in1(eq_188_in1), .out(eq_188_out));

	wire [0:0] notOp_189_in0;
	wire [0:0] notOp_189_out;
	notOp #(.WIDTH(1)) notOp_189(.in(notOp_189_in0), .out(notOp_189_out));

	wire [0:0] andOp_190_in0;
	wire [0:0] andOp_190_in1;
	wire [0:0] andOp_190_out;
	andOp #(.WIDTH(1)) andOp_190(.in0(andOp_190_in0), .in1(andOp_190_in1), .out(andOp_190_out));

	wire [31:0] eq_191_in0;
	wire [31:0] eq_191_in1;
	wire [0:0] eq_191_out;
	eq #(.WIDTH(32)) eq_191(.in0(eq_191_in0), .in1(eq_191_in1), .out(eq_191_out));

	wire [31:0] eq_192_in0;
	wire [31:0] eq_192_in1;
	wire [0:0] eq_192_out;
	eq #(.WIDTH(32)) eq_192(.in0(eq_192_in0), .in1(eq_192_in1), .out(eq_192_out));

	wire [0:0] notOp_193_in0;
	wire [0:0] notOp_193_out;
	notOp #(.WIDTH(1)) notOp_193(.in(notOp_193_in0), .out(notOp_193_out));

	wire [0:0] andOp_194_in0;
	wire [0:0] andOp_194_in1;
	wire [0:0] andOp_194_out;
	andOp #(.WIDTH(1)) andOp_194(.in0(andOp_194_in0), .in1(andOp_194_in1), .out(andOp_194_out));

	wire [31:0] eq_195_in0;
	wire [31:0] eq_195_in1;
	wire [0:0] eq_195_out;
	eq #(.WIDTH(32)) eq_195(.in0(eq_195_in0), .in1(eq_195_in1), .out(eq_195_out));

	wire [0:0] notOp_196_in0;
	wire [0:0] notOp_196_out;
	notOp #(.WIDTH(1)) notOp_196(.in(notOp_196_in0), .out(notOp_196_out));

	wire [0:0] andOp_197_in0;
	wire [0:0] andOp_197_in1;
	wire [0:0] andOp_197_out;
	andOp #(.WIDTH(1)) andOp_197(.in0(andOp_197_in0), .in1(andOp_197_in1), .out(andOp_197_out));

	wire [31:0] eq_198_in0;
	wire [31:0] eq_198_in1;
	wire [0:0] eq_198_out;
	eq #(.WIDTH(32)) eq_198(.in0(eq_198_in0), .in1(eq_198_in1), .out(eq_198_out));

	wire [31:0] eq_199_in0;
	wire [31:0] eq_199_in1;
	wire [0:0] eq_199_out;
	eq #(.WIDTH(32)) eq_199(.in0(eq_199_in0), .in1(eq_199_in1), .out(eq_199_out));

	wire [0:0] notOp_200_in0;
	wire [0:0] notOp_200_out;
	notOp #(.WIDTH(1)) notOp_200(.in(notOp_200_in0), .out(notOp_200_out));

	wire [0:0] andOp_201_in0;
	wire [0:0] andOp_201_in1;
	wire [0:0] andOp_201_out;
	andOp #(.WIDTH(1)) andOp_201(.in0(andOp_201_in0), .in1(andOp_201_in1), .out(andOp_201_out));

	wire [31:0] eq_202_in0;
	wire [31:0] eq_202_in1;
	wire [0:0] eq_202_out;
	eq #(.WIDTH(32)) eq_202(.in0(eq_202_in0), .in1(eq_202_in1), .out(eq_202_out));

	wire [31:0] eq_203_in0;
	wire [31:0] eq_203_in1;
	wire [0:0] eq_203_out;
	eq #(.WIDTH(32)) eq_203(.in0(eq_203_in0), .in1(eq_203_in1), .out(eq_203_out));

	wire [0:0] notOp_204_in0;
	wire [0:0] notOp_204_out;
	notOp #(.WIDTH(1)) notOp_204(.in(notOp_204_in0), .out(notOp_204_out));

	wire [0:0] andOp_205_in0;
	wire [0:0] andOp_205_in1;
	wire [0:0] andOp_205_out;
	andOp #(.WIDTH(1)) andOp_205(.in0(andOp_205_in0), .in1(andOp_205_in1), .out(andOp_205_out));

	wire [31:0] eq_206_in0;
	wire [31:0] eq_206_in1;
	wire [0:0] eq_206_out;
	eq #(.WIDTH(32)) eq_206(.in0(eq_206_in0), .in1(eq_206_in1), .out(eq_206_out));

	wire [0:0] notOp_207_in0;
	wire [0:0] notOp_207_out;
	notOp #(.WIDTH(1)) notOp_207(.in(notOp_207_in0), .out(notOp_207_out));

	wire [0:0] andOp_208_in0;
	wire [0:0] andOp_208_in1;
	wire [0:0] andOp_208_out;
	andOp #(.WIDTH(1)) andOp_208(.in0(andOp_208_in0), .in1(andOp_208_in1), .out(andOp_208_out));

	wire [31:0] eq_209_in0;
	wire [31:0] eq_209_in1;
	wire [0:0] eq_209_out;
	eq #(.WIDTH(32)) eq_209(.in0(eq_209_in0), .in1(eq_209_in1), .out(eq_209_out));

	wire [0:0] notOp_210_in0;
	wire [0:0] notOp_210_out;
	notOp #(.WIDTH(1)) notOp_210(.in(notOp_210_in0), .out(notOp_210_out));

	wire [0:0] andOp_211_in0;
	wire [0:0] andOp_211_in1;
	wire [0:0] andOp_211_out;
	andOp #(.WIDTH(1)) andOp_211(.in0(andOp_211_in0), .in1(andOp_211_in1), .out(andOp_211_out));

	wire [31:0] eq_212_in0;
	wire [31:0] eq_212_in1;
	wire [0:0] eq_212_out;
	eq #(.WIDTH(32)) eq_212(.in0(eq_212_in0), .in1(eq_212_in1), .out(eq_212_out));

	wire [31:0] eq_213_in0;
	wire [31:0] eq_213_in1;
	wire [0:0] eq_213_out;
	eq #(.WIDTH(32)) eq_213(.in0(eq_213_in0), .in1(eq_213_in1), .out(eq_213_out));

	wire [0:0] notOp_214_in0;
	wire [0:0] notOp_214_out;
	notOp #(.WIDTH(1)) notOp_214(.in(notOp_214_in0), .out(notOp_214_out));

	wire [0:0] andOp_215_in0;
	wire [0:0] andOp_215_in1;
	wire [0:0] andOp_215_out;
	andOp #(.WIDTH(1)) andOp_215(.in0(andOp_215_in0), .in1(andOp_215_in1), .out(andOp_215_out));

	wire [31:0] eq_216_in0;
	wire [31:0] eq_216_in1;
	wire [0:0] eq_216_out;
	eq #(.WIDTH(32)) eq_216(.in0(eq_216_in0), .in1(eq_216_in1), .out(eq_216_out));

	wire [0:0] notOp_217_in0;
	wire [0:0] notOp_217_out;
	notOp #(.WIDTH(1)) notOp_217(.in(notOp_217_in0), .out(notOp_217_out));

	wire [0:0] andOp_218_in0;
	wire [0:0] andOp_218_in1;
	wire [0:0] andOp_218_out;
	andOp #(.WIDTH(1)) andOp_218(.in0(andOp_218_in0), .in1(andOp_218_in1), .out(andOp_218_out));

	wire [31:0] eq_219_in0;
	wire [31:0] eq_219_in1;
	wire [0:0] eq_219_out;
	eq #(.WIDTH(32)) eq_219(.in0(eq_219_in0), .in1(eq_219_in1), .out(eq_219_out));

	wire [0:0] andOp_220_in0;
	wire [0:0] andOp_220_in1;
	wire [0:0] andOp_220_out;
	andOp #(.WIDTH(1)) andOp_220(.in0(andOp_220_in0), .in1(andOp_220_in1), .out(andOp_220_out));

	wire [0:0] andOp_221_in0;
	wire [0:0] andOp_221_in1;
	wire [0:0] andOp_221_out;
	andOp #(.WIDTH(1)) andOp_221(.in0(andOp_221_in0), .in1(andOp_221_in1), .out(andOp_221_out));

	wire [0:0] andOp_222_in0;
	wire [0:0] andOp_222_in1;
	wire [0:0] andOp_222_out;
	andOp #(.WIDTH(1)) andOp_222(.in0(andOp_222_in0), .in1(andOp_222_in1), .out(andOp_222_out));

	wire [0:0] andOp_223_in0;
	wire [0:0] andOp_223_in1;
	wire [0:0] andOp_223_out;
	andOp #(.WIDTH(1)) andOp_223(.in0(andOp_223_in0), .in1(andOp_223_in1), .out(andOp_223_out));

	reg [31:0] tmp_output_224_in_data;
	wire [31:0] tmp_output_224_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_224(.in_data(tmp_output_224_in_data), .out_data(tmp_output_224_out_data));

	wire [31:0] eq_225_in0;
	wire [31:0] eq_225_in1;
	wire [0:0] eq_225_out;
	eq #(.WIDTH(32)) eq_225(.in0(eq_225_in0), .in1(eq_225_in1), .out(eq_225_out));

	wire [31:0] eq_226_in0;
	wire [31:0] eq_226_in1;
	wire [0:0] eq_226_out;
	eq #(.WIDTH(32)) eq_226(.in0(eq_226_in0), .in1(eq_226_in1), .out(eq_226_out));

	wire [0:0] andOp_227_in0;
	wire [0:0] andOp_227_in1;
	wire [0:0] andOp_227_out;
	andOp #(.WIDTH(1)) andOp_227(.in0(andOp_227_in0), .in1(andOp_227_in1), .out(andOp_227_out));

	wire [0:0] andOp_228_in0;
	wire [0:0] andOp_228_in1;
	wire [0:0] andOp_228_out;
	andOp #(.WIDTH(1)) andOp_228(.in0(andOp_228_in0), .in1(andOp_228_in1), .out(andOp_228_out));

	wire [0:0] andOp_229_in0;
	wire [0:0] andOp_229_in1;
	wire [0:0] andOp_229_out;
	andOp #(.WIDTH(1)) andOp_229(.in0(andOp_229_in0), .in1(andOp_229_in1), .out(andOp_229_out));

	wire [0:0] andOp_230_in0;
	wire [0:0] andOp_230_in1;
	wire [0:0] andOp_230_out;
	andOp #(.WIDTH(1)) andOp_230(.in0(andOp_230_in0), .in1(andOp_230_in1), .out(andOp_230_out));

	wire [31:0] concat_231_in0;
	wire [31:0] concat_231_in1;
	wire [63:0] concat_231_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_231(.in0(concat_231_in0), .in1(concat_231_in1), .out(concat_231_out));

	wire [31:0] concat_232_in0;
	wire [31:0] concat_232_in1;
	wire [63:0] concat_232_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_232(.in0(concat_232_in0), .in1(concat_232_in1), .out(concat_232_out));

	wire [0:0] andOp_233_in0;
	wire [0:0] andOp_233_in1;
	wire [0:0] andOp_233_out;
	andOp #(.WIDTH(1)) andOp_233(.in0(andOp_233_in0), .in1(andOp_233_in1), .out(andOp_233_out));

	wire [0:0] andOp_234_in0;
	wire [0:0] andOp_234_in1;
	wire [0:0] andOp_234_out;
	andOp #(.WIDTH(1)) andOp_234(.in0(andOp_234_in0), .in1(andOp_234_in1), .out(andOp_234_out));

	wire [0:0] andOp_235_in0;
	wire [0:0] andOp_235_in1;
	wire [0:0] andOp_235_out;
	andOp #(.WIDTH(1)) andOp_235(.in0(andOp_235_in0), .in1(andOp_235_in1), .out(andOp_235_out));

	wire [0:0] andOp_236_in0;
	wire [0:0] andOp_236_in1;
	wire [0:0] andOp_236_out;
	andOp #(.WIDTH(1)) andOp_236(.in0(andOp_236_in0), .in1(andOp_236_in1), .out(andOp_236_out));

	wire [0:0] andOp_237_in0;
	wire [0:0] andOp_237_in1;
	wire [0:0] andOp_237_out;
	andOp #(.WIDTH(1)) andOp_237(.in0(andOp_237_in0), .in1(andOp_237_in1), .out(andOp_237_out));

	wire [0:0] andOp_238_in0;
	wire [0:0] andOp_238_in1;
	wire [0:0] andOp_238_out;
	andOp #(.WIDTH(1)) andOp_238(.in0(andOp_238_in0), .in1(andOp_238_in1), .out(andOp_238_out));

	wire [0:0] andOp_239_in0;
	wire [0:0] andOp_239_in1;
	wire [0:0] andOp_239_out;
	andOp #(.WIDTH(1)) andOp_239(.in0(andOp_239_in0), .in1(andOp_239_in1), .out(andOp_239_out));

	wire [0:0] andOp_240_in0;
	wire [0:0] andOp_240_in1;
	wire [0:0] andOp_240_out;
	andOp #(.WIDTH(1)) andOp_240(.in0(andOp_240_in0), .in1(andOp_240_in1), .out(andOp_240_out));

	wire [0:0] andOp_241_in0;
	wire [0:0] andOp_241_in1;
	wire [0:0] andOp_241_out;
	andOp #(.WIDTH(1)) andOp_241(.in0(andOp_241_in0), .in1(andOp_241_in1), .out(andOp_241_out));

	reg [31:0] tmp_output_242_in_data;
	wire [31:0] tmp_output_242_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_242(.in_data(tmp_output_242_in_data), .out_data(tmp_output_242_out_data));

	wire [31:0] eq_243_in0;
	wire [31:0] eq_243_in1;
	wire [0:0] eq_243_out;
	eq #(.WIDTH(32)) eq_243(.in0(eq_243_in0), .in1(eq_243_in1), .out(eq_243_out));

	wire [31:0] eq_244_in0;
	wire [31:0] eq_244_in1;
	wire [0:0] eq_244_out;
	eq #(.WIDTH(32)) eq_244(.in0(eq_244_in0), .in1(eq_244_in1), .out(eq_244_out));

	wire [0:0] andOp_245_in0;
	wire [0:0] andOp_245_in1;
	wire [0:0] andOp_245_out;
	andOp #(.WIDTH(1)) andOp_245(.in0(andOp_245_in0), .in1(andOp_245_in1), .out(andOp_245_out));

	wire [31:0] concat_246_in0;
	wire [31:0] concat_246_in1;
	wire [63:0] concat_246_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_246(.in0(concat_246_in0), .in1(concat_246_in1), .out(concat_246_out));

	wire [31:0] concat_247_in0;
	wire [31:0] concat_247_in1;
	wire [63:0] concat_247_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_247(.in0(concat_247_in0), .in1(concat_247_in1), .out(concat_247_out));

	wire [0:0] andOp_248_in0;
	wire [0:0] andOp_248_in1;
	wire [0:0] andOp_248_out;
	andOp #(.WIDTH(1)) andOp_248(.in0(andOp_248_in0), .in1(andOp_248_in1), .out(andOp_248_out));

	wire [0:0] andOp_249_in0;
	wire [0:0] andOp_249_in1;
	wire [0:0] andOp_249_out;
	andOp #(.WIDTH(1)) andOp_249(.in0(andOp_249_in0), .in1(andOp_249_in1), .out(andOp_249_out));

	reg [31:0] tmp_output_250_in_data;
	wire [31:0] tmp_output_250_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_250(.in_data(tmp_output_250_in_data), .out_data(tmp_output_250_out_data));

	wire [31:0] eq_251_in0;
	wire [31:0] eq_251_in1;
	wire [0:0] eq_251_out;
	eq #(.WIDTH(32)) eq_251(.in0(eq_251_in0), .in1(eq_251_in1), .out(eq_251_out));

	wire [31:0] eq_252_in0;
	wire [31:0] eq_252_in1;
	wire [0:0] eq_252_out;
	eq #(.WIDTH(32)) eq_252(.in0(eq_252_in0), .in1(eq_252_in1), .out(eq_252_out));

	wire [0:0] andOp_253_in0;
	wire [0:0] andOp_253_in1;
	wire [0:0] andOp_253_out;
	andOp #(.WIDTH(1)) andOp_253(.in0(andOp_253_in0), .in1(andOp_253_in1), .out(andOp_253_out));

	wire [0:0] andOp_254_in0;
	wire [0:0] andOp_254_in1;
	wire [0:0] andOp_254_out;
	andOp #(.WIDTH(1)) andOp_254(.in0(andOp_254_in0), .in1(andOp_254_in1), .out(andOp_254_out));

	wire [0:0] andOp_255_in0;
	wire [0:0] andOp_255_in1;
	wire [0:0] andOp_255_out;
	andOp #(.WIDTH(1)) andOp_255(.in0(andOp_255_in0), .in1(andOp_255_in1), .out(andOp_255_out));

	wire [0:0] andOp_256_in0;
	wire [0:0] andOp_256_in1;
	wire [0:0] andOp_256_out;
	andOp #(.WIDTH(1)) andOp_256(.in0(andOp_256_in0), .in1(andOp_256_in1), .out(andOp_256_out));

	reg [31:0] tmp_output_257_in_data;
	wire [31:0] tmp_output_257_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_257(.in_data(tmp_output_257_in_data), .out_data(tmp_output_257_out_data));

	wire [31:0] eq_258_in0;
	wire [31:0] eq_258_in1;
	wire [0:0] eq_258_out;
	eq #(.WIDTH(32)) eq_258(.in0(eq_258_in0), .in1(eq_258_in1), .out(eq_258_out));

	wire [31:0] eq_259_in0;
	wire [31:0] eq_259_in1;
	wire [0:0] eq_259_out;
	eq #(.WIDTH(32)) eq_259(.in0(eq_259_in0), .in1(eq_259_in1), .out(eq_259_out));

	wire [0:0] andOp_260_in0;
	wire [0:0] andOp_260_in1;
	wire [0:0] andOp_260_out;
	andOp #(.WIDTH(1)) andOp_260(.in0(andOp_260_in0), .in1(andOp_260_in1), .out(andOp_260_out));

	wire [0:0] andOp_261_in0;
	wire [0:0] andOp_261_in1;
	wire [0:0] andOp_261_out;
	andOp #(.WIDTH(1)) andOp_261(.in0(andOp_261_in0), .in1(andOp_261_in1), .out(andOp_261_out));

	wire [0:0] andOp_262_in0;
	wire [0:0] andOp_262_in1;
	wire [0:0] andOp_262_out;
	andOp #(.WIDTH(1)) andOp_262(.in0(andOp_262_in0), .in1(andOp_262_in1), .out(andOp_262_out));

	wire [0:0] andOp_263_in0;
	wire [0:0] andOp_263_in1;
	wire [0:0] andOp_263_out;
	andOp #(.WIDTH(1)) andOp_263(.in0(andOp_263_in0), .in1(andOp_263_in1), .out(andOp_263_out));

	wire [0:0] andOp_264_in0;
	wire [0:0] andOp_264_in1;
	wire [0:0] andOp_264_out;
	andOp #(.WIDTH(1)) andOp_264(.in0(andOp_264_in0), .in1(andOp_264_in1), .out(andOp_264_out));

	wire [0:0] andOp_265_in0;
	wire [0:0] andOp_265_in1;
	wire [0:0] andOp_265_out;
	andOp #(.WIDTH(1)) andOp_265(.in0(andOp_265_in0), .in1(andOp_265_in1), .out(andOp_265_out));

	wire [0:0] andOp_266_in0;
	wire [0:0] andOp_266_in1;
	wire [0:0] andOp_266_out;
	andOp #(.WIDTH(1)) andOp_266(.in0(andOp_266_in0), .in1(andOp_266_in1), .out(andOp_266_out));

	wire [0:0] andOp_267_in0;
	wire [0:0] andOp_267_in1;
	wire [0:0] andOp_267_out;
	andOp #(.WIDTH(1)) andOp_267(.in0(andOp_267_in0), .in1(andOp_267_in1), .out(andOp_267_out));

	wire [0:0] notOp_268_in0;
	wire [0:0] notOp_268_out;
	notOp #(.WIDTH(1)) notOp_268(.in(notOp_268_in0), .out(notOp_268_out));

	wire [0:0] andOp_269_in0;
	wire [0:0] andOp_269_in1;
	wire [0:0] andOp_269_out;
	andOp #(.WIDTH(1)) andOp_269(.in0(andOp_269_in0), .in1(andOp_269_in1), .out(andOp_269_out));

	wire [0:0] notOp_270_in0;
	wire [0:0] notOp_270_out;
	notOp #(.WIDTH(1)) notOp_270(.in(notOp_270_in0), .out(notOp_270_out));

	wire [0:0] andOp_271_in0;
	wire [0:0] andOp_271_in1;
	wire [0:0] andOp_271_out;
	andOp #(.WIDTH(1)) andOp_271(.in0(andOp_271_in0), .in1(andOp_271_in1), .out(andOp_271_out));

	wire [0:0] notOp_272_in0;
	wire [0:0] notOp_272_out;
	notOp #(.WIDTH(1)) notOp_272(.in(notOp_272_in0), .out(notOp_272_out));

	wire [0:0] andOp_273_in0;
	wire [0:0] andOp_273_in1;
	wire [0:0] andOp_273_out;
	andOp #(.WIDTH(1)) andOp_273(.in0(andOp_273_in0), .in1(andOp_273_in1), .out(andOp_273_out));

	wire [0:0] notOp_274_in0;
	wire [0:0] notOp_274_out;
	notOp #(.WIDTH(1)) notOp_274(.in(notOp_274_in0), .out(notOp_274_out));

	wire [0:0] andOp_275_in0;
	wire [0:0] andOp_275_in1;
	wire [0:0] andOp_275_out;
	andOp #(.WIDTH(1)) andOp_275(.in0(andOp_275_in0), .in1(andOp_275_in1), .out(andOp_275_out));

	wire [0:0] notOp_276_in0;
	wire [0:0] notOp_276_out;
	notOp #(.WIDTH(1)) notOp_276(.in(notOp_276_in0), .out(notOp_276_out));

	wire [0:0] andOp_277_in0;
	wire [0:0] andOp_277_in1;
	wire [0:0] andOp_277_out;
	andOp #(.WIDTH(1)) andOp_277(.in0(andOp_277_in0), .in1(andOp_277_in1), .out(andOp_277_out));

	wire [0:0] notOp_278_in0;
	wire [0:0] notOp_278_out;
	notOp #(.WIDTH(1)) notOp_278(.in(notOp_278_in0), .out(notOp_278_out));

	wire [0:0] andOp_279_in0;
	wire [0:0] andOp_279_in1;
	wire [0:0] andOp_279_out;
	andOp #(.WIDTH(1)) andOp_279(.in0(andOp_279_in0), .in1(andOp_279_in1), .out(andOp_279_out));

	wire [0:0] notOp_280_in0;
	wire [0:0] notOp_280_out;
	notOp #(.WIDTH(1)) notOp_280(.in(notOp_280_in0), .out(notOp_280_out));

	wire [0:0] andOp_281_in0;
	wire [0:0] andOp_281_in1;
	wire [0:0] andOp_281_out;
	andOp #(.WIDTH(1)) andOp_281(.in0(andOp_281_in0), .in1(andOp_281_in1), .out(andOp_281_out));

	wire [0:0] notOp_282_in0;
	wire [0:0] notOp_282_out;
	notOp #(.WIDTH(1)) notOp_282(.in(notOp_282_in0), .out(notOp_282_out));

	wire [0:0] andOp_283_in0;
	wire [0:0] andOp_283_in1;
	wire [0:0] andOp_283_out;
	andOp #(.WIDTH(1)) andOp_283(.in0(andOp_283_in0), .in1(andOp_283_in1), .out(andOp_283_out));

	wire [0:0] notOp_284_in0;
	wire [0:0] notOp_284_out;
	notOp #(.WIDTH(1)) notOp_284(.in(notOp_284_in0), .out(notOp_284_out));

	wire [0:0] andOp_285_in0;
	wire [0:0] andOp_285_in1;
	wire [0:0] andOp_285_out;
	andOp #(.WIDTH(1)) andOp_285(.in0(andOp_285_in0), .in1(andOp_285_in1), .out(andOp_285_out));

	wire [0:0] notOp_286_in0;
	wire [0:0] notOp_286_out;
	notOp #(.WIDTH(1)) notOp_286(.in(notOp_286_in0), .out(notOp_286_out));

	wire [0:0] andOp_287_in0;
	wire [0:0] andOp_287_in1;
	wire [0:0] andOp_287_out;
	andOp #(.WIDTH(1)) andOp_287(.in0(andOp_287_in0), .in1(andOp_287_in1), .out(andOp_287_out));

	wire [0:0] notOp_288_in0;
	wire [0:0] notOp_288_out;
	notOp #(.WIDTH(1)) notOp_288(.in(notOp_288_in0), .out(notOp_288_out));

	wire [0:0] andOp_289_in0;
	wire [0:0] andOp_289_in1;
	wire [0:0] andOp_289_out;
	andOp #(.WIDTH(1)) andOp_289(.in0(andOp_289_in0), .in1(andOp_289_in1), .out(andOp_289_out));

	wire [0:0] notOp_290_in0;
	wire [0:0] notOp_290_out;
	notOp #(.WIDTH(1)) notOp_290(.in(notOp_290_in0), .out(notOp_290_out));

	wire [0:0] andOp_291_in0;
	wire [0:0] andOp_291_in1;
	wire [0:0] andOp_291_out;
	andOp #(.WIDTH(1)) andOp_291(.in0(andOp_291_in0), .in1(andOp_291_in1), .out(andOp_291_out));

	wire [0:0] notOp_292_in0;
	wire [0:0] notOp_292_out;
	notOp #(.WIDTH(1)) notOp_292(.in(notOp_292_in0), .out(notOp_292_out));

	wire [0:0] andOp_293_in0;
	wire [0:0] andOp_293_in1;
	wire [0:0] andOp_293_out;
	andOp #(.WIDTH(1)) andOp_293(.in0(andOp_293_in0), .in1(andOp_293_in1), .out(andOp_293_out));

	wire [0:0] notOp_294_in0;
	wire [0:0] notOp_294_out;
	notOp #(.WIDTH(1)) notOp_294(.in(notOp_294_in0), .out(notOp_294_out));

	wire [0:0] andOp_295_in0;
	wire [0:0] andOp_295_in1;
	wire [0:0] andOp_295_out;
	andOp #(.WIDTH(1)) andOp_295(.in0(andOp_295_in0), .in1(andOp_295_in1), .out(andOp_295_out));

	wire [0:0] notOp_296_in0;
	wire [0:0] notOp_296_out;
	notOp #(.WIDTH(1)) notOp_296(.in(notOp_296_in0), .out(notOp_296_out));

	wire [0:0] andOp_297_in0;
	wire [0:0] andOp_297_in1;
	wire [0:0] andOp_297_out;
	andOp #(.WIDTH(1)) andOp_297(.in0(andOp_297_in0), .in1(andOp_297_in1), .out(andOp_297_out));

	wire [0:0] notOp_298_in0;
	wire [0:0] notOp_298_out;
	notOp #(.WIDTH(1)) notOp_298(.in(notOp_298_in0), .out(notOp_298_out));

	wire [0:0] andOp_299_in0;
	wire [0:0] andOp_299_in1;
	wire [0:0] andOp_299_out;
	andOp #(.WIDTH(1)) andOp_299(.in0(andOp_299_in0), .in1(andOp_299_in1), .out(andOp_299_out));

	wire [0:0] notOp_300_in0;
	wire [0:0] notOp_300_out;
	notOp #(.WIDTH(1)) notOp_300(.in(notOp_300_in0), .out(notOp_300_out));

	wire [0:0] andOp_301_in0;
	wire [0:0] andOp_301_in1;
	wire [0:0] andOp_301_out;
	andOp #(.WIDTH(1)) andOp_301(.in0(andOp_301_in0), .in1(andOp_301_in1), .out(andOp_301_out));

	wire [31:0] eq_302_in0;
	wire [31:0] eq_302_in1;
	wire [0:0] eq_302_out;
	eq #(.WIDTH(32)) eq_302(.in0(eq_302_in0), .in1(eq_302_in1), .out(eq_302_out));

	wire [31:0] eq_303_in0;
	wire [31:0] eq_303_in1;
	wire [0:0] eq_303_out;
	eq #(.WIDTH(32)) eq_303(.in0(eq_303_in0), .in1(eq_303_in1), .out(eq_303_out));

	wire [31:0] eq_304_in0;
	wire [31:0] eq_304_in1;
	wire [0:0] eq_304_out;
	eq #(.WIDTH(32)) eq_304(.in0(eq_304_in0), .in1(eq_304_in1), .out(eq_304_out));

	wire [31:0] eq_305_in0;
	wire [31:0] eq_305_in1;
	wire [0:0] eq_305_out;
	eq #(.WIDTH(32)) eq_305(.in0(eq_305_in0), .in1(eq_305_in1), .out(eq_305_out));

	wire [0:0] andOp_306_in0;
	wire [0:0] andOp_306_in1;
	wire [0:0] andOp_306_out;
	andOp #(.WIDTH(1)) andOp_306(.in0(andOp_306_in0), .in1(andOp_306_in1), .out(andOp_306_out));

	wire [31:0] eq_307_in0;
	wire [31:0] eq_307_in1;
	wire [0:0] eq_307_out;
	eq #(.WIDTH(32)) eq_307(.in0(eq_307_in0), .in1(eq_307_in1), .out(eq_307_out));

	wire [31:0] eq_308_in0;
	wire [31:0] eq_308_in1;
	wire [0:0] eq_308_out;
	eq #(.WIDTH(32)) eq_308(.in0(eq_308_in0), .in1(eq_308_in1), .out(eq_308_out));

	wire [31:0] eq_309_in0;
	wire [31:0] eq_309_in1;
	wire [0:0] eq_309_out;
	eq #(.WIDTH(32)) eq_309(.in0(eq_309_in0), .in1(eq_309_in1), .out(eq_309_out));

	wire [31:0] eq_310_in0;
	wire [31:0] eq_310_in1;
	wire [0:0] eq_310_out;
	eq #(.WIDTH(32)) eq_310(.in0(eq_310_in0), .in1(eq_310_in1), .out(eq_310_out));

	wire [0:0] andOp_311_in0;
	wire [0:0] andOp_311_in1;
	wire [0:0] andOp_311_out;
	andOp #(.WIDTH(1)) andOp_311(.in0(andOp_311_in0), .in1(andOp_311_in1), .out(andOp_311_out));

	wire [31:0] eq_312_in0;
	wire [31:0] eq_312_in1;
	wire [0:0] eq_312_out;
	eq #(.WIDTH(32)) eq_312(.in0(eq_312_in0), .in1(eq_312_in1), .out(eq_312_out));

	wire [31:0] eq_313_in0;
	wire [31:0] eq_313_in1;
	wire [0:0] eq_313_out;
	eq #(.WIDTH(32)) eq_313(.in0(eq_313_in0), .in1(eq_313_in1), .out(eq_313_out));

	wire [31:0] eq_314_in0;
	wire [31:0] eq_314_in1;
	wire [0:0] eq_314_out;
	eq #(.WIDTH(32)) eq_314(.in0(eq_314_in0), .in1(eq_314_in1), .out(eq_314_out));

	wire [31:0] eq_315_in0;
	wire [31:0] eq_315_in1;
	wire [0:0] eq_315_out;
	eq #(.WIDTH(32)) eq_315(.in0(eq_315_in0), .in1(eq_315_in1), .out(eq_315_out));

	wire [0:0] andOp_316_in0;
	wire [0:0] andOp_316_in1;
	wire [0:0] andOp_316_out;
	andOp #(.WIDTH(1)) andOp_316(.in0(andOp_316_in0), .in1(andOp_316_in1), .out(andOp_316_out));

	wire [31:0] eq_317_in0;
	wire [31:0] eq_317_in1;
	wire [0:0] eq_317_out;
	eq #(.WIDTH(32)) eq_317(.in0(eq_317_in0), .in1(eq_317_in1), .out(eq_317_out));

	wire [31:0] eq_318_in0;
	wire [31:0] eq_318_in1;
	wire [0:0] eq_318_out;
	eq #(.WIDTH(32)) eq_318(.in0(eq_318_in0), .in1(eq_318_in1), .out(eq_318_out));

	wire [31:0] eq_319_in0;
	wire [31:0] eq_319_in1;
	wire [0:0] eq_319_out;
	eq #(.WIDTH(32)) eq_319(.in0(eq_319_in0), .in1(eq_319_in1), .out(eq_319_out));

	wire [0:0] andOp_320_in0;
	wire [0:0] andOp_320_in1;
	wire [0:0] andOp_320_out;
	andOp #(.WIDTH(1)) andOp_320(.in0(andOp_320_in0), .in1(andOp_320_in1), .out(andOp_320_out));

	wire [31:0] eq_321_in0;
	wire [31:0] eq_321_in1;
	wire [0:0] eq_321_out;
	eq #(.WIDTH(32)) eq_321(.in0(eq_321_in0), .in1(eq_321_in1), .out(eq_321_out));

	wire [31:0] eq_322_in0;
	wire [31:0] eq_322_in1;
	wire [0:0] eq_322_out;
	eq #(.WIDTH(32)) eq_322(.in0(eq_322_in0), .in1(eq_322_in1), .out(eq_322_out));

	wire [31:0] eq_323_in0;
	wire [31:0] eq_323_in1;
	wire [0:0] eq_323_out;
	eq #(.WIDTH(32)) eq_323(.in0(eq_323_in0), .in1(eq_323_in1), .out(eq_323_out));

	wire [31:0] eq_324_in0;
	wire [31:0] eq_324_in1;
	wire [0:0] eq_324_out;
	eq #(.WIDTH(32)) eq_324(.in0(eq_324_in0), .in1(eq_324_in1), .out(eq_324_out));

	wire [0:0] andOp_325_in0;
	wire [0:0] andOp_325_in1;
	wire [0:0] andOp_325_out;
	andOp #(.WIDTH(1)) andOp_325(.in0(andOp_325_in0), .in1(andOp_325_in1), .out(andOp_325_out));

	wire [31:0] eq_326_in0;
	wire [31:0] eq_326_in1;
	wire [0:0] eq_326_out;
	eq #(.WIDTH(32)) eq_326(.in0(eq_326_in0), .in1(eq_326_in1), .out(eq_326_out));

	wire [31:0] eq_327_in0;
	wire [31:0] eq_327_in1;
	wire [0:0] eq_327_out;
	eq #(.WIDTH(32)) eq_327(.in0(eq_327_in0), .in1(eq_327_in1), .out(eq_327_out));

	// End Functional Units

	reg [31:0] data_store_1_0;
	reg [31:0] data_store_1_2;
	reg [31:0] data_store_1_4;
	reg [31:0] data_store_2_10;
	reg [31:0] data_store_2_6;
	reg [31:0] data_store_2_8;
	reg [31:0] data_store_3_12;
	reg [31:0] data_store_3_14;
	reg [31:0] data_store_3_16;
	reg [31:0] data_store_4_18;
	reg [31:0] data_store_4_20;
	reg [31:0] data_store_4_22;
	reg [31:0] data_store_5_24;
	reg [31:0] data_store_5_26;
	reg [31:0] data_store_5_28;
	reg [31:0] data_store_6_30;
	reg [31:0] data_store_6_32;
	reg [31:0] data_store_7_34;
	reg [31:0] data_store_7_36;
	reg [31:0] data_store_8_38;
	reg [31:0] data_store_8_40;
	reg [31:0] global_state;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_3_last_state;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;
	reg [31:0] state_4_last_state;
	reg [31:0] state_5_entry_BB_reg;
	reg [0:0] state_5_is_active;
	reg [31:0] state_5_last_BB_reg;
	reg [31:0] state_5_last_state;
	reg [31:0] state_6_entry_BB_reg;
	reg [0:0] state_6_is_active;
	reg [31:0] state_6_last_BB_reg;
	reg [31:0] state_6_last_state;
	reg [31:0] state_7_entry_BB_reg;
	reg [0:0] state_7_is_active;
	reg [31:0] state_7_last_BB_reg;
	reg [31:0] state_7_last_state;
	reg [31:0] state_8_entry_BB_reg;
	reg [0:0] state_8_is_active;
	reg [31:0] state_8_last_BB_reg;
	reg [31:0] state_8_last_state;
	reg [31:0] state_9_entry_BB_reg;
	reg [0:0] state_9_is_active;
	reg [31:0] state_9_last_BB_reg;
	reg [31:0] state_9_last_state;

	// controller for _____dlr_0___eq___alloca___dlr_builtin_fifo_32._____dlr_0___eq___alloca___dlr_builtin_fifo_32_in_data
	always @(*) begin
		if (andOp_223_out) begin 
			_____dlr_0___eq___alloca___dlr_builtin_fifo_32_in_data = tmp_output_224_out_data;
		end else begin
			_____dlr_0___eq___alloca___dlr_builtin_fifo_32_in_data = 0;
		end
	end
	// controller for _____dlr_0___eq___alloca___dlr_builtin_fifo_32._____dlr_0___eq___alloca___dlr_builtin_fifo_32_read_valid
	always @(*) begin
		if (andOp_228_out) begin 
			_____dlr_0___eq___alloca___dlr_builtin_fifo_32_read_valid = -(1'd1);
		end else begin
			_____dlr_0___eq___alloca___dlr_builtin_fifo_32_read_valid = 0;
		end
	end
	// controller for _____dlr_0___eq___alloca___dlr_builtin_fifo_32._____dlr_0___eq___alloca___dlr_builtin_fifo_32_write_valid
	always @(*) begin
		if (andOp_222_out) begin 
			_____dlr_0___eq___alloca___dlr_builtin_fifo_32_write_valid = -(1'd1);
		end else begin
			_____dlr_0___eq___alloca___dlr_builtin_fifo_32_write_valid = 0;
		end
	end
	// controller for add_add26.add_add26_in0
	// controller for add_add26.add_add26_in1
	// Insensitive connections
	assign add_add26_in0 = data_in_5_27_out_data;
	assign add_add26_in1 = tmp_output_242_out_data;
	// controller for add_add29.add_add29_in0
	// controller for add_add29.add_add29_in1
	// Insensitive connections
	assign add_add29_in0 = phi_phi28_out;
	assign add_add29_in1 = 32'd1;
	// controller for add_add5.add_add5_in0
	// controller for add_add5.add_add5_in1
	// Insensitive connections
	assign add_add5_in0 = phi_phi3_out;
	assign add_add5_in1 = 32'd1;
	// controller for andOp_101.andOp_101_in0
	// controller for andOp_101.andOp_101_in1
	// Insensitive connections
	assign andOp_101_in0 = andOp_97_out;
	assign andOp_101_in1 = notOp_100_out;
	// controller for andOp_102.andOp_102_in0
	// controller for andOp_102.andOp_102_in1
	// Insensitive connections
	assign andOp_102_in0 = bb_14_active_in_state_8_out_data;
	assign andOp_102_in1 = state_8_is_active;
	// controller for andOp_104.andOp_104_in0
	// controller for andOp_104.andOp_104_in1
	// Insensitive connections
	assign andOp_104_in0 = bb_2_active_in_state_8_out_data;
	assign andOp_104_in1 = state_8_is_active;
	// controller for andOp_106.andOp_106_in0
	// controller for andOp_106.andOp_106_in1
	// Insensitive connections
	assign andOp_106_in0 = bb_11_active_in_state_8_out_data;
	assign andOp_106_in1 = state_8_is_active;
	// controller for andOp_108.andOp_108_in0
	// controller for andOp_108.andOp_108_in1
	// Insensitive connections
	assign andOp_108_in0 = bb_3_active_in_state_8_out_data;
	assign andOp_108_in1 = state_8_is_active;
	// controller for andOp_110.andOp_110_in0
	// controller for andOp_110.andOp_110_in1
	// Insensitive connections
	assign andOp_110_in0 = andOp_108_out;
	assign andOp_110_in1 = icmp_icmp37_out;
	// controller for andOp_112.andOp_112_in0
	// controller for andOp_112.andOp_112_in1
	// Insensitive connections
	assign andOp_112_in0 = andOp_108_out;
	assign andOp_112_in1 = notOp_111_out;
	// controller for andOp_113.andOp_113_in0
	// controller for andOp_113.andOp_113_in1
	// Insensitive connections
	assign andOp_113_in0 = bb_12_active_in_state_8_out_data;
	assign andOp_113_in1 = state_8_is_active;
	// controller for andOp_162.andOp_162_in0
	// controller for andOp_162.andOp_162_in1
	// Insensitive connections
	assign andOp_162_in0 = notOp_161_out;
	assign andOp_162_in1 = andOp_46_out;
	// controller for andOp_166.andOp_166_in0
	// controller for andOp_166.andOp_166_in1
	// Insensitive connections
	assign andOp_166_in0 = notOp_165_out;
	assign andOp_166_in1 = andOp_44_out;
	// controller for andOp_171.andOp_171_in0
	// controller for andOp_171.andOp_171_in1
	// Insensitive connections
	assign andOp_171_in0 = notOp_170_out;
	assign andOp_171_in1 = andOp_64_out;
	// controller for andOp_174.andOp_174_in0
	// controller for andOp_174.andOp_174_in1
	// Insensitive connections
	assign andOp_174_in0 = notOp_173_out;
	assign andOp_174_in1 = andOp_57_out;
	// controller for andOp_177.andOp_177_in0
	// controller for andOp_177.andOp_177_in1
	// Insensitive connections
	assign andOp_177_in0 = notOp_176_out;
	assign andOp_177_in1 = andOp_53_out;
	// controller for andOp_181.andOp_181_in0
	// controller for andOp_181.andOp_181_in1
	// Insensitive connections
	assign andOp_181_in0 = notOp_180_out;
	assign andOp_181_in1 = andOp_80_out;
	// controller for andOp_184.andOp_184_in0
	// controller for andOp_184.andOp_184_in1
	// Insensitive connections
	assign andOp_184_in0 = notOp_183_out;
	assign andOp_184_in1 = andOp_70_out;
	// controller for andOp_187.andOp_187_in0
	// controller for andOp_187.andOp_187_in1
	// Insensitive connections
	assign andOp_187_in0 = notOp_186_out;
	assign andOp_187_in1 = andOp_73_out;
	// controller for andOp_190.andOp_190_in0
	// controller for andOp_190.andOp_190_in1
	// Insensitive connections
	assign andOp_190_in0 = notOp_189_out;
	assign andOp_190_in1 = andOp_84_out;
	// controller for andOp_194.andOp_194_in0
	// controller for andOp_194.andOp_194_in1
	// Insensitive connections
	assign andOp_194_in0 = notOp_193_out;
	assign andOp_194_in1 = andOp_66_out;
	// controller for andOp_197.andOp_197_in0
	// controller for andOp_197.andOp_197_in1
	// Insensitive connections
	assign andOp_197_in0 = notOp_196_out;
	assign andOp_197_in1 = andOp_88_out;
	// controller for andOp_201.andOp_201_in0
	// controller for andOp_201.andOp_201_in1
	// Insensitive connections
	assign andOp_201_in0 = notOp_200_out;
	assign andOp_201_in1 = andOp_86_out;
	// controller for andOp_205.andOp_205_in0
	// controller for andOp_205.andOp_205_in1
	// Insensitive connections
	assign andOp_205_in0 = notOp_204_out;
	assign andOp_205_in1 = andOp_113_out;
	// controller for andOp_208.andOp_208_in0
	// controller for andOp_208.andOp_208_in1
	// Insensitive connections
	assign andOp_208_in0 = notOp_207_out;
	assign andOp_208_in1 = andOp_99_out;
	// controller for andOp_211.andOp_211_in0
	// controller for andOp_211.andOp_211_in1
	// Insensitive connections
	assign andOp_211_in0 = notOp_210_out;
	assign andOp_211_in1 = andOp_95_out;
	// controller for andOp_215.andOp_215_in0
	// controller for andOp_215.andOp_215_in1
	// Insensitive connections
	assign andOp_215_in0 = notOp_214_out;
	assign andOp_215_in1 = andOp_102_out;
	// controller for andOp_218.andOp_218_in0
	// controller for andOp_218.andOp_218_in1
	// Insensitive connections
	assign andOp_218_in0 = notOp_217_out;
	assign andOp_218_in1 = andOp_104_out;
	// controller for andOp_220.andOp_220_in0
	// controller for andOp_220.andOp_220_in1
	// Insensitive connections
	assign andOp_220_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_220_in1 = state_0_is_active;
	// controller for andOp_221.andOp_221_in0
	// controller for andOp_221.andOp_221_in1
	// Insensitive connections
	assign andOp_221_in0 = bb_22_active_in_state_5_out_data;
	assign andOp_221_in1 = state_5_is_active;
	// controller for andOp_222.andOp_222_in0
	// controller for andOp_222.andOp_222_in1
	// Insensitive connections
	assign andOp_222_in0 = bb_23_active_in_state_5_out_data;
	assign andOp_222_in1 = state_5_is_active;
	// controller for andOp_223.andOp_223_in0
	// controller for andOp_223.andOp_223_in1
	// Insensitive connections
	assign andOp_223_in0 = bb_23_active_in_state_5_out_data;
	assign andOp_223_in1 = state_5_is_active;
	// controller for andOp_227.andOp_227_in0
	// controller for andOp_227.andOp_227_in1
	// Insensitive connections
	assign andOp_227_in0 = bb_10_active_in_state_6_out_data;
	assign andOp_227_in1 = state_6_is_active;
	// controller for andOp_228.andOp_228_in0
	// controller for andOp_228.andOp_228_in1
	// Insensitive connections
	assign andOp_228_in0 = bb_11_active_in_state_7_out_data;
	assign andOp_228_in1 = state_7_is_active;
	// controller for andOp_229.andOp_229_in0
	// controller for andOp_229.andOp_229_in1
	// Insensitive connections
	assign andOp_229_in0 = bb_11_active_in_state_8_out_data;
	assign andOp_229_in1 = state_8_is_active;
	// controller for andOp_230.andOp_230_in0
	// controller for andOp_230.andOp_230_in1
	// Insensitive connections
	assign andOp_230_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_230_in1 = state_1_is_active;
	// controller for andOp_233.andOp_233_in0
	// controller for andOp_233.andOp_233_in1
	// Insensitive connections
	assign andOp_233_in0 = bb_16_active_in_state_1_out_data;
	assign andOp_233_in1 = state_1_is_active;
	// controller for andOp_234.andOp_234_in0
	// controller for andOp_234.andOp_234_in1
	// Insensitive connections
	assign andOp_234_in0 = bb_17_active_in_state_2_out_data;
	assign andOp_234_in1 = state_2_is_active;
	// controller for andOp_235.andOp_235_in0
	// controller for andOp_235.andOp_235_in1
	// Insensitive connections
	assign andOp_235_in0 = bb_17_active_in_state_3_out_data;
	assign andOp_235_in1 = state_3_is_active;
	// controller for andOp_236.andOp_236_in0
	// controller for andOp_236.andOp_236_in1
	// Insensitive connections
	assign andOp_236_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_236_in1 = state_1_is_active;
	// controller for andOp_237.andOp_237_in0
	// controller for andOp_237.andOp_237_in1
	// Insensitive connections
	assign andOp_237_in0 = bb_19_active_in_state_3_out_data;
	assign andOp_237_in1 = state_3_is_active;
	// controller for andOp_238.andOp_238_in0
	// controller for andOp_238.andOp_238_in1
	// Insensitive connections
	assign andOp_238_in0 = bb_20_active_in_state_4_out_data;
	assign andOp_238_in1 = state_4_is_active;
	// controller for andOp_239.andOp_239_in0
	// controller for andOp_239.andOp_239_in1
	// Insensitive connections
	assign andOp_239_in0 = bb_20_active_in_state_5_out_data;
	assign andOp_239_in1 = state_5_is_active;
	// controller for andOp_240.andOp_240_in0
	// controller for andOp_240.andOp_240_in1
	// Insensitive connections
	assign andOp_240_in0 = bb_7_active_in_state_5_out_data;
	assign andOp_240_in1 = state_5_is_active;
	// controller for andOp_241.andOp_241_in0
	// controller for andOp_241.andOp_241_in1
	// Insensitive connections
	assign andOp_241_in0 = bb_6_active_in_state_5_out_data;
	assign andOp_241_in1 = state_5_is_active;
	// controller for andOp_245.andOp_245_in0
	// controller for andOp_245.andOp_245_in1
	// Insensitive connections
	assign andOp_245_in0 = bb_1_active_in_state_6_out_data;
	assign andOp_245_in1 = state_6_is_active;
	// controller for andOp_248.andOp_248_in0
	// controller for andOp_248.andOp_248_in1
	// Insensitive connections
	assign andOp_248_in0 = bb_1_active_in_state_6_out_data;
	assign andOp_248_in1 = state_6_is_active;
	// controller for andOp_249.andOp_249_in0
	// controller for andOp_249.andOp_249_in1
	// Insensitive connections
	assign andOp_249_in0 = bb_14_active_in_state_8_out_data;
	assign andOp_249_in1 = state_8_is_active;
	// controller for andOp_253.andOp_253_in0
	// controller for andOp_253.andOp_253_in1
	// Insensitive connections
	assign andOp_253_in0 = bb_14_active_in_state_8_out_data;
	assign andOp_253_in1 = state_8_is_active;
	// controller for andOp_254.andOp_254_in0
	// controller for andOp_254.andOp_254_in1
	// Insensitive connections
	assign andOp_254_in0 = bb_13_active_in_state_8_out_data;
	assign andOp_254_in1 = state_8_is_active;
	// controller for andOp_255.andOp_255_in0
	// controller for andOp_255.andOp_255_in1
	// Insensitive connections
	assign andOp_255_in0 = bb_3_active_in_state_8_out_data;
	assign andOp_255_in1 = state_8_is_active;
	// controller for andOp_256.andOp_256_in0
	// controller for andOp_256.andOp_256_in1
	// Insensitive connections
	assign andOp_256_in0 = bb_2_active_in_state_8_out_data;
	assign andOp_256_in1 = state_8_is_active;
	// controller for andOp_260.andOp_260_in0
	// controller for andOp_260.andOp_260_in1
	// Insensitive connections
	assign andOp_260_in0 = bb_8_active_in_state_9_out_data;
	assign andOp_260_in1 = state_9_is_active;
	// controller for andOp_261.andOp_261_in0
	// controller for andOp_261.andOp_261_in1
	// Insensitive connections
	assign andOp_261_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_261_in1 = state_0_is_active;
	// controller for andOp_262.andOp_262_in0
	// controller for andOp_262.andOp_262_in1
	// Insensitive connections
	assign andOp_262_in0 = bb_17_active_in_state_2_out_data;
	assign andOp_262_in1 = state_2_is_active;
	// controller for andOp_263.andOp_263_in0
	// controller for andOp_263.andOp_263_in1
	// Insensitive connections
	assign andOp_263_in0 = bb_20_active_in_state_4_out_data;
	assign andOp_263_in1 = state_4_is_active;
	// controller for andOp_264.andOp_264_in0
	// controller for andOp_264.andOp_264_in1
	// Insensitive connections
	assign andOp_264_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_264_in1 = state_0_is_active;
	// controller for andOp_265.andOp_265_in0
	// controller for andOp_265.andOp_265_in1
	// Insensitive connections
	assign andOp_265_in0 = bb_11_active_in_state_7_out_data;
	assign andOp_265_in1 = state_7_is_active;
	// controller for andOp_266.andOp_266_in0
	// controller for andOp_266.andOp_266_in1
	// Insensitive connections
	assign andOp_266_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_266_in1 = state_0_is_active;
	// controller for andOp_267.andOp_267_in0
	// controller for andOp_267.andOp_267_in1
	// Insensitive connections
	assign andOp_267_in0 = bb_8_active_in_state_9_out_data;
	assign andOp_267_in1 = state_9_is_active;
	// controller for andOp_269.andOp_269_in0
	// controller for andOp_269.andOp_269_in1
	// Insensitive connections
	assign andOp_269_in0 = notOp_268_out;
	assign andOp_269_in1 = 1'd1;
	// controller for andOp_271.andOp_271_in0
	// controller for andOp_271.andOp_271_in1
	// Insensitive connections
	assign andOp_271_in0 = notOp_270_out;
	assign andOp_271_in1 = andOp_269_out;
	// controller for andOp_273.andOp_273_in0
	// controller for andOp_273.andOp_273_in1
	// Insensitive connections
	assign andOp_273_in0 = notOp_272_out;
	assign andOp_273_in1 = andOp_271_out;
	// controller for andOp_275.andOp_275_in0
	// controller for andOp_275.andOp_275_in1
	// Insensitive connections
	assign andOp_275_in0 = notOp_274_out;
	assign andOp_275_in1 = 1'd1;
	// controller for andOp_277.andOp_277_in0
	// controller for andOp_277.andOp_277_in1
	// Insensitive connections
	assign andOp_277_in0 = notOp_276_out;
	assign andOp_277_in1 = 1'd1;
	// controller for andOp_279.andOp_279_in0
	// controller for andOp_279.andOp_279_in1
	// Insensitive connections
	assign andOp_279_in0 = notOp_278_out;
	assign andOp_279_in1 = andOp_277_out;
	// controller for andOp_281.andOp_281_in0
	// controller for andOp_281.andOp_281_in1
	// Insensitive connections
	assign andOp_281_in0 = notOp_280_out;
	assign andOp_281_in1 = 1'd1;
	// controller for andOp_283.andOp_283_in0
	// controller for andOp_283.andOp_283_in1
	// Insensitive connections
	assign andOp_283_in0 = notOp_282_out;
	assign andOp_283_in1 = 1'd1;
	// controller for andOp_285.andOp_285_in0
	// controller for andOp_285.andOp_285_in1
	// Insensitive connections
	assign andOp_285_in0 = notOp_284_out;
	assign andOp_285_in1 = andOp_283_out;
	// controller for andOp_287.andOp_287_in0
	// controller for andOp_287.andOp_287_in1
	// Insensitive connections
	assign andOp_287_in0 = notOp_286_out;
	assign andOp_287_in1 = 1'd1;
	// controller for andOp_289.andOp_289_in0
	// controller for andOp_289.andOp_289_in1
	// Insensitive connections
	assign andOp_289_in0 = notOp_288_out;
	assign andOp_289_in1 = andOp_287_out;
	// controller for andOp_291.andOp_291_in0
	// controller for andOp_291.andOp_291_in1
	// Insensitive connections
	assign andOp_291_in0 = notOp_290_out;
	assign andOp_291_in1 = andOp_289_out;
	// controller for andOp_293.andOp_293_in0
	// controller for andOp_293.andOp_293_in1
	// Insensitive connections
	assign andOp_293_in0 = notOp_292_out;
	assign andOp_293_in1 = 1'd1;
	// controller for andOp_295.andOp_295_in0
	// controller for andOp_295.andOp_295_in1
	// Insensitive connections
	assign andOp_295_in0 = notOp_294_out;
	assign andOp_295_in1 = 1'd1;
	// controller for andOp_297.andOp_297_in0
	// controller for andOp_297.andOp_297_in1
	// Insensitive connections
	assign andOp_297_in0 = notOp_296_out;
	assign andOp_297_in1 = andOp_295_out;
	// controller for andOp_299.andOp_299_in0
	// controller for andOp_299.andOp_299_in1
	// Insensitive connections
	assign andOp_299_in0 = notOp_298_out;
	assign andOp_299_in1 = 1'd1;
	// controller for andOp_301.andOp_301_in0
	// controller for andOp_301.andOp_301_in1
	// Insensitive connections
	assign andOp_301_in0 = notOp_300_out;
	assign andOp_301_in1 = andOp_299_out;
	// controller for andOp_306.andOp_306_in0
	// controller for andOp_306.andOp_306_in1
	// Insensitive connections
	assign andOp_306_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_306_in1 = state_1_is_active;
	// controller for andOp_311.andOp_311_in0
	// controller for andOp_311.andOp_311_in1
	// Insensitive connections
	assign andOp_311_in0 = bb_17_active_in_state_3_out_data;
	assign andOp_311_in1 = state_3_is_active;
	// controller for andOp_316.andOp_316_in0
	// controller for andOp_316.andOp_316_in1
	// Insensitive connections
	assign andOp_316_in0 = bb_6_active_in_state_5_out_data;
	assign andOp_316_in1 = state_5_is_active;
	// controller for andOp_320.andOp_320_in0
	// controller for andOp_320.andOp_320_in1
	// Insensitive connections
	assign andOp_320_in0 = bb_1_active_in_state_6_out_data;
	assign andOp_320_in1 = state_6_is_active;
	// controller for andOp_325.andOp_325_in0
	// controller for andOp_325.andOp_325_in1
	// Insensitive connections
	assign andOp_325_in0 = bb_2_active_in_state_8_out_data;
	assign andOp_325_in1 = state_8_is_active;
	// controller for andOp_42.andOp_42_in0
	// controller for andOp_42.andOp_42_in1
	// Insensitive connections
	assign andOp_42_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_42_in1 = state_0_is_active;
	// controller for andOp_44.andOp_44_in0
	// controller for andOp_44.andOp_44_in1
	// Insensitive connections
	assign andOp_44_in0 = bb_15_active_in_state_1_out_data;
	assign andOp_44_in1 = state_1_is_active;
	// controller for andOp_46.andOp_46_in0
	// controller for andOp_46.andOp_46_in1
	// Insensitive connections
	assign andOp_46_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_46_in1 = state_1_is_active;
	// controller for andOp_48.andOp_48_in0
	// controller for andOp_48.andOp_48_in1
	// Insensitive connections
	assign andOp_48_in0 = bb_16_active_in_state_1_out_data;
	assign andOp_48_in1 = state_1_is_active;
	// controller for andOp_50.andOp_50_in0
	// controller for andOp_50.andOp_50_in1
	// Insensitive connections
	assign andOp_50_in0 = andOp_48_out;
	assign andOp_50_in1 = arg_0_read_ready;
	// controller for andOp_52.andOp_52_in0
	// controller for andOp_52.andOp_52_in1
	// Insensitive connections
	assign andOp_52_in0 = andOp_48_out;
	assign andOp_52_in1 = notOp_51_out;
	// controller for andOp_53.andOp_53_in0
	// controller for andOp_53.andOp_53_in1
	// Insensitive connections
	assign andOp_53_in0 = bb_17_active_in_state_3_out_data;
	assign andOp_53_in1 = state_3_is_active;
	// controller for andOp_55.andOp_55_in0
	// controller for andOp_55.andOp_55_in1
	// Insensitive connections
	assign andOp_55_in0 = bb_17_active_in_state_3_out_data;
	assign andOp_55_in1 = state_3_is_active;
	// controller for andOp_57.andOp_57_in0
	// controller for andOp_57.andOp_57_in1
	// Insensitive connections
	assign andOp_57_in0 = bb_18_active_in_state_3_out_data;
	assign andOp_57_in1 = state_3_is_active;
	// controller for andOp_59.andOp_59_in0
	// controller for andOp_59.andOp_59_in1
	// Insensitive connections
	assign andOp_59_in0 = bb_19_active_in_state_3_out_data;
	assign andOp_59_in1 = state_3_is_active;
	// controller for andOp_61.andOp_61_in0
	// controller for andOp_61.andOp_61_in1
	// Insensitive connections
	assign andOp_61_in0 = andOp_59_out;
	assign andOp_61_in1 = arg_1_read_ready;
	// controller for andOp_63.andOp_63_in0
	// controller for andOp_63.andOp_63_in1
	// Insensitive connections
	assign andOp_63_in0 = andOp_59_out;
	assign andOp_63_in1 = notOp_62_out;
	// controller for andOp_64.andOp_64_in0
	// controller for andOp_64.andOp_64_in1
	// Insensitive connections
	assign andOp_64_in0 = bb_5_active_in_state_3_out_data;
	assign andOp_64_in1 = state_3_is_active;
	// controller for andOp_66.andOp_66_in0
	// controller for andOp_66.andOp_66_in1
	// Insensitive connections
	assign andOp_66_in0 = bb_20_active_in_state_5_out_data;
	assign andOp_66_in1 = state_5_is_active;
	// controller for andOp_68.andOp_68_in0
	// controller for andOp_68.andOp_68_in1
	// Insensitive connections
	assign andOp_68_in0 = bb_22_active_in_state_5_out_data;
	assign andOp_68_in1 = state_5_is_active;
	// controller for andOp_70.andOp_70_in0
	// controller for andOp_70.andOp_70_in1
	// Insensitive connections
	assign andOp_70_in0 = andOp_68_out;
	assign andOp_70_in1 = _____dlr_0___eq___alloca___dlr_builtin_fifo_32_write_ready;
	// controller for andOp_72.andOp_72_in0
	// controller for andOp_72.andOp_72_in1
	// Insensitive connections
	assign andOp_72_in0 = andOp_68_out;
	assign andOp_72_in1 = notOp_71_out;
	// controller for andOp_73.andOp_73_in0
	// controller for andOp_73.andOp_73_in1
	// Insensitive connections
	assign andOp_73_in0 = bb_23_active_in_state_5_out_data;
	assign andOp_73_in1 = state_5_is_active;
	// controller for andOp_75.andOp_75_in0
	// controller for andOp_75.andOp_75_in1
	// Insensitive connections
	assign andOp_75_in0 = bb_7_active_in_state_5_out_data;
	assign andOp_75_in1 = state_5_is_active;
	// controller for andOp_77.andOp_77_in0
	// controller for andOp_77.andOp_77_in1
	// Insensitive connections
	assign andOp_77_in0 = andOp_75_out;
	assign andOp_77_in1 = icmp_icmp16_out;
	// controller for andOp_79.andOp_79_in0
	// controller for andOp_79.andOp_79_in1
	// Insensitive connections
	assign andOp_79_in0 = andOp_75_out;
	assign andOp_79_in1 = notOp_78_out;
	// controller for andOp_80.andOp_80_in0
	// controller for andOp_80.andOp_80_in1
	// Insensitive connections
	assign andOp_80_in0 = bb_21_active_in_state_5_out_data;
	assign andOp_80_in1 = state_5_is_active;
	// controller for andOp_82.andOp_82_in0
	// controller for andOp_82.andOp_82_in1
	// Insensitive connections
	assign andOp_82_in0 = bb_20_active_in_state_5_out_data;
	assign andOp_82_in1 = state_5_is_active;
	// controller for andOp_84.andOp_84_in0
	// controller for andOp_84.andOp_84_in1
	// Insensitive connections
	assign andOp_84_in0 = bb_6_active_in_state_5_out_data;
	assign andOp_84_in1 = state_5_is_active;
	// controller for andOp_86.andOp_86_in0
	// controller for andOp_86.andOp_86_in1
	// Insensitive connections
	assign andOp_86_in0 = bb_9_active_in_state_6_out_data;
	assign andOp_86_in1 = state_6_is_active;
	// controller for andOp_88.andOp_88_in0
	// controller for andOp_88.andOp_88_in1
	// Insensitive connections
	assign andOp_88_in0 = bb_1_active_in_state_6_out_data;
	assign andOp_88_in1 = state_6_is_active;
	// controller for andOp_90.andOp_90_in0
	// controller for andOp_90.andOp_90_in1
	// Insensitive connections
	assign andOp_90_in0 = bb_10_active_in_state_6_out_data;
	assign andOp_90_in1 = state_6_is_active;
	// controller for andOp_92.andOp_92_in0
	// controller for andOp_92.andOp_92_in1
	// Insensitive connections
	assign andOp_92_in0 = andOp_90_out;
	assign andOp_92_in1 = _____dlr_0___eq___alloca___dlr_builtin_fifo_32_read_ready;
	// controller for andOp_94.andOp_94_in0
	// controller for andOp_94.andOp_94_in1
	// Insensitive connections
	assign andOp_94_in0 = andOp_90_out;
	assign andOp_94_in1 = notOp_93_out;
	// controller for andOp_95.andOp_95_in0
	// controller for andOp_95.andOp_95_in1
	// Insensitive connections
	assign andOp_95_in0 = bb_11_active_in_state_8_out_data;
	assign andOp_95_in1 = state_8_is_active;
	// controller for andOp_97.andOp_97_in0
	// controller for andOp_97.andOp_97_in1
	// Insensitive connections
	assign andOp_97_in0 = bb_13_active_in_state_8_out_data;
	assign andOp_97_in1 = state_8_is_active;
	// controller for andOp_99.andOp_99_in0
	// controller for andOp_99.andOp_99_in1
	// Insensitive connections
	assign andOp_99_in0 = andOp_97_out;
	assign andOp_99_in1 = arg_2_write_ready;
	// controller for arg_0.arg_0_read_valid_reg
	always @(*) begin
		if (andOp_234_out) begin 
			arg_0_read_valid_reg = -(1'd1);
		end else begin
			arg_0_read_valid_reg = 0;
		end
	end
	// controller for arg_1.arg_1_read_valid_reg
	always @(*) begin
		if (andOp_238_out) begin 
			arg_1_read_valid_reg = -(1'd1);
		end else begin
			arg_1_read_valid_reg = 0;
		end
	end
	// controller for arg_2.arg_2_in_data_reg
	always @(*) begin
		if (andOp_249_out) begin 
			arg_2_in_data_reg = tmp_output_250_out_data;
		end else begin
			arg_2_in_data_reg = 0;
		end
	end
	// controller for arg_2.arg_2_write_valid_reg
	always @(*) begin
		if (andOp_253_out) begin 
			arg_2_write_valid_reg = -(1'd1);
		end else begin
			arg_2_write_valid_reg = 0;
		end
	end
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_115_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_159_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_6.bb_10_active_in_state_6_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_6_in_data = orOp_145_out;
		end else begin
			bb_10_active_in_state_6_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_6.bb_10_predecessor_in_state_6_in_data
	always @(*) begin
		if (andOp_201_out) begin 
			bb_10_predecessor_in_state_6_in_data = 32'd9;
		end else if (eq_199_out) begin 
			bb_10_predecessor_in_state_6_in_data = state_6_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_6_in_data = 0;
		end
	end
	// controller for bb_11_active_in_state_7.bb_11_active_in_state_7_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_11_active_in_state_7_in_data = eq_146_out;
		end else begin
			bb_11_active_in_state_7_in_data = 0;
		end
	end
	// controller for bb_11_active_in_state_8.bb_11_active_in_state_8_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_11_active_in_state_8_in_data = eq_153_out;
		end else begin
			bb_11_active_in_state_8_in_data = 0;
		end
	end
	// controller for bb_11_predecessor_in_state_7.bb_11_predecessor_in_state_7_in_data
	always @(*) begin
		if (eq_202_out) begin 
			bb_11_predecessor_in_state_7_in_data = state_7_last_BB_reg;
		end else begin
			bb_11_predecessor_in_state_7_in_data = 0;
		end
	end
	// controller for bb_11_predecessor_in_state_8.bb_11_predecessor_in_state_8_in_data
	always @(*) begin
		if (eq_212_out) begin 
			bb_11_predecessor_in_state_8_in_data = state_8_last_BB_reg;
		end else begin
			bb_11_predecessor_in_state_8_in_data = 0;
		end
	end
	// controller for bb_12_active_in_state_8.bb_12_active_in_state_8_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_12_active_in_state_8_in_data = orOp_157_out;
		end else begin
			bb_12_active_in_state_8_in_data = 0;
		end
	end
	// controller for bb_12_predecessor_in_state_8.bb_12_predecessor_in_state_8_in_data
	always @(*) begin
		if (andOp_218_out) begin 
			bb_12_predecessor_in_state_8_in_data = 32'd2;
		end else if (eq_216_out) begin 
			bb_12_predecessor_in_state_8_in_data = state_8_last_BB_reg;
		end else begin
			bb_12_predecessor_in_state_8_in_data = 0;
		end
	end
	// controller for bb_13_active_in_state_8.bb_13_active_in_state_8_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_13_active_in_state_8_in_data = orOp_148_out;
		end else begin
			bb_13_active_in_state_8_in_data = 0;
		end
	end
	// controller for bb_13_predecessor_in_state_8.bb_13_predecessor_in_state_8_in_data
	always @(*) begin
		if (andOp_205_out) begin 
			bb_13_predecessor_in_state_8_in_data = 32'd12;
		end else if (eq_203_out) begin 
			bb_13_predecessor_in_state_8_in_data = state_8_last_BB_reg;
		end else begin
			bb_13_predecessor_in_state_8_in_data = 0;
		end
	end
	// controller for bb_14_active_in_state_8.bb_14_active_in_state_8_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_14_active_in_state_8_in_data = orOp_150_out;
		end else begin
			bb_14_active_in_state_8_in_data = 0;
		end
	end
	// controller for bb_14_predecessor_in_state_8.bb_14_predecessor_in_state_8_in_data
	always @(*) begin
		if (andOp_208_out) begin 
			bb_14_predecessor_in_state_8_in_data = 32'd13;
		end else if (eq_206_out) begin 
			bb_14_predecessor_in_state_8_in_data = state_8_last_BB_reg;
		end else begin
			bb_14_predecessor_in_state_8_in_data = 0;
		end
	end
	// controller for bb_15_active_in_state_1.bb_15_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_15_active_in_state_1_in_data = orOp_117_out;
		end else begin
			bb_15_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_15_predecessor_in_state_1.bb_15_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_162_out) begin 
			bb_15_predecessor_in_state_1_in_data = 32'd4;
		end else if (eq_160_out) begin 
			bb_15_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_15_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_16_active_in_state_1.bb_16_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_16_active_in_state_1_in_data = orOp_120_out;
		end else begin
			bb_16_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_16_predecessor_in_state_1.bb_16_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_166_out) begin 
			bb_16_predecessor_in_state_1_in_data = 32'd15;
		end else if (eq_164_out) begin 
			bb_16_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_16_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_17_active_in_state_2.bb_17_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_17_active_in_state_2_in_data = eq_121_out;
		end else begin
			bb_17_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_17_active_in_state_3.bb_17_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_17_active_in_state_3_in_data = eq_122_out;
		end else begin
			bb_17_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_17_predecessor_in_state_2.bb_17_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_167_out) begin 
			bb_17_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_17_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_17_predecessor_in_state_3.bb_17_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_168_out) begin 
			bb_17_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_17_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_18_active_in_state_3.bb_18_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_18_active_in_state_3_in_data = orOp_124_out;
		end else begin
			bb_18_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_18_predecessor_in_state_3.bb_18_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_171_out) begin 
			bb_18_predecessor_in_state_3_in_data = 32'd5;
		end else if (eq_169_out) begin 
			bb_18_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_18_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_19_active_in_state_3.bb_19_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_19_active_in_state_3_in_data = orOp_126_out;
		end else begin
			bb_19_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_19_predecessor_in_state_3.bb_19_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_174_out) begin 
			bb_19_predecessor_in_state_3_in_data = 32'd18;
		end else if (eq_172_out) begin 
			bb_19_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_19_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_6.bb_1_active_in_state_6_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_6_in_data = eq_143_out;
		end else begin
			bb_1_active_in_state_6_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_6.bb_1_predecessor_in_state_6_in_data
	always @(*) begin
		if (eq_198_out) begin 
			bb_1_predecessor_in_state_6_in_data = state_6_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_6_in_data = 0;
		end
	end
	// controller for bb_20_active_in_state_4.bb_20_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_20_active_in_state_4_in_data = eq_129_out;
		end else begin
			bb_20_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_20_active_in_state_5.bb_20_active_in_state_5_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_20_active_in_state_5_in_data = eq_138_out;
		end else begin
			bb_20_active_in_state_5_in_data = 0;
		end
	end
	// controller for bb_20_predecessor_in_state_4.bb_20_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_178_out) begin 
			bb_20_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_20_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_20_predecessor_in_state_5.bb_20_predecessor_in_state_5_in_data
	always @(*) begin
		if (eq_191_out) begin 
			bb_20_predecessor_in_state_5_in_data = state_5_last_BB_reg;
		end else begin
			bb_20_predecessor_in_state_5_in_data = 0;
		end
	end
	// controller for bb_21_active_in_state_5.bb_21_active_in_state_5_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_21_active_in_state_5_in_data = orOp_137_out;
		end else begin
			bb_21_active_in_state_5_in_data = 0;
		end
	end
	// controller for bb_21_predecessor_in_state_5.bb_21_predecessor_in_state_5_in_data
	always @(*) begin
		if (andOp_190_out) begin 
			bb_21_predecessor_in_state_5_in_data = 32'd6;
		end else if (eq_188_out) begin 
			bb_21_predecessor_in_state_5_in_data = state_5_last_BB_reg;
		end else begin
			bb_21_predecessor_in_state_5_in_data = 0;
		end
	end
	// controller for bb_22_active_in_state_5.bb_22_active_in_state_5_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_22_active_in_state_5_in_data = orOp_131_out;
		end else begin
			bb_22_active_in_state_5_in_data = 0;
		end
	end
	// controller for bb_22_predecessor_in_state_5.bb_22_predecessor_in_state_5_in_data
	always @(*) begin
		if (andOp_181_out) begin 
			bb_22_predecessor_in_state_5_in_data = 32'd21;
		end else if (eq_179_out) begin 
			bb_22_predecessor_in_state_5_in_data = state_5_last_BB_reg;
		end else begin
			bb_22_predecessor_in_state_5_in_data = 0;
		end
	end
	// controller for bb_23_active_in_state_5.bb_23_active_in_state_5_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_23_active_in_state_5_in_data = orOp_133_out;
		end else begin
			bb_23_active_in_state_5_in_data = 0;
		end
	end
	// controller for bb_23_predecessor_in_state_5.bb_23_predecessor_in_state_5_in_data
	always @(*) begin
		if (andOp_184_out) begin 
			bb_23_predecessor_in_state_5_in_data = 32'd22;
		end else if (eq_182_out) begin 
			bb_23_predecessor_in_state_5_in_data = state_5_last_BB_reg;
		end else begin
			bb_23_predecessor_in_state_5_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_8.bb_2_active_in_state_8_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_8_in_data = orOp_152_out;
		end else begin
			bb_2_active_in_state_8_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_8.bb_2_predecessor_in_state_8_in_data
	always @(*) begin
		if (andOp_211_out) begin 
			bb_2_predecessor_in_state_8_in_data = 32'd11;
		end else if (eq_209_out) begin 
			bb_2_predecessor_in_state_8_in_data = state_8_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_8_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_8.bb_3_active_in_state_8_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_8_in_data = orOp_155_out;
		end else begin
			bb_3_active_in_state_8_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_8.bb_3_predecessor_in_state_8_in_data
	always @(*) begin
		if (andOp_215_out) begin 
			bb_3_predecessor_in_state_8_in_data = 32'd14;
		end else if (eq_213_out) begin 
			bb_3_predecessor_in_state_8_in_data = state_8_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_8_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_1.bb_4_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_1_in_data = eq_118_out;
		end else begin
			bb_4_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_1.bb_4_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_163_out) begin 
			bb_4_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_5_active_in_state_3.bb_5_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_5_active_in_state_3_in_data = orOp_128_out;
		end else begin
			bb_5_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_5_predecessor_in_state_3.bb_5_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_177_out) begin 
			bb_5_predecessor_in_state_3_in_data = 32'd17;
		end else if (eq_175_out) begin 
			bb_5_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_5_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_6_active_in_state_5.bb_6_active_in_state_5_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_6_active_in_state_5_in_data = orOp_140_out;
		end else begin
			bb_6_active_in_state_5_in_data = 0;
		end
	end
	// controller for bb_6_predecessor_in_state_5.bb_6_predecessor_in_state_5_in_data
	always @(*) begin
		if (andOp_194_out) begin 
			bb_6_predecessor_in_state_5_in_data = 32'd20;
		end else if (eq_192_out) begin 
			bb_6_predecessor_in_state_5_in_data = state_5_last_BB_reg;
		end else begin
			bb_6_predecessor_in_state_5_in_data = 0;
		end
	end
	// controller for bb_7_active_in_state_5.bb_7_active_in_state_5_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_7_active_in_state_5_in_data = orOp_135_out;
		end else begin
			bb_7_active_in_state_5_in_data = 0;
		end
	end
	// controller for bb_7_predecessor_in_state_5.bb_7_predecessor_in_state_5_in_data
	always @(*) begin
		if (andOp_187_out) begin 
			bb_7_predecessor_in_state_5_in_data = 32'd23;
		end else if (eq_185_out) begin 
			bb_7_predecessor_in_state_5_in_data = state_5_last_BB_reg;
		end else begin
			bb_7_predecessor_in_state_5_in_data = 0;
		end
	end
	// controller for bb_8_active_in_state_9.bb_8_active_in_state_9_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_state_9_in_data = eq_158_out;
		end else begin
			bb_8_active_in_state_9_in_data = 0;
		end
	end
	// controller for bb_8_predecessor_in_state_9.bb_8_predecessor_in_state_9_in_data
	always @(*) begin
		if (eq_219_out) begin 
			bb_8_predecessor_in_state_9_in_data = state_9_last_BB_reg;
		end else begin
			bb_8_predecessor_in_state_9_in_data = 0;
		end
	end
	// controller for bb_9_active_in_state_6.bb_9_active_in_state_6_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_9_active_in_state_6_in_data = orOp_142_out;
		end else begin
			bb_9_active_in_state_6_in_data = 0;
		end
	end
	// controller for bb_9_predecessor_in_state_6.bb_9_predecessor_in_state_6_in_data
	always @(*) begin
		if (andOp_197_out) begin 
			bb_9_predecessor_in_state_6_in_data = 32'd1;
		end else if (eq_195_out) begin 
			bb_9_predecessor_in_state_6_in_data = state_6_last_BB_reg;
		end else begin
			bb_9_predecessor_in_state_6_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_42_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_43_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_6.br_10_happened_in_state_6_in_data
	always @(*) begin
		if (andOp_90_out) begin 
			br_10_happened_in_state_6_in_data = 1'd1;
		end else if (notOp_91_out) begin 
			br_10_happened_in_state_6_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_6_in_data = 0;
		end
	end
	// controller for br_11_happened_in_state_7.br_11_happened_in_state_7_in_data
	always @(*) begin
		if (andOp_95_out) begin 
			br_11_happened_in_state_7_in_data = 1'd1;
		end else if (notOp_96_out) begin 
			br_11_happened_in_state_7_in_data = 1'd0;
		end else begin
			br_11_happened_in_state_7_in_data = 0;
		end
	end
	// controller for br_11_happened_in_state_8.br_11_happened_in_state_8_in_data
	always @(*) begin
		if (andOp_106_out) begin 
			br_11_happened_in_state_8_in_data = 1'd1;
		end else if (notOp_107_out) begin 
			br_11_happened_in_state_8_in_data = 1'd0;
		end else begin
			br_11_happened_in_state_8_in_data = 0;
		end
	end
	// controller for br_12_happened_in_state_8.br_12_happened_in_state_8_in_data
	always @(*) begin
		if (andOp_113_out) begin 
			br_12_happened_in_state_8_in_data = 1'd1;
		end else if (notOp_114_out) begin 
			br_12_happened_in_state_8_in_data = 1'd0;
		end else begin
			br_12_happened_in_state_8_in_data = 0;
		end
	end
	// controller for br_13_happened_in_state_8.br_13_happened_in_state_8_in_data
	always @(*) begin
		if (andOp_97_out) begin 
			br_13_happened_in_state_8_in_data = 1'd1;
		end else if (notOp_98_out) begin 
			br_13_happened_in_state_8_in_data = 1'd0;
		end else begin
			br_13_happened_in_state_8_in_data = 0;
		end
	end
	// controller for br_14_happened_in_state_8.br_14_happened_in_state_8_in_data
	always @(*) begin
		if (andOp_102_out) begin 
			br_14_happened_in_state_8_in_data = 1'd1;
		end else if (notOp_103_out) begin 
			br_14_happened_in_state_8_in_data = 1'd0;
		end else begin
			br_14_happened_in_state_8_in_data = 0;
		end
	end
	// controller for br_15_happened_in_state_1.br_15_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_44_out) begin 
			br_15_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_45_out) begin 
			br_15_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_15_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_16_happened_in_state_1.br_16_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_48_out) begin 
			br_16_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_49_out) begin 
			br_16_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_16_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_17_happened_in_state_2.br_17_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_53_out) begin 
			br_17_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_54_out) begin 
			br_17_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_17_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_17_happened_in_state_3.br_17_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_55_out) begin 
			br_17_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_56_out) begin 
			br_17_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_17_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_18_happened_in_state_3.br_18_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_57_out) begin 
			br_18_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_58_out) begin 
			br_18_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_18_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_19_happened_in_state_3.br_19_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_59_out) begin 
			br_19_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_60_out) begin 
			br_19_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_19_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_1_happened_in_state_6.br_1_happened_in_state_6_in_data
	always @(*) begin
		if (andOp_88_out) begin 
			br_1_happened_in_state_6_in_data = 1'd1;
		end else if (notOp_89_out) begin 
			br_1_happened_in_state_6_in_data = 1'd0;
		end else begin
			br_1_happened_in_state_6_in_data = 0;
		end
	end
	// controller for br_20_happened_in_state_4.br_20_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_66_out) begin 
			br_20_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_67_out) begin 
			br_20_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_20_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_20_happened_in_state_5.br_20_happened_in_state_5_in_data
	always @(*) begin
		if (andOp_82_out) begin 
			br_20_happened_in_state_5_in_data = 1'd1;
		end else if (notOp_83_out) begin 
			br_20_happened_in_state_5_in_data = 1'd0;
		end else begin
			br_20_happened_in_state_5_in_data = 0;
		end
	end
	// controller for br_21_happened_in_state_5.br_21_happened_in_state_5_in_data
	always @(*) begin
		if (andOp_80_out) begin 
			br_21_happened_in_state_5_in_data = 1'd1;
		end else if (notOp_81_out) begin 
			br_21_happened_in_state_5_in_data = 1'd0;
		end else begin
			br_21_happened_in_state_5_in_data = 0;
		end
	end
	// controller for br_22_happened_in_state_5.br_22_happened_in_state_5_in_data
	always @(*) begin
		if (andOp_68_out) begin 
			br_22_happened_in_state_5_in_data = 1'd1;
		end else if (notOp_69_out) begin 
			br_22_happened_in_state_5_in_data = 1'd0;
		end else begin
			br_22_happened_in_state_5_in_data = 0;
		end
	end
	// controller for br_23_happened_in_state_5.br_23_happened_in_state_5_in_data
	always @(*) begin
		if (andOp_73_out) begin 
			br_23_happened_in_state_5_in_data = 1'd1;
		end else if (notOp_74_out) begin 
			br_23_happened_in_state_5_in_data = 1'd0;
		end else begin
			br_23_happened_in_state_5_in_data = 0;
		end
	end
	// controller for br_2_happened_in_state_8.br_2_happened_in_state_8_in_data
	always @(*) begin
		if (andOp_104_out) begin 
			br_2_happened_in_state_8_in_data = 1'd1;
		end else if (notOp_105_out) begin 
			br_2_happened_in_state_8_in_data = 1'd0;
		end else begin
			br_2_happened_in_state_8_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_8.br_3_happened_in_state_8_in_data
	always @(*) begin
		if (andOp_108_out) begin 
			br_3_happened_in_state_8_in_data = 1'd1;
		end else if (notOp_109_out) begin 
			br_3_happened_in_state_8_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_8_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_1.br_4_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_46_out) begin 
			br_4_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_47_out) begin 
			br_4_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_5_happened_in_state_3.br_5_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_64_out) begin 
			br_5_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_65_out) begin 
			br_5_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_5_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_6_happened_in_state_5.br_6_happened_in_state_5_in_data
	always @(*) begin
		if (andOp_84_out) begin 
			br_6_happened_in_state_5_in_data = 1'd1;
		end else if (notOp_85_out) begin 
			br_6_happened_in_state_5_in_data = 1'd0;
		end else begin
			br_6_happened_in_state_5_in_data = 0;
		end
	end
	// controller for br_7_happened_in_state_5.br_7_happened_in_state_5_in_data
	always @(*) begin
		if (andOp_75_out) begin 
			br_7_happened_in_state_5_in_data = 1'd1;
		end else if (notOp_76_out) begin 
			br_7_happened_in_state_5_in_data = 1'd0;
		end else begin
			br_7_happened_in_state_5_in_data = 0;
		end
	end
	// controller for br_9_happened_in_state_6.br_9_happened_in_state_6_in_data
	always @(*) begin
		if (andOp_86_out) begin 
			br_9_happened_in_state_6_in_data = 1'd1;
		end else if (notOp_87_out) begin 
			br_9_happened_in_state_6_in_data = 1'd0;
		end else begin
			br_9_happened_in_state_6_in_data = 0;
		end
	end
	// controller for concat_231.concat_231_in0
	// controller for concat_231.concat_231_in1
	// Insensitive connections
	assign concat_231_in0 = data_in_1_1_out_data;
	assign concat_231_in1 = 32'd0;
	// controller for concat_232.concat_232_in0
	// controller for concat_232.concat_232_in1
	// Insensitive connections
	assign concat_232_in0 = 32'd7;
	assign concat_232_in1 = 32'd0;
	// controller for concat_246.concat_246_in0
	// controller for concat_246.concat_246_in1
	// Insensitive connections
	assign concat_246_in0 = data_in_6_33_out_data;
	assign concat_246_in1 = 32'd0;
	// controller for concat_247.concat_247_in0
	// controller for concat_247.concat_247_in1
	// Insensitive connections
	assign concat_247_in0 = 32'd3;
	assign concat_247_in1 = 32'd7;
	// controller for data_in_1_1.data_in_1_1_in_data
	always @(*) begin
		if (eq_303_out) begin 
			data_in_1_1_in_data = 32'd0;
		end else if (eq_304_out) begin 
			data_in_1_1_in_data = data_store_1_0;
		end else if (eq_305_out) begin 
			data_in_1_1_in_data = data_store_5_24;
		end else begin
			data_in_1_1_in_data = 0;
		end
	end
	// controller for data_in_1_3.data_in_1_3_in_data
	always @(*) begin
		if (eq_303_out) begin 
			data_in_1_3_in_data = 32'd0;
		end else if (eq_304_out) begin 
			data_in_1_3_in_data = data_store_1_2;
		end else if (eq_305_out) begin 
			data_in_1_3_in_data = data_store_5_26;
		end else begin
			data_in_1_3_in_data = 0;
		end
	end
	// controller for data_in_1_5.data_in_1_5_in_data
	always @(*) begin
		if (eq_303_out) begin 
			data_in_1_5_in_data = 32'd0;
		end else if (eq_304_out) begin 
			data_in_1_5_in_data = data_store_1_4;
		end else if (eq_305_out) begin 
			data_in_1_5_in_data = data_store_5_28;
		end else begin
			data_in_1_5_in_data = 0;
		end
	end
	// controller for data_in_2_11.data_in_2_11_in_data
	always @(*) begin
		if (eq_307_out) begin 
			data_in_2_11_in_data = data_store_1_4;
		end else if (eq_308_out) begin 
			data_in_2_11_in_data = data_store_2_10;
		end else begin
			data_in_2_11_in_data = 0;
		end
	end
	// controller for data_in_2_7.data_in_2_7_in_data
	always @(*) begin
		if (eq_307_out) begin 
			data_in_2_7_in_data = data_store_1_0;
		end else if (eq_308_out) begin 
			data_in_2_7_in_data = data_store_2_6;
		end else begin
			data_in_2_7_in_data = 0;
		end
	end
	// controller for data_in_2_9.data_in_2_9_in_data
	always @(*) begin
		if (eq_307_out) begin 
			data_in_2_9_in_data = data_store_1_2;
		end else if (eq_308_out) begin 
			data_in_2_9_in_data = data_store_2_8;
		end else begin
			data_in_2_9_in_data = 0;
		end
	end
	// controller for data_in_3_13.data_in_3_13_in_data
	always @(*) begin
		if (eq_309_out) begin 
			data_in_3_13_in_data = data_store_2_6;
		end else if (eq_310_out) begin 
			data_in_3_13_in_data = data_store_3_12;
		end else begin
			data_in_3_13_in_data = 0;
		end
	end
	// controller for data_in_3_15.data_in_3_15_in_data
	always @(*) begin
		if (eq_309_out) begin 
			data_in_3_15_in_data = data_store_2_8;
		end else if (eq_310_out) begin 
			data_in_3_15_in_data = data_store_3_14;
		end else begin
			data_in_3_15_in_data = 0;
		end
	end
	// controller for data_in_3_17.data_in_3_17_in_data
	always @(*) begin
		if (eq_309_out) begin 
			data_in_3_17_in_data = data_store_2_10;
		end else if (eq_310_out) begin 
			data_in_3_17_in_data = data_store_3_16;
		end else begin
			data_in_3_17_in_data = 0;
		end
	end
	// controller for data_in_4_19.data_in_4_19_in_data
	always @(*) begin
		if (eq_312_out) begin 
			data_in_4_19_in_data = data_store_3_12;
		end else if (eq_313_out) begin 
			data_in_4_19_in_data = data_store_4_18;
		end else begin
			data_in_4_19_in_data = 0;
		end
	end
	// controller for data_in_4_21.data_in_4_21_in_data
	always @(*) begin
		if (eq_312_out) begin 
			data_in_4_21_in_data = data_store_3_14;
		end else if (eq_313_out) begin 
			data_in_4_21_in_data = data_store_4_20;
		end else begin
			data_in_4_21_in_data = 0;
		end
	end
	// controller for data_in_4_23.data_in_4_23_in_data
	always @(*) begin
		if (eq_312_out) begin 
			data_in_4_23_in_data = data_store_3_16;
		end else if (eq_313_out) begin 
			data_in_4_23_in_data = data_store_4_22;
		end else begin
			data_in_4_23_in_data = 0;
		end
	end
	// controller for data_in_5_25.data_in_5_25_in_data
	always @(*) begin
		if (eq_314_out) begin 
			data_in_5_25_in_data = data_store_4_18;
		end else if (eq_315_out) begin 
			data_in_5_25_in_data = data_store_5_24;
		end else begin
			data_in_5_25_in_data = 0;
		end
	end
	// controller for data_in_5_27.data_in_5_27_in_data
	always @(*) begin
		if (eq_314_out) begin 
			data_in_5_27_in_data = data_store_4_20;
		end else if (eq_315_out) begin 
			data_in_5_27_in_data = data_store_5_26;
		end else begin
			data_in_5_27_in_data = 0;
		end
	end
	// controller for data_in_5_29.data_in_5_29_in_data
	always @(*) begin
		if (eq_314_out) begin 
			data_in_5_29_in_data = data_store_4_22;
		end else if (eq_315_out) begin 
			data_in_5_29_in_data = data_store_5_28;
		end else begin
			data_in_5_29_in_data = 0;
		end
	end
	// controller for data_in_6_31.data_in_6_31_in_data
	always @(*) begin
		if (eq_317_out) begin 
			data_in_6_31_in_data = 32'd0;
		end else if (eq_318_out) begin 
			data_in_6_31_in_data = data_store_6_30;
		end else if (eq_319_out) begin 
			data_in_6_31_in_data = data_store_8_38;
		end else begin
			data_in_6_31_in_data = 0;
		end
	end
	// controller for data_in_6_33.data_in_6_33_in_data
	always @(*) begin
		if (eq_317_out) begin 
			data_in_6_33_in_data = 32'd0;
		end else if (eq_318_out) begin 
			data_in_6_33_in_data = data_store_6_32;
		end else if (eq_319_out) begin 
			data_in_6_33_in_data = data_store_8_40;
		end else begin
			data_in_6_33_in_data = 0;
		end
	end
	// controller for data_in_7_35.data_in_7_35_in_data
	always @(*) begin
		if (eq_321_out) begin 
			data_in_7_35_in_data = data_store_6_30;
		end else if (eq_322_out) begin 
			data_in_7_35_in_data = data_store_7_34;
		end else begin
			data_in_7_35_in_data = 0;
		end
	end
	// controller for data_in_7_37.data_in_7_37_in_data
	always @(*) begin
		if (eq_321_out) begin 
			data_in_7_37_in_data = data_store_6_32;
		end else if (eq_322_out) begin 
			data_in_7_37_in_data = data_store_7_36;
		end else begin
			data_in_7_37_in_data = 0;
		end
	end
	// controller for data_in_8_39.data_in_8_39_in_data
	always @(*) begin
		if (eq_323_out) begin 
			data_in_8_39_in_data = data_store_7_34;
		end else if (eq_324_out) begin 
			data_in_8_39_in_data = data_store_8_38;
		end else begin
			data_in_8_39_in_data = 0;
		end
	end
	// controller for data_in_8_41.data_in_8_41_in_data
	always @(*) begin
		if (eq_323_out) begin 
			data_in_8_41_in_data = data_store_7_36;
		end else if (eq_324_out) begin 
			data_in_8_41_in_data = data_store_8_40;
		end else begin
			data_in_8_41_in_data = 0;
		end
	end
	// controller for eq_115.eq_115_in0
	// controller for eq_115.eq_115_in1
	// Insensitive connections
	assign eq_115_in0 = 32'd0;
	assign eq_115_in1 = state_0_entry_BB_reg;
	// controller for eq_116.eq_116_in0
	// controller for eq_116.eq_116_in1
	// Insensitive connections
	assign eq_116_in0 = 32'd15;
	assign eq_116_in1 = state_1_entry_BB_reg;
	// controller for eq_118.eq_118_in0
	// controller for eq_118.eq_118_in1
	// Insensitive connections
	assign eq_118_in0 = 32'd4;
	assign eq_118_in1 = state_1_entry_BB_reg;
	// controller for eq_119.eq_119_in0
	// controller for eq_119.eq_119_in1
	// Insensitive connections
	assign eq_119_in0 = 32'd16;
	assign eq_119_in1 = state_1_entry_BB_reg;
	// controller for eq_121.eq_121_in0
	// controller for eq_121.eq_121_in1
	// Insensitive connections
	assign eq_121_in0 = 32'd17;
	assign eq_121_in1 = state_2_entry_BB_reg;
	// controller for eq_122.eq_122_in0
	// controller for eq_122.eq_122_in1
	// Insensitive connections
	assign eq_122_in0 = 32'd17;
	assign eq_122_in1 = state_3_entry_BB_reg;
	// controller for eq_123.eq_123_in0
	// controller for eq_123.eq_123_in1
	// Insensitive connections
	assign eq_123_in0 = 32'd18;
	assign eq_123_in1 = state_3_entry_BB_reg;
	// controller for eq_125.eq_125_in0
	// controller for eq_125.eq_125_in1
	// Insensitive connections
	assign eq_125_in0 = 32'd19;
	assign eq_125_in1 = state_3_entry_BB_reg;
	// controller for eq_127.eq_127_in0
	// controller for eq_127.eq_127_in1
	// Insensitive connections
	assign eq_127_in0 = 32'd5;
	assign eq_127_in1 = state_3_entry_BB_reg;
	// controller for eq_129.eq_129_in0
	// controller for eq_129.eq_129_in1
	// Insensitive connections
	assign eq_129_in0 = 32'd20;
	assign eq_129_in1 = state_4_entry_BB_reg;
	// controller for eq_130.eq_130_in0
	// controller for eq_130.eq_130_in1
	// Insensitive connections
	assign eq_130_in0 = 32'd22;
	assign eq_130_in1 = state_5_entry_BB_reg;
	// controller for eq_132.eq_132_in0
	// controller for eq_132.eq_132_in1
	// Insensitive connections
	assign eq_132_in0 = 32'd23;
	assign eq_132_in1 = state_5_entry_BB_reg;
	// controller for eq_134.eq_134_in0
	// controller for eq_134.eq_134_in1
	// Insensitive connections
	assign eq_134_in0 = 32'd7;
	assign eq_134_in1 = state_5_entry_BB_reg;
	// controller for eq_136.eq_136_in0
	// controller for eq_136.eq_136_in1
	// Insensitive connections
	assign eq_136_in0 = 32'd21;
	assign eq_136_in1 = state_5_entry_BB_reg;
	// controller for eq_138.eq_138_in0
	// controller for eq_138.eq_138_in1
	// Insensitive connections
	assign eq_138_in0 = 32'd20;
	assign eq_138_in1 = state_5_entry_BB_reg;
	// controller for eq_139.eq_139_in0
	// controller for eq_139.eq_139_in1
	// Insensitive connections
	assign eq_139_in0 = 32'd6;
	assign eq_139_in1 = state_5_entry_BB_reg;
	// controller for eq_141.eq_141_in0
	// controller for eq_141.eq_141_in1
	// Insensitive connections
	assign eq_141_in0 = 32'd9;
	assign eq_141_in1 = state_6_entry_BB_reg;
	// controller for eq_143.eq_143_in0
	// controller for eq_143.eq_143_in1
	// Insensitive connections
	assign eq_143_in0 = 32'd1;
	assign eq_143_in1 = state_6_entry_BB_reg;
	// controller for eq_144.eq_144_in0
	// controller for eq_144.eq_144_in1
	// Insensitive connections
	assign eq_144_in0 = 32'd10;
	assign eq_144_in1 = state_6_entry_BB_reg;
	// controller for eq_146.eq_146_in0
	// controller for eq_146.eq_146_in1
	// Insensitive connections
	assign eq_146_in0 = 32'd11;
	assign eq_146_in1 = state_7_entry_BB_reg;
	// controller for eq_147.eq_147_in0
	// controller for eq_147.eq_147_in1
	// Insensitive connections
	assign eq_147_in0 = 32'd13;
	assign eq_147_in1 = state_8_entry_BB_reg;
	// controller for eq_149.eq_149_in0
	// controller for eq_149.eq_149_in1
	// Insensitive connections
	assign eq_149_in0 = 32'd14;
	assign eq_149_in1 = state_8_entry_BB_reg;
	// controller for eq_151.eq_151_in0
	// controller for eq_151.eq_151_in1
	// Insensitive connections
	assign eq_151_in0 = 32'd2;
	assign eq_151_in1 = state_8_entry_BB_reg;
	// controller for eq_153.eq_153_in0
	// controller for eq_153.eq_153_in1
	// Insensitive connections
	assign eq_153_in0 = 32'd11;
	assign eq_153_in1 = state_8_entry_BB_reg;
	// controller for eq_154.eq_154_in0
	// controller for eq_154.eq_154_in1
	// Insensitive connections
	assign eq_154_in0 = 32'd3;
	assign eq_154_in1 = state_8_entry_BB_reg;
	// controller for eq_156.eq_156_in0
	// controller for eq_156.eq_156_in1
	// Insensitive connections
	assign eq_156_in0 = 32'd12;
	assign eq_156_in1 = state_8_entry_BB_reg;
	// controller for eq_158.eq_158_in0
	// controller for eq_158.eq_158_in1
	// Insensitive connections
	assign eq_158_in0 = 32'd8;
	assign eq_158_in1 = state_9_entry_BB_reg;
	// controller for eq_159.eq_159_in0
	// controller for eq_159.eq_159_in1
	// Insensitive connections
	assign eq_159_in0 = 32'd0;
	assign eq_159_in1 = state_0_entry_BB_reg;
	// controller for eq_160.eq_160_in0
	// controller for eq_160.eq_160_in1
	// Insensitive connections
	assign eq_160_in0 = 32'd15;
	assign eq_160_in1 = state_1_entry_BB_reg;
	// controller for eq_163.eq_163_in0
	// controller for eq_163.eq_163_in1
	// Insensitive connections
	assign eq_163_in0 = 32'd4;
	assign eq_163_in1 = state_1_entry_BB_reg;
	// controller for eq_164.eq_164_in0
	// controller for eq_164.eq_164_in1
	// Insensitive connections
	assign eq_164_in0 = 32'd16;
	assign eq_164_in1 = state_1_entry_BB_reg;
	// controller for eq_167.eq_167_in0
	// controller for eq_167.eq_167_in1
	// Insensitive connections
	assign eq_167_in0 = 32'd17;
	assign eq_167_in1 = state_2_entry_BB_reg;
	// controller for eq_168.eq_168_in0
	// controller for eq_168.eq_168_in1
	// Insensitive connections
	assign eq_168_in0 = 32'd17;
	assign eq_168_in1 = state_3_entry_BB_reg;
	// controller for eq_169.eq_169_in0
	// controller for eq_169.eq_169_in1
	// Insensitive connections
	assign eq_169_in0 = 32'd18;
	assign eq_169_in1 = state_3_entry_BB_reg;
	// controller for eq_172.eq_172_in0
	// controller for eq_172.eq_172_in1
	// Insensitive connections
	assign eq_172_in0 = 32'd19;
	assign eq_172_in1 = state_3_entry_BB_reg;
	// controller for eq_175.eq_175_in0
	// controller for eq_175.eq_175_in1
	// Insensitive connections
	assign eq_175_in0 = 32'd5;
	assign eq_175_in1 = state_3_entry_BB_reg;
	// controller for eq_178.eq_178_in0
	// controller for eq_178.eq_178_in1
	// Insensitive connections
	assign eq_178_in0 = 32'd20;
	assign eq_178_in1 = state_4_entry_BB_reg;
	// controller for eq_179.eq_179_in0
	// controller for eq_179.eq_179_in1
	// Insensitive connections
	assign eq_179_in0 = 32'd22;
	assign eq_179_in1 = state_5_entry_BB_reg;
	// controller for eq_182.eq_182_in0
	// controller for eq_182.eq_182_in1
	// Insensitive connections
	assign eq_182_in0 = 32'd23;
	assign eq_182_in1 = state_5_entry_BB_reg;
	// controller for eq_185.eq_185_in0
	// controller for eq_185.eq_185_in1
	// Insensitive connections
	assign eq_185_in0 = 32'd7;
	assign eq_185_in1 = state_5_entry_BB_reg;
	// controller for eq_188.eq_188_in0
	// controller for eq_188.eq_188_in1
	// Insensitive connections
	assign eq_188_in0 = 32'd21;
	assign eq_188_in1 = state_5_entry_BB_reg;
	// controller for eq_191.eq_191_in0
	// controller for eq_191.eq_191_in1
	// Insensitive connections
	assign eq_191_in0 = 32'd20;
	assign eq_191_in1 = state_5_entry_BB_reg;
	// controller for eq_192.eq_192_in0
	// controller for eq_192.eq_192_in1
	// Insensitive connections
	assign eq_192_in0 = 32'd6;
	assign eq_192_in1 = state_5_entry_BB_reg;
	// controller for eq_195.eq_195_in0
	// controller for eq_195.eq_195_in1
	// Insensitive connections
	assign eq_195_in0 = 32'd9;
	assign eq_195_in1 = state_6_entry_BB_reg;
	// controller for eq_198.eq_198_in0
	// controller for eq_198.eq_198_in1
	// Insensitive connections
	assign eq_198_in0 = 32'd1;
	assign eq_198_in1 = state_6_entry_BB_reg;
	// controller for eq_199.eq_199_in0
	// controller for eq_199.eq_199_in1
	// Insensitive connections
	assign eq_199_in0 = 32'd10;
	assign eq_199_in1 = state_6_entry_BB_reg;
	// controller for eq_202.eq_202_in0
	// controller for eq_202.eq_202_in1
	// Insensitive connections
	assign eq_202_in0 = 32'd11;
	assign eq_202_in1 = state_7_entry_BB_reg;
	// controller for eq_203.eq_203_in0
	// controller for eq_203.eq_203_in1
	// Insensitive connections
	assign eq_203_in0 = 32'd13;
	assign eq_203_in1 = state_8_entry_BB_reg;
	// controller for eq_206.eq_206_in0
	// controller for eq_206.eq_206_in1
	// Insensitive connections
	assign eq_206_in0 = 32'd14;
	assign eq_206_in1 = state_8_entry_BB_reg;
	// controller for eq_209.eq_209_in0
	// controller for eq_209.eq_209_in1
	// Insensitive connections
	assign eq_209_in0 = 32'd2;
	assign eq_209_in1 = state_8_entry_BB_reg;
	// controller for eq_212.eq_212_in0
	// controller for eq_212.eq_212_in1
	// Insensitive connections
	assign eq_212_in0 = 32'd11;
	assign eq_212_in1 = state_8_entry_BB_reg;
	// controller for eq_213.eq_213_in0
	// controller for eq_213.eq_213_in1
	// Insensitive connections
	assign eq_213_in0 = 32'd3;
	assign eq_213_in1 = state_8_entry_BB_reg;
	// controller for eq_216.eq_216_in0
	// controller for eq_216.eq_216_in1
	// Insensitive connections
	assign eq_216_in0 = 32'd12;
	assign eq_216_in1 = state_8_entry_BB_reg;
	// controller for eq_219.eq_219_in0
	// controller for eq_219.eq_219_in1
	// Insensitive connections
	assign eq_219_in0 = 32'd8;
	assign eq_219_in1 = state_9_entry_BB_reg;
	// controller for eq_225.eq_225_in0
	// controller for eq_225.eq_225_in1
	// Insensitive connections
	assign eq_225_in0 = 32'd22;
	assign eq_225_in1 = state_5_entry_BB_reg;
	// controller for eq_226.eq_226_in0
	// controller for eq_226.eq_226_in1
	// Insensitive connections
	assign eq_226_in0 = 32'd20;
	assign eq_226_in1 = state_5_entry_BB_reg;
	// controller for eq_243.eq_243_in0
	// controller for eq_243.eq_243_in1
	// Insensitive connections
	assign eq_243_in0 = 32'd22;
	assign eq_243_in1 = state_5_entry_BB_reg;
	// controller for eq_244.eq_244_in0
	// controller for eq_244.eq_244_in1
	// Insensitive connections
	assign eq_244_in0 = 32'd20;
	assign eq_244_in1 = state_5_entry_BB_reg;
	// controller for eq_251.eq_251_in0
	// controller for eq_251.eq_251_in1
	// Insensitive connections
	assign eq_251_in0 = 32'd13;
	assign eq_251_in1 = state_8_entry_BB_reg;
	// controller for eq_252.eq_252_in0
	// controller for eq_252.eq_252_in1
	// Insensitive connections
	assign eq_252_in0 = 32'd11;
	assign eq_252_in1 = state_8_entry_BB_reg;
	// controller for eq_258.eq_258_in0
	// controller for eq_258.eq_258_in1
	// Insensitive connections
	assign eq_258_in0 = 32'd13;
	assign eq_258_in1 = state_8_entry_BB_reg;
	// controller for eq_259.eq_259_in0
	// controller for eq_259.eq_259_in1
	// Insensitive connections
	assign eq_259_in0 = 32'd11;
	assign eq_259_in1 = state_8_entry_BB_reg;
	// controller for eq_302.eq_302_in0
	// controller for eq_302.eq_302_in1
	// Insensitive connections
	assign eq_302_in0 = 32'd0;
	assign eq_302_in1 = state_0_last_state;
	// controller for eq_303.eq_303_in0
	// controller for eq_303.eq_303_in1
	// Insensitive connections
	assign eq_303_in0 = 32'd0;
	assign eq_303_in1 = state_1_last_state;
	// controller for eq_304.eq_304_in0
	// controller for eq_304.eq_304_in1
	// Insensitive connections
	assign eq_304_in0 = 32'd1;
	assign eq_304_in1 = state_1_last_state;
	// controller for eq_305.eq_305_in0
	// controller for eq_305.eq_305_in1
	// Insensitive connections
	assign eq_305_in0 = 32'd5;
	assign eq_305_in1 = state_1_last_state;
	// controller for eq_307.eq_307_in0
	// controller for eq_307.eq_307_in1
	// Insensitive connections
	assign eq_307_in0 = 32'd1;
	assign eq_307_in1 = state_2_last_state;
	// controller for eq_308.eq_308_in0
	// controller for eq_308.eq_308_in1
	// Insensitive connections
	assign eq_308_in0 = 32'd2;
	assign eq_308_in1 = state_2_last_state;
	// controller for eq_309.eq_309_in0
	// controller for eq_309.eq_309_in1
	// Insensitive connections
	assign eq_309_in0 = 32'd2;
	assign eq_309_in1 = state_3_last_state;
	// controller for eq_310.eq_310_in0
	// controller for eq_310.eq_310_in1
	// Insensitive connections
	assign eq_310_in0 = 32'd3;
	assign eq_310_in1 = state_3_last_state;
	// controller for eq_312.eq_312_in0
	// controller for eq_312.eq_312_in1
	// Insensitive connections
	assign eq_312_in0 = 32'd3;
	assign eq_312_in1 = state_4_last_state;
	// controller for eq_313.eq_313_in0
	// controller for eq_313.eq_313_in1
	// Insensitive connections
	assign eq_313_in0 = 32'd4;
	assign eq_313_in1 = state_4_last_state;
	// controller for eq_314.eq_314_in0
	// controller for eq_314.eq_314_in1
	// Insensitive connections
	assign eq_314_in0 = 32'd4;
	assign eq_314_in1 = state_5_last_state;
	// controller for eq_315.eq_315_in0
	// controller for eq_315.eq_315_in1
	// Insensitive connections
	assign eq_315_in0 = 32'd5;
	assign eq_315_in1 = state_5_last_state;
	// controller for eq_317.eq_317_in0
	// controller for eq_317.eq_317_in1
	// Insensitive connections
	assign eq_317_in0 = 32'd5;
	assign eq_317_in1 = state_6_last_state;
	// controller for eq_318.eq_318_in0
	// controller for eq_318.eq_318_in1
	// Insensitive connections
	assign eq_318_in0 = 32'd6;
	assign eq_318_in1 = state_6_last_state;
	// controller for eq_319.eq_319_in0
	// controller for eq_319.eq_319_in1
	// Insensitive connections
	assign eq_319_in0 = 32'd8;
	assign eq_319_in1 = state_6_last_state;
	// controller for eq_321.eq_321_in0
	// controller for eq_321.eq_321_in1
	// Insensitive connections
	assign eq_321_in0 = 32'd6;
	assign eq_321_in1 = state_7_last_state;
	// controller for eq_322.eq_322_in0
	// controller for eq_322.eq_322_in1
	// Insensitive connections
	assign eq_322_in0 = 32'd7;
	assign eq_322_in1 = state_7_last_state;
	// controller for eq_323.eq_323_in0
	// controller for eq_323.eq_323_in1
	// Insensitive connections
	assign eq_323_in0 = 32'd7;
	assign eq_323_in1 = state_8_last_state;
	// controller for eq_324.eq_324_in0
	// controller for eq_324.eq_324_in1
	// Insensitive connections
	assign eq_324_in0 = 32'd8;
	assign eq_324_in1 = state_8_last_state;
	// controller for eq_326.eq_326_in0
	// controller for eq_326.eq_326_in1
	// Insensitive connections
	assign eq_326_in0 = 32'd8;
	assign eq_326_in1 = state_9_last_state;
	// controller for eq_327.eq_327_in0
	// controller for eq_327.eq_327_in1
	// Insensitive connections
	assign eq_327_in0 = 32'd9;
	assign eq_327_in1 = state_9_last_state;
	// controller for icmp_icmp16.icmp_icmp16_in0
	// controller for icmp_icmp16.icmp_icmp16_in1
	// Insensitive connections
	assign icmp_icmp16_in0 = data_in_5_25_out_data;
	assign icmp_icmp16_in1 = 32'd15;
	// controller for icmp_icmp37.icmp_icmp37_in0
	// controller for icmp_icmp37.icmp_icmp37_in1
	// Insensitive connections
	assign icmp_icmp37_in0 = data_in_8_41_out_data;
	assign icmp_icmp37_in1 = 32'd15;
	// controller for mul_mul39.mul_mul39_in0
	// controller for mul_mul39.mul_mul39_in1
	// Insensitive connections
	assign mul_mul39_in0 = 32'd2;
	assign mul_mul39_in1 = tmp_output_257_out_data;
	// controller for notOp_100.notOp_100_in0
	// Insensitive connections
	assign notOp_100_in0 = arg_2_write_ready;
	// controller for notOp_103.notOp_103_in0
	// Insensitive connections
	assign notOp_103_in0 = andOp_102_out;
	// controller for notOp_105.notOp_105_in0
	// Insensitive connections
	assign notOp_105_in0 = andOp_104_out;
	// controller for notOp_107.notOp_107_in0
	// Insensitive connections
	assign notOp_107_in0 = andOp_106_out;
	// controller for notOp_109.notOp_109_in0
	// Insensitive connections
	assign notOp_109_in0 = andOp_108_out;
	// controller for notOp_111.notOp_111_in0
	// Insensitive connections
	assign notOp_111_in0 = icmp_icmp37_out;
	// controller for notOp_114.notOp_114_in0
	// Insensitive connections
	assign notOp_114_in0 = andOp_113_out;
	// controller for notOp_161.notOp_161_in0
	// Insensitive connections
	assign notOp_161_in0 = eq_160_out;
	// controller for notOp_165.notOp_165_in0
	// Insensitive connections
	assign notOp_165_in0 = eq_164_out;
	// controller for notOp_170.notOp_170_in0
	// Insensitive connections
	assign notOp_170_in0 = eq_169_out;
	// controller for notOp_173.notOp_173_in0
	// Insensitive connections
	assign notOp_173_in0 = eq_172_out;
	// controller for notOp_176.notOp_176_in0
	// Insensitive connections
	assign notOp_176_in0 = eq_175_out;
	// controller for notOp_180.notOp_180_in0
	// Insensitive connections
	assign notOp_180_in0 = eq_179_out;
	// controller for notOp_183.notOp_183_in0
	// Insensitive connections
	assign notOp_183_in0 = eq_182_out;
	// controller for notOp_186.notOp_186_in0
	// Insensitive connections
	assign notOp_186_in0 = eq_185_out;
	// controller for notOp_189.notOp_189_in0
	// Insensitive connections
	assign notOp_189_in0 = eq_188_out;
	// controller for notOp_193.notOp_193_in0
	// Insensitive connections
	assign notOp_193_in0 = eq_192_out;
	// controller for notOp_196.notOp_196_in0
	// Insensitive connections
	assign notOp_196_in0 = eq_195_out;
	// controller for notOp_200.notOp_200_in0
	// Insensitive connections
	assign notOp_200_in0 = eq_199_out;
	// controller for notOp_204.notOp_204_in0
	// Insensitive connections
	assign notOp_204_in0 = eq_203_out;
	// controller for notOp_207.notOp_207_in0
	// Insensitive connections
	assign notOp_207_in0 = eq_206_out;
	// controller for notOp_210.notOp_210_in0
	// Insensitive connections
	assign notOp_210_in0 = eq_209_out;
	// controller for notOp_214.notOp_214_in0
	// Insensitive connections
	assign notOp_214_in0 = eq_213_out;
	// controller for notOp_217.notOp_217_in0
	// Insensitive connections
	assign notOp_217_in0 = eq_216_out;
	// controller for notOp_268.notOp_268_in0
	// Insensitive connections
	assign notOp_268_in0 = andOp_261_out;
	// controller for notOp_270.notOp_270_in0
	// Insensitive connections
	assign notOp_270_in0 = andOp_52_out;
	// controller for notOp_272.notOp_272_in0
	// Insensitive connections
	assign notOp_272_in0 = andOp_77_out;
	// controller for notOp_274.notOp_274_in0
	// Insensitive connections
	assign notOp_274_in0 = andOp_50_out;
	// controller for notOp_276.notOp_276_in0
	// Insensitive connections
	assign notOp_276_in0 = andOp_262_out;
	// controller for notOp_278.notOp_278_in0
	// Insensitive connections
	assign notOp_278_in0 = andOp_63_out;
	// controller for notOp_280.notOp_280_in0
	// Insensitive connections
	assign notOp_280_in0 = andOp_61_out;
	// controller for notOp_282.notOp_282_in0
	// Insensitive connections
	assign notOp_282_in0 = andOp_263_out;
	// controller for notOp_284.notOp_284_in0
	// Insensitive connections
	assign notOp_284_in0 = andOp_72_out;
	// controller for notOp_286.notOp_286_in0
	// Insensitive connections
	assign notOp_286_in0 = andOp_110_out;
	// controller for notOp_288.notOp_288_in0
	// Insensitive connections
	assign notOp_288_in0 = andOp_264_out;
	// controller for notOp_290.notOp_290_in0
	// Insensitive connections
	assign notOp_290_in0 = andOp_94_out;
	// controller for notOp_292.notOp_292_in0
	// Insensitive connections
	assign notOp_292_in0 = andOp_92_out;
	// controller for notOp_294.notOp_294_in0
	// Insensitive connections
	assign notOp_294_in0 = andOp_101_out;
	// controller for notOp_296.notOp_296_in0
	// Insensitive connections
	assign notOp_296_in0 = andOp_265_out;
	// controller for notOp_298.notOp_298_in0
	// Insensitive connections
	assign notOp_298_in0 = andOp_266_out;
	// controller for notOp_300.notOp_300_in0
	// Insensitive connections
	assign notOp_300_in0 = andOp_267_out;
	// controller for notOp_43.notOp_43_in0
	// Insensitive connections
	assign notOp_43_in0 = andOp_42_out;
	// controller for notOp_45.notOp_45_in0
	// Insensitive connections
	assign notOp_45_in0 = andOp_44_out;
	// controller for notOp_47.notOp_47_in0
	// Insensitive connections
	assign notOp_47_in0 = andOp_46_out;
	// controller for notOp_49.notOp_49_in0
	// Insensitive connections
	assign notOp_49_in0 = andOp_48_out;
	// controller for notOp_51.notOp_51_in0
	// Insensitive connections
	assign notOp_51_in0 = arg_0_read_ready;
	// controller for notOp_54.notOp_54_in0
	// Insensitive connections
	assign notOp_54_in0 = andOp_53_out;
	// controller for notOp_56.notOp_56_in0
	// Insensitive connections
	assign notOp_56_in0 = andOp_55_out;
	// controller for notOp_58.notOp_58_in0
	// Insensitive connections
	assign notOp_58_in0 = andOp_57_out;
	// controller for notOp_60.notOp_60_in0
	// Insensitive connections
	assign notOp_60_in0 = andOp_59_out;
	// controller for notOp_62.notOp_62_in0
	// Insensitive connections
	assign notOp_62_in0 = arg_1_read_ready;
	// controller for notOp_65.notOp_65_in0
	// Insensitive connections
	assign notOp_65_in0 = andOp_64_out;
	// controller for notOp_67.notOp_67_in0
	// Insensitive connections
	assign notOp_67_in0 = andOp_66_out;
	// controller for notOp_69.notOp_69_in0
	// Insensitive connections
	assign notOp_69_in0 = andOp_68_out;
	// controller for notOp_71.notOp_71_in0
	// Insensitive connections
	assign notOp_71_in0 = _____dlr_0___eq___alloca___dlr_builtin_fifo_32_write_ready;
	// controller for notOp_74.notOp_74_in0
	// Insensitive connections
	assign notOp_74_in0 = andOp_73_out;
	// controller for notOp_76.notOp_76_in0
	// Insensitive connections
	assign notOp_76_in0 = andOp_75_out;
	// controller for notOp_78.notOp_78_in0
	// Insensitive connections
	assign notOp_78_in0 = icmp_icmp16_out;
	// controller for notOp_81.notOp_81_in0
	// Insensitive connections
	assign notOp_81_in0 = andOp_80_out;
	// controller for notOp_83.notOp_83_in0
	// Insensitive connections
	assign notOp_83_in0 = andOp_82_out;
	// controller for notOp_85.notOp_85_in0
	// Insensitive connections
	assign notOp_85_in0 = andOp_84_out;
	// controller for notOp_87.notOp_87_in0
	// Insensitive connections
	assign notOp_87_in0 = andOp_86_out;
	// controller for notOp_89.notOp_89_in0
	// Insensitive connections
	assign notOp_89_in0 = andOp_88_out;
	// controller for notOp_91.notOp_91_in0
	// Insensitive connections
	assign notOp_91_in0 = andOp_90_out;
	// controller for notOp_93.notOp_93_in0
	// Insensitive connections
	assign notOp_93_in0 = _____dlr_0___eq___alloca___dlr_builtin_fifo_32_read_ready;
	// controller for notOp_96.notOp_96_in0
	// Insensitive connections
	assign notOp_96_in0 = andOp_95_out;
	// controller for notOp_98.notOp_98_in0
	// Insensitive connections
	assign notOp_98_in0 = andOp_97_out;
	// controller for orOp_117.orOp_117_in0
	// controller for orOp_117.orOp_117_in1
	// Insensitive connections
	assign orOp_117_in0 = eq_116_out;
	assign orOp_117_in1 = andOp_46_out;
	// controller for orOp_120.orOp_120_in0
	// controller for orOp_120.orOp_120_in1
	// Insensitive connections
	assign orOp_120_in0 = eq_119_out;
	assign orOp_120_in1 = andOp_44_out;
	// controller for orOp_124.orOp_124_in0
	// controller for orOp_124.orOp_124_in1
	// Insensitive connections
	assign orOp_124_in0 = eq_123_out;
	assign orOp_124_in1 = andOp_64_out;
	// controller for orOp_126.orOp_126_in0
	// controller for orOp_126.orOp_126_in1
	// Insensitive connections
	assign orOp_126_in0 = eq_125_out;
	assign orOp_126_in1 = andOp_57_out;
	// controller for orOp_128.orOp_128_in0
	// controller for orOp_128.orOp_128_in1
	// Insensitive connections
	assign orOp_128_in0 = eq_127_out;
	assign orOp_128_in1 = andOp_53_out;
	// controller for orOp_131.orOp_131_in0
	// controller for orOp_131.orOp_131_in1
	// Insensitive connections
	assign orOp_131_in0 = eq_130_out;
	assign orOp_131_in1 = andOp_80_out;
	// controller for orOp_133.orOp_133_in0
	// controller for orOp_133.orOp_133_in1
	// Insensitive connections
	assign orOp_133_in0 = eq_132_out;
	assign orOp_133_in1 = andOp_70_out;
	// controller for orOp_135.orOp_135_in0
	// controller for orOp_135.orOp_135_in1
	// Insensitive connections
	assign orOp_135_in0 = eq_134_out;
	assign orOp_135_in1 = andOp_73_out;
	// controller for orOp_137.orOp_137_in0
	// controller for orOp_137.orOp_137_in1
	// Insensitive connections
	assign orOp_137_in0 = eq_136_out;
	assign orOp_137_in1 = andOp_84_out;
	// controller for orOp_140.orOp_140_in0
	// controller for orOp_140.orOp_140_in1
	// Insensitive connections
	assign orOp_140_in0 = eq_139_out;
	assign orOp_140_in1 = andOp_66_out;
	// controller for orOp_142.orOp_142_in0
	// controller for orOp_142.orOp_142_in1
	// Insensitive connections
	assign orOp_142_in0 = eq_141_out;
	assign orOp_142_in1 = andOp_88_out;
	// controller for orOp_145.orOp_145_in0
	// controller for orOp_145.orOp_145_in1
	// Insensitive connections
	assign orOp_145_in0 = eq_144_out;
	assign orOp_145_in1 = andOp_86_out;
	// controller for orOp_148.orOp_148_in0
	// controller for orOp_148.orOp_148_in1
	// Insensitive connections
	assign orOp_148_in0 = eq_147_out;
	assign orOp_148_in1 = andOp_113_out;
	// controller for orOp_150.orOp_150_in0
	// controller for orOp_150.orOp_150_in1
	// Insensitive connections
	assign orOp_150_in0 = eq_149_out;
	assign orOp_150_in1 = andOp_99_out;
	// controller for orOp_152.orOp_152_in0
	// controller for orOp_152.orOp_152_in1
	// Insensitive connections
	assign orOp_152_in0 = eq_151_out;
	assign orOp_152_in1 = andOp_95_out;
	// controller for orOp_155.orOp_155_in0
	// controller for orOp_155.orOp_155_in1
	// Insensitive connections
	assign orOp_155_in0 = eq_154_out;
	assign orOp_155_in1 = andOp_102_out;
	// controller for orOp_157.orOp_157_in0
	// controller for orOp_157.orOp_157_in1
	// Insensitive connections
	assign orOp_157_in0 = eq_156_out;
	assign orOp_157_in1 = andOp_104_out;
	// controller for phi_phi28.phi_phi28_in
	// controller for phi_phi28.phi_phi28_last_block
	// controller for phi_phi28.phi_phi28_s
	// Insensitive connections
	assign phi_phi28_in = concat_246_out;
	assign phi_phi28_last_block = bb_1_predecessor_in_state_6_out_data;
	assign phi_phi28_s = concat_247_out;
	// controller for phi_phi3.phi_phi3_in
	// controller for phi_phi3.phi_phi3_last_block
	// controller for phi_phi3.phi_phi3_s
	// Insensitive connections
	assign phi_phi3_in = concat_231_out;
	assign phi_phi3_last_block = bb_4_predecessor_in_state_1_out_data;
	assign phi_phi3_s = concat_232_out;
	// controller for ret47.valid_reg
	always @(*) begin
		if (andOp_260_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// controller for tmp_output_224.tmp_output_224_in_data
	always @(*) begin
		if (eq_225_out) begin 
			tmp_output_224_in_data = data_in_5_29_out_data;
		end else if (eq_226_out) begin 
			tmp_output_224_in_data = add_add26_out;
		end else begin
			tmp_output_224_in_data = 0;
		end
	end
	// controller for tmp_output_242.tmp_output_242_in_data
	always @(*) begin
		if (eq_244_out) begin 
			tmp_output_242_in_data = arg_1_out_data;
		end else begin
			tmp_output_242_in_data = 0;
		end
	end
	// controller for tmp_output_250.tmp_output_250_in_data
	always @(*) begin
		if (eq_251_out) begin 
			tmp_output_250_in_data = data_in_8_39_out_data;
		end else if (eq_252_out) begin 
			tmp_output_250_in_data = mul_mul39_out;
		end else begin
			tmp_output_250_in_data = 0;
		end
	end
	// controller for tmp_output_257.tmp_output_257_in_data
	always @(*) begin
		if (eq_259_out) begin 
			tmp_output_257_in_data = _____dlr_0___eq___alloca___dlr_builtin_fifo_32_out_data;
		end else begin
			tmp_output_257_in_data = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			data_store_1_0 <= 0;
		end else begin
			if (andOp_306_out) begin
				data_store_1_0 <= add_add5_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_2 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_2 <= data_in_1_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_4 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_4 <= data_in_1_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_10 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_10 <= data_in_2_11_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_6 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_6 <= data_in_2_7_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_8 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_8 <= data_in_2_9_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_12 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_12 <= data_in_3_13_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_14 <= 0;
		end else begin
			if (andOp_311_out) begin
				data_store_3_14 <= arg_0_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_16 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_16 <= data_in_3_17_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_18 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_18 <= data_in_4_19_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_20 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_20 <= data_in_4_21_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_22 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_22 <= data_in_4_23_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_24 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_24 <= data_in_5_25_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_26 <= 0;
		end else begin
			if (state_5_is_active) begin
				data_store_5_26 <= data_in_5_27_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_5_28 <= 0;
		end else begin
			if (andOp_316_out) begin
				data_store_5_28 <= add_add26_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_30 <= 0;
		end else begin
			if (state_6_is_active) begin
				data_store_6_30 <= data_in_6_31_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_6_32 <= 0;
		end else begin
			if (andOp_320_out) begin
				data_store_6_32 <= add_add29_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_7_34 <= 0;
		end else begin
			if (state_7_is_active) begin
				data_store_7_34 <= data_in_7_35_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_7_36 <= 0;
		end else begin
			if (state_7_is_active) begin
				data_store_7_36 <= data_in_7_37_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_8_38 <= 0;
		end else begin
			if (andOp_325_out) begin
				data_store_8_38 <= mul_mul39_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_8_40 <= 0;
		end else begin
			if (state_8_is_active) begin
				data_store_8_40 <= data_in_8_41_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_101_out) begin
				global_state <= 32'd8;
			end
			if (andOp_110_out) begin
				global_state <= 32'd6;
			end
			if (andOp_261_out) begin
				global_state <= 32'd1;
			end
			if (andOp_262_out) begin
				global_state <= 32'd3;
			end
			if (andOp_263_out) begin
				global_state <= 32'd5;
			end
			if (andOp_264_out) begin
				global_state <= 32'd6;
			end
			if (andOp_265_out) begin
				global_state <= 32'd8;
			end
			if (andOp_266_out) begin
				global_state <= 32'd9;
			end
			if (andOp_267_out) begin
				global_state <= 32'd9;
			end
			if (andOp_50_out) begin
				global_state <= 32'd2;
			end
			if (andOp_52_out) begin
				global_state <= 32'd1;
			end
			if (andOp_61_out) begin
				global_state <= 32'd4;
			end
			if (andOp_63_out) begin
				global_state <= 32'd3;
			end
			if (andOp_72_out) begin
				global_state <= 32'd5;
			end
			if (andOp_77_out) begin
				global_state <= 32'd1;
			end
			if (andOp_92_out) begin
				global_state <= 32'd7;
			end
			if (andOp_94_out) begin
				global_state <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (1'd1) begin
				state_0_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_261_out) begin
				state_1_entry_BB_reg <= 32'd4;
			end
			if (andOp_52_out) begin
				state_1_entry_BB_reg <= 32'd16;
			end
			if (andOp_77_out) begin
				state_1_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 1;
		end else begin
			if (andOp_261_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_273_out) begin
				state_1_is_active <= 1'd0;
			end
			if (andOp_52_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_77_out) begin
				state_1_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_261_out) begin
				state_1_last_BB_reg <= 32'd0;
			end
			if (andOp_52_out) begin
				state_1_last_BB_reg <= 32'd16;
			end
			if (andOp_77_out) begin
				state_1_last_BB_reg <= 32'd7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_261_out) begin
				state_1_last_state <= 32'd0;
			end
			if (andOp_52_out) begin
				state_1_last_state <= 32'd1;
			end
			if (andOp_77_out) begin
				state_1_last_state <= 32'd5;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_50_out) begin
				state_2_entry_BB_reg <= 32'd17;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_275_out) begin
				state_2_is_active <= 1'd0;
			end
			if (andOp_50_out) begin
				state_2_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_50_out) begin
				state_2_last_BB_reg <= 32'd16;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_50_out) begin
				state_2_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_262_out) begin
				state_3_entry_BB_reg <= 32'd17;
			end
			if (andOp_63_out) begin
				state_3_entry_BB_reg <= 32'd19;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_262_out) begin
				state_3_is_active <= 1'd1;
			end
			if (andOp_279_out) begin
				state_3_is_active <= 1'd0;
			end
			if (andOp_63_out) begin
				state_3_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_262_out) begin
				state_3_last_BB_reg <= bb_17_predecessor_in_state_2_out_data;
			end
			if (andOp_63_out) begin
				state_3_last_BB_reg <= 32'd19;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_state <= 0;
		end else begin
			if (andOp_262_out) begin
				state_3_last_state <= 32'd2;
			end
			if (andOp_63_out) begin
				state_3_last_state <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_61_out) begin
				state_4_entry_BB_reg <= 32'd20;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_281_out) begin
				state_4_is_active <= 1'd0;
			end
			if (andOp_61_out) begin
				state_4_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_61_out) begin
				state_4_last_BB_reg <= 32'd19;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_state <= 0;
		end else begin
			if (andOp_61_out) begin
				state_4_last_state <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_entry_BB_reg <= 0;
		end else begin
			if (andOp_263_out) begin
				state_5_entry_BB_reg <= 32'd20;
			end
			if (andOp_72_out) begin
				state_5_entry_BB_reg <= 32'd22;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_is_active <= 0;
		end else begin
			if (andOp_263_out) begin
				state_5_is_active <= 1'd1;
			end
			if (andOp_285_out) begin
				state_5_is_active <= 1'd0;
			end
			if (andOp_72_out) begin
				state_5_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_last_BB_reg <= 0;
		end else begin
			if (andOp_263_out) begin
				state_5_last_BB_reg <= bb_20_predecessor_in_state_4_out_data;
			end
			if (andOp_72_out) begin
				state_5_last_BB_reg <= 32'd22;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_5_last_state <= 0;
		end else begin
			if (andOp_263_out) begin
				state_5_last_state <= 32'd4;
			end
			if (andOp_72_out) begin
				state_5_last_state <= 32'd5;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_entry_BB_reg <= 0;
		end else begin
			if (andOp_110_out) begin
				state_6_entry_BB_reg <= 32'd1;
			end
			if (andOp_264_out) begin
				state_6_entry_BB_reg <= 32'd1;
			end
			if (andOp_94_out) begin
				state_6_entry_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_is_active <= 1;
		end else begin
			if (andOp_110_out) begin
				state_6_is_active <= 1'd1;
			end
			if (andOp_264_out) begin
				state_6_is_active <= 1'd1;
			end
			if (andOp_291_out) begin
				state_6_is_active <= 1'd0;
			end
			if (andOp_94_out) begin
				state_6_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_last_BB_reg <= 0;
		end else begin
			if (andOp_110_out) begin
				state_6_last_BB_reg <= 32'd3;
			end
			if (andOp_264_out) begin
				state_6_last_BB_reg <= 32'd7;
			end
			if (andOp_94_out) begin
				state_6_last_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_6_last_state <= 0;
		end else begin
			if (andOp_110_out) begin
				state_6_last_state <= 32'd8;
			end
			if (andOp_264_out) begin
				state_6_last_state <= 32'd5;
			end
			if (andOp_94_out) begin
				state_6_last_state <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_entry_BB_reg <= 0;
		end else begin
			if (andOp_92_out) begin
				state_7_entry_BB_reg <= 32'd11;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_is_active <= 0;
		end else begin
			if (andOp_293_out) begin
				state_7_is_active <= 1'd0;
			end
			if (andOp_92_out) begin
				state_7_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_last_BB_reg <= 0;
		end else begin
			if (andOp_92_out) begin
				state_7_last_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_7_last_state <= 0;
		end else begin
			if (andOp_92_out) begin
				state_7_last_state <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_8_entry_BB_reg <= 0;
		end else begin
			if (andOp_101_out) begin
				state_8_entry_BB_reg <= 32'd13;
			end
			if (andOp_265_out) begin
				state_8_entry_BB_reg <= 32'd11;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_8_is_active <= 0;
		end else begin
			if (andOp_101_out) begin
				state_8_is_active <= 1'd1;
			end
			if (andOp_265_out) begin
				state_8_is_active <= 1'd1;
			end
			if (andOp_297_out) begin
				state_8_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_8_last_BB_reg <= 0;
		end else begin
			if (andOp_101_out) begin
				state_8_last_BB_reg <= 32'd13;
			end
			if (andOp_265_out) begin
				state_8_last_BB_reg <= bb_11_predecessor_in_state_7_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_8_last_state <= 0;
		end else begin
			if (andOp_101_out) begin
				state_8_last_state <= 32'd8;
			end
			if (andOp_265_out) begin
				state_8_last_state <= 32'd7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_9_entry_BB_reg <= 0;
		end else begin
			if (andOp_266_out) begin
				state_9_entry_BB_reg <= 32'd8;
			end
			if (andOp_267_out) begin
				state_9_entry_BB_reg <= 32'd8;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_9_is_active <= 1;
		end else begin
			if (andOp_266_out) begin
				state_9_is_active <= 1'd1;
			end
			if (andOp_267_out) begin
				state_9_is_active <= 1'd1;
			end
			if (andOp_301_out) begin
				state_9_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_9_last_BB_reg <= 0;
		end else begin
			if (andOp_266_out) begin
				state_9_last_BB_reg <= 32'd3;
			end
			if (andOp_267_out) begin
				state_9_last_BB_reg <= bb_8_predecessor_in_state_9_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_9_last_state <= 0;
		end else begin
			if (andOp_266_out) begin
				state_9_last_state <= 32'd8;
			end
			if (andOp_267_out) begin
				state_9_last_state <= 32'd9;
			end
		end
	end

endmodule

