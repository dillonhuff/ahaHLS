module channel_reduce_4(input [0:0] clk, input [0:0] rst, output [0:0] valid, output [31:0] out_in_data, output [0:0] out_read_valid, output [0:0] out_rst, output [0:0] out_write_valid, input [31:0] out_out_data, input [0:0] out_read_ready, input [0:0] out_write_ready, output [31:0] in_in_data, output [0:0] in_read_valid, output [0:0] in_rst, output [0:0] in_write_valid, input [31:0] in_out_data, input [0:0] in_read_ready, input [0:0] in_write_ready);

	reg [0:0] valid_reg;
	reg [31:0] out_in_data_reg;
	reg [0:0] out_read_valid_reg;
	reg [0:0] out_rst_reg;
	reg [0:0] out_write_valid_reg;
	reg [31:0] in_in_data_reg;
	reg [0:0] in_read_valid_reg;
	reg [0:0] in_rst_reg;
	reg [0:0] in_write_valid_reg;

	assign valid = valid_reg;
	assign out_in_data = out_in_data_reg;
	assign out_read_valid = out_read_valid_reg;
	assign out_rst = out_rst_reg;
	assign out_write_valid = out_write_valid_reg;
	assign in_in_data = in_in_data_reg;
	assign in_read_valid = in_read_valid_reg;
	assign in_rst = in_rst_reg;
	assign in_write_valid = in_write_valid_reg;

	// Start debug wires and ports

	initial begin
	end





	// End debug wires and ports

	// Start Functional Units
	add alloca_0();

	add bitcast_1();

	add call_2();

	reg [31:0] raddr_ram_0_reg;
	reg [31:0] waddr_ram_0_reg;
	reg [31:0] wdata_ram_0_reg;
	reg [0:0] wen_ram_0_reg;
	wire [31:0] rdata_ram_0;
	register #(.WIDTH(32)) ram_0(.clk(clk), .raddr(raddr_ram_0_reg), .rdata(rdata_ram_0), .rst(rst), .waddr(waddr_ram_0_reg), .wdata(wdata_ram_0_reg), .wen(wen_ram_0_reg));

	br_dummy br_unit();

	add call_18();

	reg [63:0] phi_in_phi_5;
	reg [31:0] phi_last_block_phi_5;
	reg [63:0] phi_s_phi_5;
	wire [31:0] phi_out_phi_5;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_5(.in(phi_in_phi_5), .last_block(phi_last_block_phi_5), .out(phi_out_phi_5), .s(phi_s_phi_5));

	reg [31:0] add_in0_add_12;
	reg [31:0] add_in1_add_12;
	wire [31:0] add_out_add_12;
	add #(.WIDTH(32)) add_add_12(.in0(add_in0_add_12), .in1(add_in1_add_12), .out(add_out_add_12));

	reg [31:0] add_in0_add_14;
	reg [31:0] add_in1_add_14;
	wire [31:0] add_out_add_14;
	add #(.WIDTH(32)) add_add_14(.in0(add_in0_add_14), .in1(add_in1_add_14), .out(add_out_add_14));

	reg [31:0] cmp_in0_icmp_15;
	reg [31:0] cmp_in1_icmp_15;
	wire [0:0] cmp_out_icmp_15;
	eq #(.WIDTH(32)) icmp_15(.in0(cmp_in0_icmp_15), .in1(cmp_in1_icmp_15), .out(cmp_out_icmp_15));

	reg [31:0] data_in_1_1_in_data;
	wire [31:0] data_in_1_1_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_1(.in_data(data_in_1_1_in_data), .out_data(data_in_1_1_out_data));

	reg [31:0] data_in_1_3_in_data;
	wire [31:0] data_in_1_3_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_3(.in_data(data_in_1_3_in_data), .out_data(data_in_1_3_out_data));

	reg [0:0] data_in_1_5_in_data;
	wire [0:0] data_in_1_5_out_data;
	hls_wire #(.WIDTH(1)) data_in_1_5(.in_data(data_in_1_5_in_data), .out_data(data_in_1_5_out_data));

	reg [31:0] data_in_1_7_in_data;
	wire [31:0] data_in_1_7_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_7(.in_data(data_in_1_7_in_data), .out_data(data_in_1_7_out_data));

	reg [31:0] data_in_2_9_in_data;
	wire [31:0] data_in_2_9_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_9(.in_data(data_in_2_9_in_data), .out_data(data_in_2_9_out_data));

	reg [31:0] data_in_2_11_in_data;
	wire [31:0] data_in_2_11_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_11(.in_data(data_in_2_11_in_data), .out_data(data_in_2_11_out_data));

	reg [0:0] data_in_2_13_in_data;
	wire [0:0] data_in_2_13_out_data;
	hls_wire #(.WIDTH(1)) data_in_2_13(.in_data(data_in_2_13_in_data), .out_data(data_in_2_13_out_data));

	reg [31:0] data_in_2_15_in_data;
	wire [31:0] data_in_2_15_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_15(.in_data(data_in_2_15_in_data), .out_data(data_in_2_15_out_data));

	reg [31:0] data_in_3_17_in_data;
	wire [31:0] data_in_3_17_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_17(.in_data(data_in_3_17_in_data), .out_data(data_in_3_17_out_data));

	reg [31:0] data_in_3_19_in_data;
	wire [31:0] data_in_3_19_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_19(.in_data(data_in_3_19_in_data), .out_data(data_in_3_19_out_data));

	reg [0:0] data_in_3_21_in_data;
	wire [0:0] data_in_3_21_out_data;
	hls_wire #(.WIDTH(1)) data_in_3_21(.in_data(data_in_3_21_in_data), .out_data(data_in_3_21_out_data));

	reg [31:0] data_in_3_23_in_data;
	wire [31:0] data_in_3_23_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_23(.in_data(data_in_3_23_in_data), .out_data(data_in_3_23_out_data));

	reg [31:0] data_in_4_25_in_data;
	wire [31:0] data_in_4_25_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_25(.in_data(data_in_4_25_in_data), .out_data(data_in_4_25_out_data));

	reg [31:0] data_in_4_27_in_data;
	wire [31:0] data_in_4_27_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_27(.in_data(data_in_4_27_in_data), .out_data(data_in_4_27_out_data));

	reg [0:0] data_in_4_29_in_data;
	wire [0:0] data_in_4_29_out_data;
	hls_wire #(.WIDTH(1)) data_in_4_29(.in_data(data_in_4_29_in_data), .out_data(data_in_4_29_out_data));

	reg [31:0] data_in_4_31_in_data;
	wire [31:0] data_in_4_31_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_31(.in_data(data_in_4_31_in_data), .out_data(data_in_4_31_out_data));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] bb_0_active_in_state_1_in_data;
	wire [0:0] bb_0_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_1(.in_data(bb_0_active_in_state_1_in_data), .out_data(bb_0_active_in_state_1_out_data));

	reg [31:0] bb_0_predecessor_in_state_1_in_data;
	wire [31:0] bb_0_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_1(.in_data(bb_0_predecessor_in_state_1_in_data), .out_data(bb_0_predecessor_in_state_1_out_data));

	reg [0:0] bb_3_active_in_state_1_in_data;
	wire [0:0] bb_3_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_1(.in_data(bb_3_active_in_state_1_in_data), .out_data(bb_3_active_in_state_1_out_data));

	reg [31:0] bb_3_predecessor_in_state_1_in_data;
	wire [31:0] bb_3_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_1(.in_data(bb_3_predecessor_in_state_1_in_data), .out_data(bb_3_predecessor_in_state_1_out_data));

	reg [0:0] bb_9_active_in_state_1_in_data;
	wire [0:0] bb_9_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_9_active_in_state_1(.in_data(bb_9_active_in_state_1_in_data), .out_data(bb_9_active_in_state_1_out_data));

	reg [31:0] bb_9_predecessor_in_state_1_in_data;
	wire [31:0] bb_9_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_9_predecessor_in_state_1(.in_data(bb_9_predecessor_in_state_1_in_data), .out_data(bb_9_predecessor_in_state_1_out_data));

	reg [0:0] bb_8_active_in_state_1_in_data;
	wire [0:0] bb_8_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active_in_state_1(.in_data(bb_8_active_in_state_1_in_data), .out_data(bb_8_active_in_state_1_out_data));

	reg [31:0] bb_8_predecessor_in_state_1_in_data;
	wire [31:0] bb_8_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor_in_state_1(.in_data(bb_8_predecessor_in_state_1_in_data), .out_data(bb_8_predecessor_in_state_1_out_data));

	reg [0:0] bb_10_active_in_state_2_in_data;
	wire [0:0] bb_10_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_2(.in_data(bb_10_active_in_state_2_in_data), .out_data(bb_10_active_in_state_2_out_data));

	reg [31:0] bb_10_predecessor_in_state_2_in_data;
	wire [31:0] bb_10_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_2(.in_data(bb_10_predecessor_in_state_2_in_data), .out_data(bb_10_predecessor_in_state_2_out_data));

	reg [0:0] bb_10_active_in_state_3_in_data;
	wire [0:0] bb_10_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_3(.in_data(bb_10_active_in_state_3_in_data), .out_data(bb_10_active_in_state_3_out_data));

	reg [31:0] bb_10_predecessor_in_state_3_in_data;
	wire [31:0] bb_10_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_3(.in_data(bb_10_predecessor_in_state_3_in_data), .out_data(bb_10_predecessor_in_state_3_out_data));

	reg [0:0] bb_4_active_in_state_3_in_data;
	wire [0:0] bb_4_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_3(.in_data(bb_4_active_in_state_3_in_data), .out_data(bb_4_active_in_state_3_out_data));

	reg [31:0] bb_4_predecessor_in_state_3_in_data;
	wire [31:0] bb_4_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_3(.in_data(bb_4_predecessor_in_state_3_in_data), .out_data(bb_4_predecessor_in_state_3_out_data));

	reg [0:0] bb_1_active_in_state_4_in_data;
	wire [0:0] bb_1_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_4(.in_data(bb_1_active_in_state_4_in_data), .out_data(bb_1_active_in_state_4_out_data));

	reg [31:0] bb_1_predecessor_in_state_4_in_data;
	wire [31:0] bb_1_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_4(.in_data(bb_1_predecessor_in_state_4_in_data), .out_data(bb_1_predecessor_in_state_4_out_data));

	reg [0:0] bb_2_active_in_state_4_in_data;
	wire [0:0] bb_2_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_4(.in_data(bb_2_active_in_state_4_in_data), .out_data(bb_2_active_in_state_4_out_data));

	reg [31:0] bb_2_predecessor_in_state_4_in_data;
	wire [31:0] bb_2_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_4(.in_data(bb_2_predecessor_in_state_4_in_data), .out_data(bb_2_predecessor_in_state_4_out_data));

	reg [0:0] bb_5_active_in_state_4_in_data;
	wire [0:0] bb_5_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_5_active_in_state_4(.in_data(bb_5_active_in_state_4_in_data), .out_data(bb_5_active_in_state_4_out_data));

	reg [31:0] bb_5_predecessor_in_state_4_in_data;
	wire [31:0] bb_5_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_5_predecessor_in_state_4(.in_data(bb_5_predecessor_in_state_4_in_data), .out_data(bb_5_predecessor_in_state_4_out_data));

	reg [0:0] bb_6_active_in_state_4_in_data;
	wire [0:0] bb_6_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_6_active_in_state_4(.in_data(bb_6_active_in_state_4_in_data), .out_data(bb_6_active_in_state_4_out_data));

	reg [31:0] bb_6_predecessor_in_state_4_in_data;
	wire [31:0] bb_6_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_6_predecessor_in_state_4(.in_data(bb_6_predecessor_in_state_4_in_data), .out_data(bb_6_predecessor_in_state_4_out_data));

	reg [0:0] bb_7_active_in_state_4_in_data;
	wire [0:0] bb_7_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_7_active_in_state_4(.in_data(bb_7_active_in_state_4_in_data), .out_data(bb_7_active_in_state_4_out_data));

	reg [31:0] bb_7_predecessor_in_state_4_in_data;
	wire [31:0] bb_7_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_7_predecessor_in_state_4(.in_data(bb_7_predecessor_in_state_4_in_data), .out_data(bb_7_predecessor_in_state_4_out_data));

	reg [0:0] bb_4_active_in_state_4_in_data;
	wire [0:0] bb_4_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_4(.in_data(bb_4_active_in_state_4_in_data), .out_data(bb_4_active_in_state_4_out_data));

	reg [31:0] bb_4_predecessor_in_state_4_in_data;
	wire [31:0] bb_4_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_4(.in_data(bb_4_predecessor_in_state_4_in_data), .out_data(bb_4_predecessor_in_state_4_out_data));

	reg [0:0] andOp_32_in0;
	reg [0:0] andOp_32_in1;
	wire [0:0] andOp_32_out;
	andOp #(.WIDTH(1)) andOp_32(.in0(andOp_32_in0), .in1(andOp_32_in1), .out(andOp_32_out));

	reg [0:0] andOp_33_in0;
	reg [0:0] andOp_33_in1;
	wire [0:0] andOp_33_out;
	andOp #(.WIDTH(1)) andOp_33(.in0(andOp_33_in0), .in1(andOp_33_in1), .out(andOp_33_out));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] notOp_34_in0;
	wire [0:0] notOp_34_out;
	notOp #(.WIDTH(1)) notOp_34(.in(notOp_34_in0), .out(notOp_34_out));

	reg [0:0] andOp_35_in0;
	reg [0:0] andOp_35_in1;
	wire [0:0] andOp_35_out;
	andOp #(.WIDTH(1)) andOp_35(.in0(andOp_35_in0), .in1(andOp_35_in1), .out(andOp_35_out));

	reg [0:0] andOp_36_in0;
	reg [0:0] andOp_36_in1;
	wire [0:0] andOp_36_out;
	andOp #(.WIDTH(1)) andOp_36(.in0(andOp_36_in0), .in1(andOp_36_in1), .out(andOp_36_out));

	reg [0:0] br_0_happened_in_state_1_in_data;
	wire [0:0] br_0_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_1(.in_data(br_0_happened_in_state_1_in_data), .out_data(br_0_happened_in_state_1_out_data));

	reg [0:0] notOp_37_in0;
	wire [0:0] notOp_37_out;
	notOp #(.WIDTH(1)) notOp_37(.in(notOp_37_in0), .out(notOp_37_out));

	reg [0:0] andOp_38_in0;
	reg [0:0] andOp_38_in1;
	wire [0:0] andOp_38_out;
	andOp #(.WIDTH(1)) andOp_38(.in0(andOp_38_in0), .in1(andOp_38_in1), .out(andOp_38_out));

	reg [0:0] andOp_39_in0;
	reg [0:0] andOp_39_in1;
	wire [0:0] andOp_39_out;
	andOp #(.WIDTH(1)) andOp_39(.in0(andOp_39_in0), .in1(andOp_39_in1), .out(andOp_39_out));

	reg [0:0] br_3_happened_in_state_1_in_data;
	wire [0:0] br_3_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_1(.in_data(br_3_happened_in_state_1_in_data), .out_data(br_3_happened_in_state_1_out_data));

	reg [0:0] notOp_40_in0;
	wire [0:0] notOp_40_out;
	notOp #(.WIDTH(1)) notOp_40(.in(notOp_40_in0), .out(notOp_40_out));

	reg [0:0] andOp_41_in0;
	reg [0:0] andOp_41_in1;
	wire [0:0] andOp_41_out;
	andOp #(.WIDTH(1)) andOp_41(.in0(andOp_41_in0), .in1(andOp_41_in1), .out(andOp_41_out));

	reg [0:0] andOp_42_in0;
	reg [0:0] andOp_42_in1;
	wire [0:0] andOp_42_out;
	andOp #(.WIDTH(1)) andOp_42(.in0(andOp_42_in0), .in1(andOp_42_in1), .out(andOp_42_out));

	reg [0:0] br_9_happened_in_state_1_in_data;
	wire [0:0] br_9_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_9_happened_in_state_1(.in_data(br_9_happened_in_state_1_in_data), .out_data(br_9_happened_in_state_1_out_data));

	reg [0:0] notOp_43_in0;
	wire [0:0] notOp_43_out;
	notOp #(.WIDTH(1)) notOp_43(.in(notOp_43_in0), .out(notOp_43_out));

	reg [0:0] andOp_44_in0;
	reg [0:0] andOp_44_in1;
	wire [0:0] andOp_44_out;
	andOp #(.WIDTH(1)) andOp_44(.in0(andOp_44_in0), .in1(andOp_44_in1), .out(andOp_44_out));

	reg [0:0] notOp_45_in0;
	wire [0:0] notOp_45_out;
	notOp #(.WIDTH(1)) notOp_45(.in(notOp_45_in0), .out(notOp_45_out));

	reg [0:0] andOp_46_in0;
	reg [0:0] andOp_46_in1;
	wire [0:0] andOp_46_out;
	andOp #(.WIDTH(1)) andOp_46(.in0(andOp_46_in0), .in1(andOp_46_in1), .out(andOp_46_out));

	reg [0:0] andOp_47_in0;
	reg [0:0] andOp_47_in1;
	wire [0:0] andOp_47_out;
	andOp #(.WIDTH(1)) andOp_47(.in0(andOp_47_in0), .in1(andOp_47_in1), .out(andOp_47_out));

	reg [0:0] andOp_48_in0;
	reg [0:0] andOp_48_in1;
	wire [0:0] andOp_48_out;
	andOp #(.WIDTH(1)) andOp_48(.in0(andOp_48_in0), .in1(andOp_48_in1), .out(andOp_48_out));

	reg [0:0] br_8_happened_in_state_1_in_data;
	wire [0:0] br_8_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_8_happened_in_state_1(.in_data(br_8_happened_in_state_1_in_data), .out_data(br_8_happened_in_state_1_out_data));

	reg [0:0] notOp_49_in0;
	wire [0:0] notOp_49_out;
	notOp #(.WIDTH(1)) notOp_49(.in(notOp_49_in0), .out(notOp_49_out));

	reg [0:0] andOp_50_in0;
	reg [0:0] andOp_50_in1;
	wire [0:0] andOp_50_out;
	andOp #(.WIDTH(1)) andOp_50(.in0(andOp_50_in0), .in1(andOp_50_in1), .out(andOp_50_out));

	reg [0:0] andOp_51_in0;
	reg [0:0] andOp_51_in1;
	wire [0:0] andOp_51_out;
	andOp #(.WIDTH(1)) andOp_51(.in0(andOp_51_in0), .in1(andOp_51_in1), .out(andOp_51_out));

	reg [0:0] br_10_happened_in_state_2_in_data;
	wire [0:0] br_10_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_2(.in_data(br_10_happened_in_state_2_in_data), .out_data(br_10_happened_in_state_2_out_data));

	reg [0:0] notOp_52_in0;
	wire [0:0] notOp_52_out;
	notOp #(.WIDTH(1)) notOp_52(.in(notOp_52_in0), .out(notOp_52_out));

	reg [0:0] andOp_53_in0;
	reg [0:0] andOp_53_in1;
	wire [0:0] andOp_53_out;
	andOp #(.WIDTH(1)) andOp_53(.in0(andOp_53_in0), .in1(andOp_53_in1), .out(andOp_53_out));

	reg [0:0] andOp_54_in0;
	reg [0:0] andOp_54_in1;
	wire [0:0] andOp_54_out;
	andOp #(.WIDTH(1)) andOp_54(.in0(andOp_54_in0), .in1(andOp_54_in1), .out(andOp_54_out));

	reg [0:0] br_10_happened_in_state_3_in_data;
	wire [0:0] br_10_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_3(.in_data(br_10_happened_in_state_3_in_data), .out_data(br_10_happened_in_state_3_out_data));

	reg [0:0] notOp_55_in0;
	wire [0:0] notOp_55_out;
	notOp #(.WIDTH(1)) notOp_55(.in(notOp_55_in0), .out(notOp_55_out));

	reg [0:0] andOp_56_in0;
	reg [0:0] andOp_56_in1;
	wire [0:0] andOp_56_out;
	andOp #(.WIDTH(1)) andOp_56(.in0(andOp_56_in0), .in1(andOp_56_in1), .out(andOp_56_out));

	reg [0:0] andOp_57_in0;
	reg [0:0] andOp_57_in1;
	wire [0:0] andOp_57_out;
	andOp #(.WIDTH(1)) andOp_57(.in0(andOp_57_in0), .in1(andOp_57_in1), .out(andOp_57_out));

	reg [0:0] br_4_happened_in_state_3_in_data;
	wire [0:0] br_4_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_3(.in_data(br_4_happened_in_state_3_in_data), .out_data(br_4_happened_in_state_3_out_data));

	reg [0:0] notOp_58_in0;
	wire [0:0] notOp_58_out;
	notOp #(.WIDTH(1)) notOp_58(.in(notOp_58_in0), .out(notOp_58_out));

	reg [0:0] andOp_59_in0;
	reg [0:0] andOp_59_in1;
	wire [0:0] andOp_59_out;
	andOp #(.WIDTH(1)) andOp_59(.in0(andOp_59_in0), .in1(andOp_59_in1), .out(andOp_59_out));

	reg [0:0] notOp_60_in0;
	wire [0:0] notOp_60_out;
	notOp #(.WIDTH(1)) notOp_60(.in(notOp_60_in0), .out(notOp_60_out));

	reg [0:0] andOp_61_in0;
	reg [0:0] andOp_61_in1;
	wire [0:0] andOp_61_out;
	andOp #(.WIDTH(1)) andOp_61(.in0(andOp_61_in0), .in1(andOp_61_in1), .out(andOp_61_out));

	reg [0:0] andOp_62_in0;
	reg [0:0] andOp_62_in1;
	wire [0:0] andOp_62_out;
	andOp #(.WIDTH(1)) andOp_62(.in0(andOp_62_in0), .in1(andOp_62_in1), .out(andOp_62_out));

	reg [0:0] andOp_63_in0;
	reg [0:0] andOp_63_in1;
	wire [0:0] andOp_63_out;
	andOp #(.WIDTH(1)) andOp_63(.in0(andOp_63_in0), .in1(andOp_63_in1), .out(andOp_63_out));

	reg [0:0] br_1_happened_in_state_4_in_data;
	wire [0:0] br_1_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened_in_state_4(.in_data(br_1_happened_in_state_4_in_data), .out_data(br_1_happened_in_state_4_out_data));

	reg [0:0] notOp_64_in0;
	wire [0:0] notOp_64_out;
	notOp #(.WIDTH(1)) notOp_64(.in(notOp_64_in0), .out(notOp_64_out));

	reg [0:0] andOp_65_in0;
	reg [0:0] andOp_65_in1;
	wire [0:0] andOp_65_out;
	andOp #(.WIDTH(1)) andOp_65(.in0(andOp_65_in0), .in1(andOp_65_in1), .out(andOp_65_out));

	reg [0:0] andOp_66_in0;
	reg [0:0] andOp_66_in1;
	wire [0:0] andOp_66_out;
	andOp #(.WIDTH(1)) andOp_66(.in0(andOp_66_in0), .in1(andOp_66_in1), .out(andOp_66_out));

	reg [0:0] br_5_happened_in_state_4_in_data;
	wire [0:0] br_5_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_5_happened_in_state_4(.in_data(br_5_happened_in_state_4_in_data), .out_data(br_5_happened_in_state_4_out_data));

	reg [0:0] notOp_67_in0;
	wire [0:0] notOp_67_out;
	notOp #(.WIDTH(1)) notOp_67(.in(notOp_67_in0), .out(notOp_67_out));

	reg [0:0] andOp_68_in0;
	reg [0:0] andOp_68_in1;
	wire [0:0] andOp_68_out;
	andOp #(.WIDTH(1)) andOp_68(.in0(andOp_68_in0), .in1(andOp_68_in1), .out(andOp_68_out));

	reg [0:0] andOp_69_in0;
	reg [0:0] andOp_69_in1;
	wire [0:0] andOp_69_out;
	andOp #(.WIDTH(1)) andOp_69(.in0(andOp_69_in0), .in1(andOp_69_in1), .out(andOp_69_out));

	reg [0:0] br_6_happened_in_state_4_in_data;
	wire [0:0] br_6_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_6_happened_in_state_4(.in_data(br_6_happened_in_state_4_in_data), .out_data(br_6_happened_in_state_4_out_data));

	reg [0:0] notOp_70_in0;
	wire [0:0] notOp_70_out;
	notOp #(.WIDTH(1)) notOp_70(.in(notOp_70_in0), .out(notOp_70_out));

	reg [0:0] andOp_71_in0;
	reg [0:0] andOp_71_in1;
	wire [0:0] andOp_71_out;
	andOp #(.WIDTH(1)) andOp_71(.in0(andOp_71_in0), .in1(andOp_71_in1), .out(andOp_71_out));

	reg [0:0] notOp_72_in0;
	wire [0:0] notOp_72_out;
	notOp #(.WIDTH(1)) notOp_72(.in(notOp_72_in0), .out(notOp_72_out));

	reg [0:0] andOp_73_in0;
	reg [0:0] andOp_73_in1;
	wire [0:0] andOp_73_out;
	andOp #(.WIDTH(1)) andOp_73(.in0(andOp_73_in0), .in1(andOp_73_in1), .out(andOp_73_out));

	reg [0:0] andOp_74_in0;
	reg [0:0] andOp_74_in1;
	wire [0:0] andOp_74_out;
	andOp #(.WIDTH(1)) andOp_74(.in0(andOp_74_in0), .in1(andOp_74_in1), .out(andOp_74_out));

	reg [0:0] andOp_75_in0;
	reg [0:0] andOp_75_in1;
	wire [0:0] andOp_75_out;
	andOp #(.WIDTH(1)) andOp_75(.in0(andOp_75_in0), .in1(andOp_75_in1), .out(andOp_75_out));

	reg [0:0] br_7_happened_in_state_4_in_data;
	wire [0:0] br_7_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_7_happened_in_state_4(.in_data(br_7_happened_in_state_4_in_data), .out_data(br_7_happened_in_state_4_out_data));

	reg [0:0] notOp_76_in0;
	wire [0:0] notOp_76_out;
	notOp #(.WIDTH(1)) notOp_76(.in(notOp_76_in0), .out(notOp_76_out));

	reg [0:0] andOp_77_in0;
	reg [0:0] andOp_77_in1;
	wire [0:0] andOp_77_out;
	andOp #(.WIDTH(1)) andOp_77(.in0(andOp_77_in0), .in1(andOp_77_in1), .out(andOp_77_out));

	reg [0:0] andOp_78_in0;
	reg [0:0] andOp_78_in1;
	wire [0:0] andOp_78_out;
	andOp #(.WIDTH(1)) andOp_78(.in0(andOp_78_in0), .in1(andOp_78_in1), .out(andOp_78_out));

	reg [0:0] br_4_happened_in_state_4_in_data;
	wire [0:0] br_4_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_4(.in_data(br_4_happened_in_state_4_in_data), .out_data(br_4_happened_in_state_4_out_data));

	reg [0:0] notOp_79_in0;
	wire [0:0] notOp_79_out;
	notOp #(.WIDTH(1)) notOp_79(.in(notOp_79_in0), .out(notOp_79_out));

	reg [0:0] andOp_80_in0;
	reg [0:0] andOp_80_in1;
	wire [0:0] andOp_80_out;
	andOp #(.WIDTH(1)) andOp_80(.in0(andOp_80_in0), .in1(andOp_80_in1), .out(andOp_80_out));

	reg [0:0] notOp_81_in0;
	wire [0:0] notOp_81_out;
	notOp #(.WIDTH(1)) notOp_81(.in(notOp_81_in0), .out(notOp_81_out));

	reg [0:0] andOp_82_in0;
	reg [0:0] andOp_82_in1;
	wire [0:0] andOp_82_out;
	andOp #(.WIDTH(1)) andOp_82(.in0(andOp_82_in0), .in1(andOp_82_in1), .out(andOp_82_out));

	reg [31:0] eq_83_in0;
	reg [31:0] eq_83_in1;
	wire [0:0] eq_83_out;
	eq #(.WIDTH(32)) eq_83(.in0(eq_83_in0), .in1(eq_83_in1), .out(eq_83_out));

	reg [31:0] eq_84_in0;
	reg [31:0] eq_84_in1;
	wire [0:0] eq_84_out;
	eq #(.WIDTH(32)) eq_84(.in0(eq_84_in0), .in1(eq_84_in1), .out(eq_84_out));

	reg [31:0] eq_85_in0;
	reg [31:0] eq_85_in1;
	wire [0:0] eq_85_out;
	eq #(.WIDTH(32)) eq_85(.in0(eq_85_in0), .in1(eq_85_in1), .out(eq_85_out));

	reg [0:0] orOp_86_in0;
	reg [0:0] orOp_86_in1;
	wire [0:0] orOp_86_out;
	orOp #(.WIDTH(1)) orOp_86(.in0(orOp_86_in0), .in1(orOp_86_in1), .out(orOp_86_out));

	reg [31:0] eq_87_in0;
	reg [31:0] eq_87_in1;
	wire [0:0] eq_87_out;
	eq #(.WIDTH(32)) eq_87(.in0(eq_87_in0), .in1(eq_87_in1), .out(eq_87_out));

	reg [0:0] orOp_88_in0;
	reg [0:0] orOp_88_in1;
	wire [0:0] orOp_88_out;
	orOp #(.WIDTH(1)) orOp_88(.in0(orOp_88_in0), .in1(orOp_88_in1), .out(orOp_88_out));

	reg [31:0] eq_89_in0;
	reg [31:0] eq_89_in1;
	wire [0:0] eq_89_out;
	eq #(.WIDTH(32)) eq_89(.in0(eq_89_in0), .in1(eq_89_in1), .out(eq_89_out));

	reg [0:0] orOp_90_in0;
	reg [0:0] orOp_90_in1;
	wire [0:0] orOp_90_out;
	orOp #(.WIDTH(1)) orOp_90(.in0(orOp_90_in0), .in1(orOp_90_in1), .out(orOp_90_out));

	reg [31:0] eq_91_in0;
	reg [31:0] eq_91_in1;
	wire [0:0] eq_91_out;
	eq #(.WIDTH(32)) eq_91(.in0(eq_91_in0), .in1(eq_91_in1), .out(eq_91_out));

	reg [31:0] eq_92_in0;
	reg [31:0] eq_92_in1;
	wire [0:0] eq_92_out;
	eq #(.WIDTH(32)) eq_92(.in0(eq_92_in0), .in1(eq_92_in1), .out(eq_92_out));

	reg [31:0] eq_93_in0;
	reg [31:0] eq_93_in1;
	wire [0:0] eq_93_out;
	eq #(.WIDTH(32)) eq_93(.in0(eq_93_in0), .in1(eq_93_in1), .out(eq_93_out));

	reg [0:0] orOp_94_in0;
	reg [0:0] orOp_94_in1;
	wire [0:0] orOp_94_out;
	orOp #(.WIDTH(1)) orOp_94(.in0(orOp_94_in0), .in1(orOp_94_in1), .out(orOp_94_out));

	reg [31:0] eq_95_in0;
	reg [31:0] eq_95_in1;
	wire [0:0] eq_95_out;
	eq #(.WIDTH(32)) eq_95(.in0(eq_95_in0), .in1(eq_95_in1), .out(eq_95_out));

	reg [0:0] orOp_96_in0;
	reg [0:0] orOp_96_in1;
	wire [0:0] orOp_96_out;
	orOp #(.WIDTH(1)) orOp_96(.in0(orOp_96_in0), .in1(orOp_96_in1), .out(orOp_96_out));

	reg [31:0] eq_97_in0;
	reg [31:0] eq_97_in1;
	wire [0:0] eq_97_out;
	eq #(.WIDTH(32)) eq_97(.in0(eq_97_in0), .in1(eq_97_in1), .out(eq_97_out));

	reg [0:0] orOp_98_in0;
	reg [0:0] orOp_98_in1;
	wire [0:0] orOp_98_out;
	orOp #(.WIDTH(1)) orOp_98(.in0(orOp_98_in0), .in1(orOp_98_in1), .out(orOp_98_out));

	reg [31:0] eq_99_in0;
	reg [31:0] eq_99_in1;
	wire [0:0] eq_99_out;
	eq #(.WIDTH(32)) eq_99(.in0(eq_99_in0), .in1(eq_99_in1), .out(eq_99_out));

	reg [0:0] orOp_100_in0;
	reg [0:0] orOp_100_in1;
	wire [0:0] orOp_100_out;
	orOp #(.WIDTH(1)) orOp_100(.in0(orOp_100_in0), .in1(orOp_100_in1), .out(orOp_100_out));

	reg [31:0] eq_101_in0;
	reg [31:0] eq_101_in1;
	wire [0:0] eq_101_out;
	eq #(.WIDTH(32)) eq_101(.in0(eq_101_in0), .in1(eq_101_in1), .out(eq_101_out));

	reg [0:0] orOp_102_in0;
	reg [0:0] orOp_102_in1;
	wire [0:0] orOp_102_out;
	orOp #(.WIDTH(1)) orOp_102(.in0(orOp_102_in0), .in1(orOp_102_in1), .out(orOp_102_out));

	reg [31:0] eq_103_in0;
	reg [31:0] eq_103_in1;
	wire [0:0] eq_103_out;
	eq #(.WIDTH(32)) eq_103(.in0(eq_103_in0), .in1(eq_103_in1), .out(eq_103_out));

	reg [0:0] orOp_104_in0;
	reg [0:0] orOp_104_in1;
	wire [0:0] orOp_104_out;
	orOp #(.WIDTH(1)) orOp_104(.in0(orOp_104_in0), .in1(orOp_104_in1), .out(orOp_104_out));

	reg [31:0] eq_105_in0;
	reg [31:0] eq_105_in1;
	wire [0:0] eq_105_out;
	eq #(.WIDTH(32)) eq_105(.in0(eq_105_in0), .in1(eq_105_in1), .out(eq_105_out));

	reg [31:0] eq_106_in0;
	reg [31:0] eq_106_in1;
	wire [0:0] eq_106_out;
	eq #(.WIDTH(32)) eq_106(.in0(eq_106_in0), .in1(eq_106_in1), .out(eq_106_out));

	reg [31:0] eq_107_in0;
	reg [31:0] eq_107_in1;
	wire [0:0] eq_107_out;
	eq #(.WIDTH(32)) eq_107(.in0(eq_107_in0), .in1(eq_107_in1), .out(eq_107_out));

	reg [31:0] eq_108_in0;
	reg [31:0] eq_108_in1;
	wire [0:0] eq_108_out;
	eq #(.WIDTH(32)) eq_108(.in0(eq_108_in0), .in1(eq_108_in1), .out(eq_108_out));

	reg [0:0] notOp_109_in0;
	wire [0:0] notOp_109_out;
	notOp #(.WIDTH(1)) notOp_109(.in(notOp_109_in0), .out(notOp_109_out));

	reg [0:0] andOp_110_in0;
	reg [0:0] andOp_110_in1;
	wire [0:0] andOp_110_out;
	andOp #(.WIDTH(1)) andOp_110(.in0(andOp_110_in0), .in1(andOp_110_in1), .out(andOp_110_out));

	reg [31:0] eq_111_in0;
	reg [31:0] eq_111_in1;
	wire [0:0] eq_111_out;
	eq #(.WIDTH(32)) eq_111(.in0(eq_111_in0), .in1(eq_111_in1), .out(eq_111_out));

	reg [0:0] notOp_112_in0;
	wire [0:0] notOp_112_out;
	notOp #(.WIDTH(1)) notOp_112(.in(notOp_112_in0), .out(notOp_112_out));

	reg [0:0] andOp_113_in0;
	reg [0:0] andOp_113_in1;
	wire [0:0] andOp_113_out;
	andOp #(.WIDTH(1)) andOp_113(.in0(andOp_113_in0), .in1(andOp_113_in1), .out(andOp_113_out));

	reg [31:0] eq_114_in0;
	reg [31:0] eq_114_in1;
	wire [0:0] eq_114_out;
	eq #(.WIDTH(32)) eq_114(.in0(eq_114_in0), .in1(eq_114_in1), .out(eq_114_out));

	reg [0:0] notOp_115_in0;
	wire [0:0] notOp_115_out;
	notOp #(.WIDTH(1)) notOp_115(.in(notOp_115_in0), .out(notOp_115_out));

	reg [0:0] andOp_116_in0;
	reg [0:0] andOp_116_in1;
	wire [0:0] andOp_116_out;
	andOp #(.WIDTH(1)) andOp_116(.in0(andOp_116_in0), .in1(andOp_116_in1), .out(andOp_116_out));

	reg [31:0] eq_117_in0;
	reg [31:0] eq_117_in1;
	wire [0:0] eq_117_out;
	eq #(.WIDTH(32)) eq_117(.in0(eq_117_in0), .in1(eq_117_in1), .out(eq_117_out));

	reg [31:0] eq_118_in0;
	reg [31:0] eq_118_in1;
	wire [0:0] eq_118_out;
	eq #(.WIDTH(32)) eq_118(.in0(eq_118_in0), .in1(eq_118_in1), .out(eq_118_out));

	reg [31:0] eq_119_in0;
	reg [31:0] eq_119_in1;
	wire [0:0] eq_119_out;
	eq #(.WIDTH(32)) eq_119(.in0(eq_119_in0), .in1(eq_119_in1), .out(eq_119_out));

	reg [0:0] notOp_120_in0;
	wire [0:0] notOp_120_out;
	notOp #(.WIDTH(1)) notOp_120(.in(notOp_120_in0), .out(notOp_120_out));

	reg [0:0] andOp_121_in0;
	reg [0:0] andOp_121_in1;
	wire [0:0] andOp_121_out;
	andOp #(.WIDTH(1)) andOp_121(.in0(andOp_121_in0), .in1(andOp_121_in1), .out(andOp_121_out));

	reg [31:0] eq_122_in0;
	reg [31:0] eq_122_in1;
	wire [0:0] eq_122_out;
	eq #(.WIDTH(32)) eq_122(.in0(eq_122_in0), .in1(eq_122_in1), .out(eq_122_out));

	reg [0:0] notOp_123_in0;
	wire [0:0] notOp_123_out;
	notOp #(.WIDTH(1)) notOp_123(.in(notOp_123_in0), .out(notOp_123_out));

	reg [0:0] andOp_124_in0;
	reg [0:0] andOp_124_in1;
	wire [0:0] andOp_124_out;
	andOp #(.WIDTH(1)) andOp_124(.in0(andOp_124_in0), .in1(andOp_124_in1), .out(andOp_124_out));

	reg [31:0] eq_125_in0;
	reg [31:0] eq_125_in1;
	wire [0:0] eq_125_out;
	eq #(.WIDTH(32)) eq_125(.in0(eq_125_in0), .in1(eq_125_in1), .out(eq_125_out));

	reg [0:0] notOp_126_in0;
	wire [0:0] notOp_126_out;
	notOp #(.WIDTH(1)) notOp_126(.in(notOp_126_in0), .out(notOp_126_out));

	reg [0:0] andOp_127_in0;
	reg [0:0] andOp_127_in1;
	wire [0:0] andOp_127_out;
	andOp #(.WIDTH(1)) andOp_127(.in0(andOp_127_in0), .in1(andOp_127_in1), .out(andOp_127_out));

	reg [31:0] eq_128_in0;
	reg [31:0] eq_128_in1;
	wire [0:0] eq_128_out;
	eq #(.WIDTH(32)) eq_128(.in0(eq_128_in0), .in1(eq_128_in1), .out(eq_128_out));

	reg [0:0] notOp_129_in0;
	wire [0:0] notOp_129_out;
	notOp #(.WIDTH(1)) notOp_129(.in(notOp_129_in0), .out(notOp_129_out));

	reg [0:0] andOp_130_in0;
	reg [0:0] andOp_130_in1;
	wire [0:0] andOp_130_out;
	andOp #(.WIDTH(1)) andOp_130(.in0(andOp_130_in0), .in1(andOp_130_in1), .out(andOp_130_out));

	reg [31:0] eq_131_in0;
	reg [31:0] eq_131_in1;
	wire [0:0] eq_131_out;
	eq #(.WIDTH(32)) eq_131(.in0(eq_131_in0), .in1(eq_131_in1), .out(eq_131_out));

	reg [0:0] notOp_132_in0;
	wire [0:0] notOp_132_out;
	notOp #(.WIDTH(1)) notOp_132(.in(notOp_132_in0), .out(notOp_132_out));

	reg [0:0] andOp_133_in0;
	reg [0:0] andOp_133_in1;
	wire [0:0] andOp_133_out;
	andOp #(.WIDTH(1)) andOp_133(.in0(andOp_133_in0), .in1(andOp_133_in1), .out(andOp_133_out));

	reg [31:0] eq_134_in0;
	reg [31:0] eq_134_in1;
	wire [0:0] eq_134_out;
	eq #(.WIDTH(32)) eq_134(.in0(eq_134_in0), .in1(eq_134_in1), .out(eq_134_out));

	reg [0:0] notOp_135_in0;
	wire [0:0] notOp_135_out;
	notOp #(.WIDTH(1)) notOp_135(.in(notOp_135_in0), .out(notOp_135_out));

	reg [0:0] andOp_136_in0;
	reg [0:0] andOp_136_in1;
	wire [0:0] andOp_136_out;
	andOp #(.WIDTH(1)) andOp_136(.in0(andOp_136_in0), .in1(andOp_136_in1), .out(andOp_136_out));

	reg [31:0] eq_137_in0;
	reg [31:0] eq_137_in1;
	wire [0:0] eq_137_out;
	eq #(.WIDTH(32)) eq_137(.in0(eq_137_in0), .in1(eq_137_in1), .out(eq_137_out));

	reg [0:0] andOp_138_in0;
	reg [0:0] andOp_138_in1;
	wire [0:0] andOp_138_out;
	andOp #(.WIDTH(1)) andOp_138(.in0(andOp_138_in0), .in1(andOp_138_in1), .out(andOp_138_out));

	reg [0:0] andOp_139_in0;
	reg [0:0] andOp_139_in1;
	wire [0:0] andOp_139_out;
	andOp #(.WIDTH(1)) andOp_139(.in0(andOp_139_in0), .in1(andOp_139_in1), .out(andOp_139_out));

	reg [0:0] andOp_140_in0;
	reg [0:0] andOp_140_in1;
	wire [0:0] andOp_140_out;
	andOp #(.WIDTH(1)) andOp_140(.in0(andOp_140_in0), .in1(andOp_140_in1), .out(andOp_140_out));

	reg [0:0] andOp_141_in0;
	reg [0:0] andOp_141_in1;
	wire [0:0] andOp_141_out;
	andOp #(.WIDTH(1)) andOp_141(.in0(andOp_141_in0), .in1(andOp_141_in1), .out(andOp_141_out));

	reg [0:0] andOp_142_in0;
	reg [0:0] andOp_142_in1;
	wire [0:0] andOp_142_out;
	andOp #(.WIDTH(1)) andOp_142(.in0(andOp_142_in0), .in1(andOp_142_in1), .out(andOp_142_out));

	reg [0:0] andOp_143_in0;
	reg [0:0] andOp_143_in1;
	wire [0:0] andOp_143_out;
	andOp #(.WIDTH(1)) andOp_143(.in0(andOp_143_in0), .in1(andOp_143_in1), .out(andOp_143_out));

	reg [0:0] andOp_144_in0;
	reg [0:0] andOp_144_in1;
	wire [0:0] andOp_144_out;
	andOp #(.WIDTH(1)) andOp_144(.in0(andOp_144_in0), .in1(andOp_144_in1), .out(andOp_144_out));

	reg [0:0] andOp_145_in0;
	reg [0:0] andOp_145_in1;
	wire [0:0] andOp_145_out;
	andOp #(.WIDTH(1)) andOp_145(.in0(andOp_145_in0), .in1(andOp_145_in1), .out(andOp_145_out));

	reg [31:0] concat_146_in0;
	reg [31:0] concat_146_in1;
	wire [63:0] concat_146_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_146(.in0(concat_146_in0), .in1(concat_146_in1), .out(concat_146_out));

	reg [31:0] concat_147_in0;
	reg [31:0] concat_147_in1;
	wire [63:0] concat_147_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_147(.in0(concat_147_in0), .in1(concat_147_in1), .out(concat_147_out));

	reg [0:0] andOp_148_in0;
	reg [0:0] andOp_148_in1;
	wire [0:0] andOp_148_out;
	andOp #(.WIDTH(1)) andOp_148(.in0(andOp_148_in0), .in1(andOp_148_in1), .out(andOp_148_out));

	reg [0:0] andOp_149_in0;
	reg [0:0] andOp_149_in1;
	wire [0:0] andOp_149_out;
	andOp #(.WIDTH(1)) andOp_149(.in0(andOp_149_in0), .in1(andOp_149_in1), .out(andOp_149_out));

	reg [0:0] andOp_150_in0;
	reg [0:0] andOp_150_in1;
	wire [0:0] andOp_150_out;
	andOp #(.WIDTH(1)) andOp_150(.in0(andOp_150_in0), .in1(andOp_150_in1), .out(andOp_150_out));

	reg [0:0] andOp_151_in0;
	reg [0:0] andOp_151_in1;
	wire [0:0] andOp_151_out;
	andOp #(.WIDTH(1)) andOp_151(.in0(andOp_151_in0), .in1(andOp_151_in1), .out(andOp_151_out));

	reg [31:0] tmp_output_152_in_data;
	wire [31:0] tmp_output_152_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_152(.in_data(tmp_output_152_in_data), .out_data(tmp_output_152_out_data));

	reg [31:0] eq_153_in0;
	reg [31:0] eq_153_in1;
	wire [0:0] eq_153_out;
	eq #(.WIDTH(32)) eq_153(.in0(eq_153_in0), .in1(eq_153_in1), .out(eq_153_out));

	reg [0:0] andOp_154_in0;
	reg [0:0] andOp_154_in1;
	wire [0:0] andOp_154_out;
	andOp #(.WIDTH(1)) andOp_154(.in0(andOp_154_in0), .in1(andOp_154_in1), .out(andOp_154_out));

	reg [0:0] andOp_155_in0;
	reg [0:0] andOp_155_in1;
	wire [0:0] andOp_155_out;
	andOp #(.WIDTH(1)) andOp_155(.in0(andOp_155_in0), .in1(andOp_155_in1), .out(andOp_155_out));

	reg [0:0] andOp_156_in0;
	reg [0:0] andOp_156_in1;
	wire [0:0] andOp_156_out;
	andOp #(.WIDTH(1)) andOp_156(.in0(andOp_156_in0), .in1(andOp_156_in1), .out(andOp_156_out));

	reg [0:0] andOp_157_in0;
	reg [0:0] andOp_157_in1;
	wire [0:0] andOp_157_out;
	andOp #(.WIDTH(1)) andOp_157(.in0(andOp_157_in0), .in1(andOp_157_in1), .out(andOp_157_out));

	reg [0:0] andOp_158_in0;
	reg [0:0] andOp_158_in1;
	wire [0:0] andOp_158_out;
	andOp #(.WIDTH(1)) andOp_158(.in0(andOp_158_in0), .in1(andOp_158_in1), .out(andOp_158_out));

	reg [0:0] andOp_159_in0;
	reg [0:0] andOp_159_in1;
	wire [0:0] andOp_159_out;
	andOp #(.WIDTH(1)) andOp_159(.in0(andOp_159_in0), .in1(andOp_159_in1), .out(andOp_159_out));

	reg [0:0] andOp_160_in0;
	reg [0:0] andOp_160_in1;
	wire [0:0] andOp_160_out;
	andOp #(.WIDTH(1)) andOp_160(.in0(andOp_160_in0), .in1(andOp_160_in1), .out(andOp_160_out));

	reg [0:0] andOp_161_in0;
	reg [0:0] andOp_161_in1;
	wire [0:0] andOp_161_out;
	andOp #(.WIDTH(1)) andOp_161(.in0(andOp_161_in0), .in1(andOp_161_in1), .out(andOp_161_out));

	reg [0:0] andOp_162_in0;
	reg [0:0] andOp_162_in1;
	wire [0:0] andOp_162_out;
	andOp #(.WIDTH(1)) andOp_162(.in0(andOp_162_in0), .in1(andOp_162_in1), .out(andOp_162_out));

	reg [0:0] andOp_163_in0;
	reg [0:0] andOp_163_in1;
	wire [0:0] andOp_163_out;
	andOp #(.WIDTH(1)) andOp_163(.in0(andOp_163_in0), .in1(andOp_163_in1), .out(andOp_163_out));

	reg [0:0] andOp_164_in0;
	reg [0:0] andOp_164_in1;
	wire [0:0] andOp_164_out;
	andOp #(.WIDTH(1)) andOp_164(.in0(andOp_164_in0), .in1(andOp_164_in1), .out(andOp_164_out));

	reg [0:0] notOp_165_in0;
	wire [0:0] notOp_165_out;
	notOp #(.WIDTH(1)) notOp_165(.in(notOp_165_in0), .out(notOp_165_out));

	reg [0:0] andOp_166_in0;
	reg [0:0] andOp_166_in1;
	wire [0:0] andOp_166_out;
	andOp #(.WIDTH(1)) andOp_166(.in0(andOp_166_in0), .in1(andOp_166_in1), .out(andOp_166_out));

	reg [0:0] notOp_167_in0;
	wire [0:0] notOp_167_out;
	notOp #(.WIDTH(1)) notOp_167(.in(notOp_167_in0), .out(notOp_167_out));

	reg [0:0] andOp_168_in0;
	reg [0:0] andOp_168_in1;
	wire [0:0] andOp_168_out;
	andOp #(.WIDTH(1)) andOp_168(.in0(andOp_168_in0), .in1(andOp_168_in1), .out(andOp_168_out));

	reg [0:0] notOp_169_in0;
	wire [0:0] notOp_169_out;
	notOp #(.WIDTH(1)) notOp_169(.in(notOp_169_in0), .out(notOp_169_out));

	reg [0:0] andOp_170_in0;
	reg [0:0] andOp_170_in1;
	wire [0:0] andOp_170_out;
	andOp #(.WIDTH(1)) andOp_170(.in0(andOp_170_in0), .in1(andOp_170_in1), .out(andOp_170_out));

	reg [0:0] notOp_171_in0;
	wire [0:0] notOp_171_out;
	notOp #(.WIDTH(1)) notOp_171(.in(notOp_171_in0), .out(notOp_171_out));

	reg [0:0] andOp_172_in0;
	reg [0:0] andOp_172_in1;
	wire [0:0] andOp_172_out;
	andOp #(.WIDTH(1)) andOp_172(.in0(andOp_172_in0), .in1(andOp_172_in1), .out(andOp_172_out));

	reg [0:0] notOp_173_in0;
	wire [0:0] notOp_173_out;
	notOp #(.WIDTH(1)) notOp_173(.in(notOp_173_in0), .out(notOp_173_out));

	reg [0:0] andOp_174_in0;
	reg [0:0] andOp_174_in1;
	wire [0:0] andOp_174_out;
	andOp #(.WIDTH(1)) andOp_174(.in0(andOp_174_in0), .in1(andOp_174_in1), .out(andOp_174_out));

	reg [0:0] notOp_175_in0;
	wire [0:0] notOp_175_out;
	notOp #(.WIDTH(1)) notOp_175(.in(notOp_175_in0), .out(notOp_175_out));

	reg [0:0] andOp_176_in0;
	reg [0:0] andOp_176_in1;
	wire [0:0] andOp_176_out;
	andOp #(.WIDTH(1)) andOp_176(.in0(andOp_176_in0), .in1(andOp_176_in1), .out(andOp_176_out));

	reg [0:0] notOp_177_in0;
	wire [0:0] notOp_177_out;
	notOp #(.WIDTH(1)) notOp_177(.in(notOp_177_in0), .out(notOp_177_out));

	reg [0:0] andOp_178_in0;
	reg [0:0] andOp_178_in1;
	wire [0:0] andOp_178_out;
	andOp #(.WIDTH(1)) andOp_178(.in0(andOp_178_in0), .in1(andOp_178_in1), .out(andOp_178_out));

	reg [0:0] notOp_179_in0;
	wire [0:0] notOp_179_out;
	notOp #(.WIDTH(1)) notOp_179(.in(notOp_179_in0), .out(notOp_179_out));

	reg [0:0] andOp_180_in0;
	reg [0:0] andOp_180_in1;
	wire [0:0] andOp_180_out;
	andOp #(.WIDTH(1)) andOp_180(.in0(andOp_180_in0), .in1(andOp_180_in1), .out(andOp_180_out));

	reg [31:0] eq_181_in0;
	reg [31:0] eq_181_in1;
	wire [0:0] eq_181_out;
	eq #(.WIDTH(32)) eq_181(.in0(eq_181_in0), .in1(eq_181_in1), .out(eq_181_out));

	reg [31:0] eq_182_in0;
	reg [31:0] eq_182_in1;
	wire [0:0] eq_182_out;
	eq #(.WIDTH(32)) eq_182(.in0(eq_182_in0), .in1(eq_182_in1), .out(eq_182_out));

	reg [31:0] eq_183_in0;
	reg [31:0] eq_183_in1;
	wire [0:0] eq_183_out;
	eq #(.WIDTH(32)) eq_183(.in0(eq_183_in0), .in1(eq_183_in1), .out(eq_183_out));

	reg [31:0] eq_184_in0;
	reg [31:0] eq_184_in1;
	wire [0:0] eq_184_out;
	eq #(.WIDTH(32)) eq_184(.in0(eq_184_in0), .in1(eq_184_in1), .out(eq_184_out));

	reg [0:0] andOp_185_in0;
	reg [0:0] andOp_185_in1;
	wire [0:0] andOp_185_out;
	andOp #(.WIDTH(1)) andOp_185(.in0(andOp_185_in0), .in1(andOp_185_in1), .out(andOp_185_out));

	reg [31:0] eq_186_in0;
	reg [31:0] eq_186_in1;
	wire [0:0] eq_186_out;
	eq #(.WIDTH(32)) eq_186(.in0(eq_186_in0), .in1(eq_186_in1), .out(eq_186_out));

	reg [0:0] andOp_187_in0;
	reg [0:0] andOp_187_in1;
	wire [0:0] andOp_187_out;
	andOp #(.WIDTH(1)) andOp_187(.in0(andOp_187_in0), .in1(andOp_187_in1), .out(andOp_187_out));

	reg [0:0] notOp_188_in0;
	wire [0:0] notOp_188_out;
	notOp #(.WIDTH(1)) notOp_188(.in(notOp_188_in0), .out(notOp_188_out));

	reg [0:0] andOp_189_in0;
	reg [0:0] andOp_189_in1;
	wire [0:0] andOp_189_out;
	andOp #(.WIDTH(1)) andOp_189(.in0(andOp_189_in0), .in1(andOp_189_in1), .out(andOp_189_out));

	reg [0:0] notOp_190_in0;
	wire [0:0] notOp_190_out;
	notOp #(.WIDTH(1)) notOp_190(.in(notOp_190_in0), .out(notOp_190_out));

	reg [0:0] andOp_191_in0;
	reg [0:0] andOp_191_in1;
	wire [0:0] andOp_191_out;
	andOp #(.WIDTH(1)) andOp_191(.in0(andOp_191_in0), .in1(andOp_191_in1), .out(andOp_191_out));

	reg [0:0] notOp_192_in0;
	wire [0:0] notOp_192_out;
	notOp #(.WIDTH(1)) notOp_192(.in(notOp_192_in0), .out(notOp_192_out));

	reg [0:0] andOp_193_in0;
	reg [0:0] andOp_193_in1;
	wire [0:0] andOp_193_out;
	andOp #(.WIDTH(1)) andOp_193(.in0(andOp_193_in0), .in1(andOp_193_in1), .out(andOp_193_out));

	reg [0:0] andOp_194_in0;
	reg [0:0] andOp_194_in1;
	wire [0:0] andOp_194_out;
	andOp #(.WIDTH(1)) andOp_194(.in0(andOp_194_in0), .in1(andOp_194_in1), .out(andOp_194_out));

	reg [31:0] eq_195_in0;
	reg [31:0] eq_195_in1;
	wire [0:0] eq_195_out;
	eq #(.WIDTH(32)) eq_195(.in0(eq_195_in0), .in1(eq_195_in1), .out(eq_195_out));

	reg [0:0] andOp_196_in0;
	reg [0:0] andOp_196_in1;
	wire [0:0] andOp_196_out;
	andOp #(.WIDTH(1)) andOp_196(.in0(andOp_196_in0), .in1(andOp_196_in1), .out(andOp_196_out));

	reg [0:0] notOp_197_in0;
	wire [0:0] notOp_197_out;
	notOp #(.WIDTH(1)) notOp_197(.in(notOp_197_in0), .out(notOp_197_out));

	reg [0:0] andOp_198_in0;
	reg [0:0] andOp_198_in1;
	wire [0:0] andOp_198_out;
	andOp #(.WIDTH(1)) andOp_198(.in0(andOp_198_in0), .in1(andOp_198_in1), .out(andOp_198_out));

	reg [0:0] notOp_199_in0;
	wire [0:0] notOp_199_out;
	notOp #(.WIDTH(1)) notOp_199(.in(notOp_199_in0), .out(notOp_199_out));

	reg [0:0] andOp_200_in0;
	reg [0:0] andOp_200_in1;
	wire [0:0] andOp_200_out;
	andOp #(.WIDTH(1)) andOp_200(.in0(andOp_200_in0), .in1(andOp_200_in1), .out(andOp_200_out));

	reg [0:0] notOp_201_in0;
	wire [0:0] notOp_201_out;
	notOp #(.WIDTH(1)) notOp_201(.in(notOp_201_in0), .out(notOp_201_out));

	reg [0:0] andOp_202_in0;
	reg [0:0] andOp_202_in1;
	wire [0:0] andOp_202_out;
	andOp #(.WIDTH(1)) andOp_202(.in0(andOp_202_in0), .in1(andOp_202_in1), .out(andOp_202_out));

	reg [0:0] andOp_203_in0;
	reg [0:0] andOp_203_in1;
	wire [0:0] andOp_203_out;
	andOp #(.WIDTH(1)) andOp_203(.in0(andOp_203_in0), .in1(andOp_203_in1), .out(andOp_203_out));

	reg [31:0] eq_204_in0;
	reg [31:0] eq_204_in1;
	wire [0:0] eq_204_out;
	eq #(.WIDTH(32)) eq_204(.in0(eq_204_in0), .in1(eq_204_in1), .out(eq_204_out));

	reg [0:0] andOp_205_in0;
	reg [0:0] andOp_205_in1;
	wire [0:0] andOp_205_out;
	andOp #(.WIDTH(1)) andOp_205(.in0(andOp_205_in0), .in1(andOp_205_in1), .out(andOp_205_out));

	reg [0:0] notOp_206_in0;
	wire [0:0] notOp_206_out;
	notOp #(.WIDTH(1)) notOp_206(.in(notOp_206_in0), .out(notOp_206_out));

	reg [0:0] andOp_207_in0;
	reg [0:0] andOp_207_in1;
	wire [0:0] andOp_207_out;
	andOp #(.WIDTH(1)) andOp_207(.in0(andOp_207_in0), .in1(andOp_207_in1), .out(andOp_207_out));

	reg [0:0] notOp_208_in0;
	wire [0:0] notOp_208_out;
	notOp #(.WIDTH(1)) notOp_208(.in(notOp_208_in0), .out(notOp_208_out));

	reg [0:0] andOp_209_in0;
	reg [0:0] andOp_209_in1;
	wire [0:0] andOp_209_out;
	andOp #(.WIDTH(1)) andOp_209(.in0(andOp_209_in0), .in1(andOp_209_in1), .out(andOp_209_out));

	reg [0:0] notOp_210_in0;
	wire [0:0] notOp_210_out;
	notOp #(.WIDTH(1)) notOp_210(.in(notOp_210_in0), .out(notOp_210_out));

	reg [0:0] andOp_211_in0;
	reg [0:0] andOp_211_in1;
	wire [0:0] andOp_211_out;
	andOp #(.WIDTH(1)) andOp_211(.in0(andOp_211_in0), .in1(andOp_211_in1), .out(andOp_211_out));

	reg [0:0] andOp_212_in0;
	reg [0:0] andOp_212_in1;
	wire [0:0] andOp_212_out;
	andOp #(.WIDTH(1)) andOp_212(.in0(andOp_212_in0), .in1(andOp_212_in1), .out(andOp_212_out));

	reg [31:0] eq_213_in0;
	reg [31:0] eq_213_in1;
	wire [0:0] eq_213_out;
	eq #(.WIDTH(32)) eq_213(.in0(eq_213_in0), .in1(eq_213_in1), .out(eq_213_out));

	reg [0:0] andOp_214_in0;
	reg [0:0] andOp_214_in1;
	wire [0:0] andOp_214_out;
	andOp #(.WIDTH(1)) andOp_214(.in0(andOp_214_in0), .in1(andOp_214_in1), .out(andOp_214_out));

	reg [0:0] notOp_215_in0;
	wire [0:0] notOp_215_out;
	notOp #(.WIDTH(1)) notOp_215(.in(notOp_215_in0), .out(notOp_215_out));

	reg [0:0] andOp_216_in0;
	reg [0:0] andOp_216_in1;
	wire [0:0] andOp_216_out;
	andOp #(.WIDTH(1)) andOp_216(.in0(andOp_216_in0), .in1(andOp_216_in1), .out(andOp_216_out));

	reg [0:0] notOp_217_in0;
	wire [0:0] notOp_217_out;
	notOp #(.WIDTH(1)) notOp_217(.in(notOp_217_in0), .out(notOp_217_out));

	reg [0:0] andOp_218_in0;
	reg [0:0] andOp_218_in1;
	wire [0:0] andOp_218_out;
	andOp #(.WIDTH(1)) andOp_218(.in0(andOp_218_in0), .in1(andOp_218_in1), .out(andOp_218_out));

	reg [0:0] notOp_219_in0;
	wire [0:0] notOp_219_out;
	notOp #(.WIDTH(1)) notOp_219(.in(notOp_219_in0), .out(notOp_219_out));

	reg [0:0] andOp_220_in0;
	reg [0:0] andOp_220_in1;
	wire [0:0] andOp_220_out;
	andOp #(.WIDTH(1)) andOp_220(.in0(andOp_220_in0), .in1(andOp_220_in1), .out(andOp_220_out));

	reg [31:0] eq_221_in0;
	reg [31:0] eq_221_in1;
	wire [0:0] eq_221_out;
	eq #(.WIDTH(32)) eq_221(.in0(eq_221_in0), .in1(eq_221_in1), .out(eq_221_out));

	reg [31:0] eq_222_in0;
	reg [31:0] eq_222_in1;
	wire [0:0] eq_222_out;
	eq #(.WIDTH(32)) eq_222(.in0(eq_222_in0), .in1(eq_222_in1), .out(eq_222_out));

	reg [0:0] andOp_223_in0;
	reg [0:0] andOp_223_in1;
	wire [0:0] andOp_223_out;
	andOp #(.WIDTH(1)) andOp_223(.in0(andOp_223_in0), .in1(andOp_223_in1), .out(andOp_223_out));

	reg [31:0] eq_224_in0;
	reg [31:0] eq_224_in1;
	wire [0:0] eq_224_out;
	eq #(.WIDTH(32)) eq_224(.in0(eq_224_in0), .in1(eq_224_in1), .out(eq_224_out));

	reg [0:0] andOp_225_in0;
	reg [0:0] andOp_225_in1;
	wire [0:0] andOp_225_out;
	andOp #(.WIDTH(1)) andOp_225(.in0(andOp_225_in0), .in1(andOp_225_in1), .out(andOp_225_out));

	reg [0:0] notOp_226_in0;
	wire [0:0] notOp_226_out;
	notOp #(.WIDTH(1)) notOp_226(.in(notOp_226_in0), .out(notOp_226_out));

	reg [0:0] andOp_227_in0;
	reg [0:0] andOp_227_in1;
	wire [0:0] andOp_227_out;
	andOp #(.WIDTH(1)) andOp_227(.in0(andOp_227_in0), .in1(andOp_227_in1), .out(andOp_227_out));

	reg [0:0] notOp_228_in0;
	wire [0:0] notOp_228_out;
	notOp #(.WIDTH(1)) notOp_228(.in(notOp_228_in0), .out(notOp_228_out));

	reg [0:0] andOp_229_in0;
	reg [0:0] andOp_229_in1;
	wire [0:0] andOp_229_out;
	andOp #(.WIDTH(1)) andOp_229(.in0(andOp_229_in0), .in1(andOp_229_in1), .out(andOp_229_out));

	reg [0:0] notOp_230_in0;
	wire [0:0] notOp_230_out;
	notOp #(.WIDTH(1)) notOp_230(.in(notOp_230_in0), .out(notOp_230_out));

	reg [0:0] andOp_231_in0;
	reg [0:0] andOp_231_in1;
	wire [0:0] andOp_231_out;
	andOp #(.WIDTH(1)) andOp_231(.in0(andOp_231_in0), .in1(andOp_231_in1), .out(andOp_231_out));

	reg [0:0] andOp_232_in0;
	reg [0:0] andOp_232_in1;
	wire [0:0] andOp_232_out;
	andOp #(.WIDTH(1)) andOp_232(.in0(andOp_232_in0), .in1(andOp_232_in1), .out(andOp_232_out));

	reg [31:0] eq_233_in0;
	reg [31:0] eq_233_in1;
	wire [0:0] eq_233_out;
	eq #(.WIDTH(32)) eq_233(.in0(eq_233_in0), .in1(eq_233_in1), .out(eq_233_out));

	reg [0:0] andOp_234_in0;
	reg [0:0] andOp_234_in1;
	wire [0:0] andOp_234_out;
	andOp #(.WIDTH(1)) andOp_234(.in0(andOp_234_in0), .in1(andOp_234_in1), .out(andOp_234_out));

	reg [0:0] notOp_235_in0;
	wire [0:0] notOp_235_out;
	notOp #(.WIDTH(1)) notOp_235(.in(notOp_235_in0), .out(notOp_235_out));

	reg [0:0] andOp_236_in0;
	reg [0:0] andOp_236_in1;
	wire [0:0] andOp_236_out;
	andOp #(.WIDTH(1)) andOp_236(.in0(andOp_236_in0), .in1(andOp_236_in1), .out(andOp_236_out));

	reg [0:0] notOp_237_in0;
	wire [0:0] notOp_237_out;
	notOp #(.WIDTH(1)) notOp_237(.in(notOp_237_in0), .out(notOp_237_out));

	reg [0:0] andOp_238_in0;
	reg [0:0] andOp_238_in1;
	wire [0:0] andOp_238_out;
	andOp #(.WIDTH(1)) andOp_238(.in0(andOp_238_in0), .in1(andOp_238_in1), .out(andOp_238_out));

	reg [0:0] notOp_239_in0;
	wire [0:0] notOp_239_out;
	notOp #(.WIDTH(1)) notOp_239(.in(notOp_239_in0), .out(notOp_239_out));

	reg [0:0] andOp_240_in0;
	reg [0:0] andOp_240_in1;
	wire [0:0] andOp_240_out;
	andOp #(.WIDTH(1)) andOp_240(.in0(andOp_240_in0), .in1(andOp_240_in1), .out(andOp_240_out));

	reg [0:0] andOp_241_in0;
	reg [0:0] andOp_241_in1;
	wire [0:0] andOp_241_out;
	andOp #(.WIDTH(1)) andOp_241(.in0(andOp_241_in0), .in1(andOp_241_in1), .out(andOp_241_out));

	reg [31:0] eq_242_in0;
	reg [31:0] eq_242_in1;
	wire [0:0] eq_242_out;
	eq #(.WIDTH(32)) eq_242(.in0(eq_242_in0), .in1(eq_242_in1), .out(eq_242_out));

	reg [0:0] andOp_243_in0;
	reg [0:0] andOp_243_in1;
	wire [0:0] andOp_243_out;
	andOp #(.WIDTH(1)) andOp_243(.in0(andOp_243_in0), .in1(andOp_243_in1), .out(andOp_243_out));

	reg [0:0] notOp_244_in0;
	wire [0:0] notOp_244_out;
	notOp #(.WIDTH(1)) notOp_244(.in(notOp_244_in0), .out(notOp_244_out));

	reg [0:0] andOp_245_in0;
	reg [0:0] andOp_245_in1;
	wire [0:0] andOp_245_out;
	andOp #(.WIDTH(1)) andOp_245(.in0(andOp_245_in0), .in1(andOp_245_in1), .out(andOp_245_out));

	reg [0:0] notOp_246_in0;
	wire [0:0] notOp_246_out;
	notOp #(.WIDTH(1)) notOp_246(.in(notOp_246_in0), .out(notOp_246_out));

	reg [0:0] andOp_247_in0;
	reg [0:0] andOp_247_in1;
	wire [0:0] andOp_247_out;
	andOp #(.WIDTH(1)) andOp_247(.in0(andOp_247_in0), .in1(andOp_247_in1), .out(andOp_247_out));

	reg [0:0] notOp_248_in0;
	wire [0:0] notOp_248_out;
	notOp #(.WIDTH(1)) notOp_248(.in(notOp_248_in0), .out(notOp_248_out));

	reg [0:0] andOp_249_in0;
	reg [0:0] andOp_249_in1;
	wire [0:0] andOp_249_out;
	andOp #(.WIDTH(1)) andOp_249(.in0(andOp_249_in0), .in1(andOp_249_in1), .out(andOp_249_out));

	reg [0:0] andOp_250_in0;
	reg [0:0] andOp_250_in1;
	wire [0:0] andOp_250_out;
	andOp #(.WIDTH(1)) andOp_250(.in0(andOp_250_in0), .in1(andOp_250_in1), .out(andOp_250_out));

	reg [31:0] eq_251_in0;
	reg [31:0] eq_251_in1;
	wire [0:0] eq_251_out;
	eq #(.WIDTH(32)) eq_251(.in0(eq_251_in0), .in1(eq_251_in1), .out(eq_251_out));

	reg [0:0] andOp_252_in0;
	reg [0:0] andOp_252_in1;
	wire [0:0] andOp_252_out;
	andOp #(.WIDTH(1)) andOp_252(.in0(andOp_252_in0), .in1(andOp_252_in1), .out(andOp_252_out));

	reg [0:0] notOp_253_in0;
	wire [0:0] notOp_253_out;
	notOp #(.WIDTH(1)) notOp_253(.in(notOp_253_in0), .out(notOp_253_out));

	reg [0:0] andOp_254_in0;
	reg [0:0] andOp_254_in1;
	wire [0:0] andOp_254_out;
	andOp #(.WIDTH(1)) andOp_254(.in0(andOp_254_in0), .in1(andOp_254_in1), .out(andOp_254_out));

	reg [0:0] notOp_255_in0;
	wire [0:0] notOp_255_out;
	notOp #(.WIDTH(1)) notOp_255(.in(notOp_255_in0), .out(notOp_255_out));

	reg [0:0] andOp_256_in0;
	reg [0:0] andOp_256_in1;
	wire [0:0] andOp_256_out;
	andOp #(.WIDTH(1)) andOp_256(.in0(andOp_256_in0), .in1(andOp_256_in1), .out(andOp_256_out));

	reg [0:0] notOp_257_in0;
	wire [0:0] notOp_257_out;
	notOp #(.WIDTH(1)) notOp_257(.in(notOp_257_in0), .out(notOp_257_out));

	reg [0:0] andOp_258_in0;
	reg [0:0] andOp_258_in1;
	wire [0:0] andOp_258_out;
	andOp #(.WIDTH(1)) andOp_258(.in0(andOp_258_in0), .in1(andOp_258_in1), .out(andOp_258_out));

	reg [31:0] eq_259_in0;
	reg [31:0] eq_259_in1;
	wire [0:0] eq_259_out;
	eq #(.WIDTH(32)) eq_259(.in0(eq_259_in0), .in1(eq_259_in1), .out(eq_259_out));

	reg [31:0] eq_260_in0;
	reg [31:0] eq_260_in1;
	wire [0:0] eq_260_out;
	eq #(.WIDTH(32)) eq_260(.in0(eq_260_in0), .in1(eq_260_in1), .out(eq_260_out));

	reg [0:0] andOp_261_in0;
	reg [0:0] andOp_261_in1;
	wire [0:0] andOp_261_out;
	andOp #(.WIDTH(1)) andOp_261(.in0(andOp_261_in0), .in1(andOp_261_in1), .out(andOp_261_out));

	reg [31:0] eq_262_in0;
	reg [31:0] eq_262_in1;
	wire [0:0] eq_262_out;
	eq #(.WIDTH(32)) eq_262(.in0(eq_262_in0), .in1(eq_262_in1), .out(eq_262_out));

	reg [0:0] andOp_263_in0;
	reg [0:0] andOp_263_in1;
	wire [0:0] andOp_263_out;
	andOp #(.WIDTH(1)) andOp_263(.in0(andOp_263_in0), .in1(andOp_263_in1), .out(andOp_263_out));

	reg [0:0] notOp_264_in0;
	wire [0:0] notOp_264_out;
	notOp #(.WIDTH(1)) notOp_264(.in(notOp_264_in0), .out(notOp_264_out));

	reg [0:0] andOp_265_in0;
	reg [0:0] andOp_265_in1;
	wire [0:0] andOp_265_out;
	andOp #(.WIDTH(1)) andOp_265(.in0(andOp_265_in0), .in1(andOp_265_in1), .out(andOp_265_out));

	reg [0:0] notOp_266_in0;
	wire [0:0] notOp_266_out;
	notOp #(.WIDTH(1)) notOp_266(.in(notOp_266_in0), .out(notOp_266_out));

	reg [0:0] andOp_267_in0;
	reg [0:0] andOp_267_in1;
	wire [0:0] andOp_267_out;
	andOp #(.WIDTH(1)) andOp_267(.in0(andOp_267_in0), .in1(andOp_267_in1), .out(andOp_267_out));

	reg [0:0] notOp_268_in0;
	wire [0:0] notOp_268_out;
	notOp #(.WIDTH(1)) notOp_268(.in(notOp_268_in0), .out(notOp_268_out));

	reg [0:0] andOp_269_in0;
	reg [0:0] andOp_269_in1;
	wire [0:0] andOp_269_out;
	andOp #(.WIDTH(1)) andOp_269(.in0(andOp_269_in0), .in1(andOp_269_in1), .out(andOp_269_out));

	reg [0:0] andOp_270_in0;
	reg [0:0] andOp_270_in1;
	wire [0:0] andOp_270_out;
	andOp #(.WIDTH(1)) andOp_270(.in0(andOp_270_in0), .in1(andOp_270_in1), .out(andOp_270_out));

	reg [31:0] eq_271_in0;
	reg [31:0] eq_271_in1;
	wire [0:0] eq_271_out;
	eq #(.WIDTH(32)) eq_271(.in0(eq_271_in0), .in1(eq_271_in1), .out(eq_271_out));

	reg [0:0] andOp_272_in0;
	reg [0:0] andOp_272_in1;
	wire [0:0] andOp_272_out;
	andOp #(.WIDTH(1)) andOp_272(.in0(andOp_272_in0), .in1(andOp_272_in1), .out(andOp_272_out));

	reg [0:0] notOp_273_in0;
	wire [0:0] notOp_273_out;
	notOp #(.WIDTH(1)) notOp_273(.in(notOp_273_in0), .out(notOp_273_out));

	reg [0:0] andOp_274_in0;
	reg [0:0] andOp_274_in1;
	wire [0:0] andOp_274_out;
	andOp #(.WIDTH(1)) andOp_274(.in0(andOp_274_in0), .in1(andOp_274_in1), .out(andOp_274_out));

	reg [0:0] notOp_275_in0;
	wire [0:0] notOp_275_out;
	notOp #(.WIDTH(1)) notOp_275(.in(notOp_275_in0), .out(notOp_275_out));

	reg [0:0] andOp_276_in0;
	reg [0:0] andOp_276_in1;
	wire [0:0] andOp_276_out;
	andOp #(.WIDTH(1)) andOp_276(.in0(andOp_276_in0), .in1(andOp_276_in1), .out(andOp_276_out));

	reg [0:0] notOp_277_in0;
	wire [0:0] notOp_277_out;
	notOp #(.WIDTH(1)) notOp_277(.in(notOp_277_in0), .out(notOp_277_out));

	reg [0:0] andOp_278_in0;
	reg [0:0] andOp_278_in1;
	wire [0:0] andOp_278_out;
	andOp #(.WIDTH(1)) andOp_278(.in0(andOp_278_in0), .in1(andOp_278_in1), .out(andOp_278_out));

	reg [0:0] andOp_279_in0;
	reg [0:0] andOp_279_in1;
	wire [0:0] andOp_279_out;
	andOp #(.WIDTH(1)) andOp_279(.in0(andOp_279_in0), .in1(andOp_279_in1), .out(andOp_279_out));

	reg [31:0] eq_280_in0;
	reg [31:0] eq_280_in1;
	wire [0:0] eq_280_out;
	eq #(.WIDTH(32)) eq_280(.in0(eq_280_in0), .in1(eq_280_in1), .out(eq_280_out));

	reg [0:0] andOp_281_in0;
	reg [0:0] andOp_281_in1;
	wire [0:0] andOp_281_out;
	andOp #(.WIDTH(1)) andOp_281(.in0(andOp_281_in0), .in1(andOp_281_in1), .out(andOp_281_out));

	reg [0:0] notOp_282_in0;
	wire [0:0] notOp_282_out;
	notOp #(.WIDTH(1)) notOp_282(.in(notOp_282_in0), .out(notOp_282_out));

	reg [0:0] andOp_283_in0;
	reg [0:0] andOp_283_in1;
	wire [0:0] andOp_283_out;
	andOp #(.WIDTH(1)) andOp_283(.in0(andOp_283_in0), .in1(andOp_283_in1), .out(andOp_283_out));

	reg [0:0] notOp_284_in0;
	wire [0:0] notOp_284_out;
	notOp #(.WIDTH(1)) notOp_284(.in(notOp_284_in0), .out(notOp_284_out));

	reg [0:0] andOp_285_in0;
	reg [0:0] andOp_285_in1;
	wire [0:0] andOp_285_out;
	andOp #(.WIDTH(1)) andOp_285(.in0(andOp_285_in0), .in1(andOp_285_in1), .out(andOp_285_out));

	reg [0:0] notOp_286_in0;
	wire [0:0] notOp_286_out;
	notOp #(.WIDTH(1)) notOp_286(.in(notOp_286_in0), .out(notOp_286_out));

	reg [0:0] andOp_287_in0;
	reg [0:0] andOp_287_in1;
	wire [0:0] andOp_287_out;
	andOp #(.WIDTH(1)) andOp_287(.in0(andOp_287_in0), .in1(andOp_287_in1), .out(andOp_287_out));

	reg [0:0] andOp_288_in0;
	reg [0:0] andOp_288_in1;
	wire [0:0] andOp_288_out;
	andOp #(.WIDTH(1)) andOp_288(.in0(andOp_288_in0), .in1(andOp_288_in1), .out(andOp_288_out));

	reg [31:0] eq_289_in0;
	reg [31:0] eq_289_in1;
	wire [0:0] eq_289_out;
	eq #(.WIDTH(32)) eq_289(.in0(eq_289_in0), .in1(eq_289_in1), .out(eq_289_out));

	reg [0:0] andOp_290_in0;
	reg [0:0] andOp_290_in1;
	wire [0:0] andOp_290_out;
	andOp #(.WIDTH(1)) andOp_290(.in0(andOp_290_in0), .in1(andOp_290_in1), .out(andOp_290_out));

	reg [0:0] notOp_291_in0;
	wire [0:0] notOp_291_out;
	notOp #(.WIDTH(1)) notOp_291(.in(notOp_291_in0), .out(notOp_291_out));

	reg [0:0] andOp_292_in0;
	reg [0:0] andOp_292_in1;
	wire [0:0] andOp_292_out;
	andOp #(.WIDTH(1)) andOp_292(.in0(andOp_292_in0), .in1(andOp_292_in1), .out(andOp_292_out));

	reg [0:0] notOp_293_in0;
	wire [0:0] notOp_293_out;
	notOp #(.WIDTH(1)) notOp_293(.in(notOp_293_in0), .out(notOp_293_out));

	reg [0:0] andOp_294_in0;
	reg [0:0] andOp_294_in1;
	wire [0:0] andOp_294_out;
	andOp #(.WIDTH(1)) andOp_294(.in0(andOp_294_in0), .in1(andOp_294_in1), .out(andOp_294_out));

	reg [0:0] notOp_295_in0;
	wire [0:0] notOp_295_out;
	notOp #(.WIDTH(1)) notOp_295(.in(notOp_295_in0), .out(notOp_295_out));

	reg [0:0] andOp_296_in0;
	reg [0:0] andOp_296_in1;
	wire [0:0] andOp_296_out;
	andOp #(.WIDTH(1)) andOp_296(.in0(andOp_296_in0), .in1(andOp_296_in1), .out(andOp_296_out));

	reg [31:0] eq_297_in0;
	reg [31:0] eq_297_in1;
	wire [0:0] eq_297_out;
	eq #(.WIDTH(32)) eq_297(.in0(eq_297_in0), .in1(eq_297_in1), .out(eq_297_out));

	reg [31:0] eq_298_in0;
	reg [31:0] eq_298_in1;
	wire [0:0] eq_298_out;
	eq #(.WIDTH(32)) eq_298(.in0(eq_298_in0), .in1(eq_298_in1), .out(eq_298_out));

	reg [0:0] andOp_299_in0;
	reg [0:0] andOp_299_in1;
	wire [0:0] andOp_299_out;
	andOp #(.WIDTH(1)) andOp_299(.in0(andOp_299_in0), .in1(andOp_299_in1), .out(andOp_299_out));

	reg [31:0] eq_300_in0;
	reg [31:0] eq_300_in1;
	wire [0:0] eq_300_out;
	eq #(.WIDTH(32)) eq_300(.in0(eq_300_in0), .in1(eq_300_in1), .out(eq_300_out));

	reg [0:0] andOp_301_in0;
	reg [0:0] andOp_301_in1;
	wire [0:0] andOp_301_out;
	andOp #(.WIDTH(1)) andOp_301(.in0(andOp_301_in0), .in1(andOp_301_in1), .out(andOp_301_out));

	reg [0:0] notOp_302_in0;
	wire [0:0] notOp_302_out;
	notOp #(.WIDTH(1)) notOp_302(.in(notOp_302_in0), .out(notOp_302_out));

	reg [0:0] andOp_303_in0;
	reg [0:0] andOp_303_in1;
	wire [0:0] andOp_303_out;
	andOp #(.WIDTH(1)) andOp_303(.in0(andOp_303_in0), .in1(andOp_303_in1), .out(andOp_303_out));

	reg [0:0] notOp_304_in0;
	wire [0:0] notOp_304_out;
	notOp #(.WIDTH(1)) notOp_304(.in(notOp_304_in0), .out(notOp_304_out));

	reg [0:0] andOp_305_in0;
	reg [0:0] andOp_305_in1;
	wire [0:0] andOp_305_out;
	andOp #(.WIDTH(1)) andOp_305(.in0(andOp_305_in0), .in1(andOp_305_in1), .out(andOp_305_out));

	reg [0:0] notOp_306_in0;
	wire [0:0] notOp_306_out;
	notOp #(.WIDTH(1)) notOp_306(.in(notOp_306_in0), .out(notOp_306_out));

	reg [0:0] andOp_307_in0;
	reg [0:0] andOp_307_in1;
	wire [0:0] andOp_307_out;
	andOp #(.WIDTH(1)) andOp_307(.in0(andOp_307_in0), .in1(andOp_307_in1), .out(andOp_307_out));

	reg [0:0] andOp_308_in0;
	reg [0:0] andOp_308_in1;
	wire [0:0] andOp_308_out;
	andOp #(.WIDTH(1)) andOp_308(.in0(andOp_308_in0), .in1(andOp_308_in1), .out(andOp_308_out));

	reg [31:0] eq_309_in0;
	reg [31:0] eq_309_in1;
	wire [0:0] eq_309_out;
	eq #(.WIDTH(32)) eq_309(.in0(eq_309_in0), .in1(eq_309_in1), .out(eq_309_out));

	reg [0:0] andOp_310_in0;
	reg [0:0] andOp_310_in1;
	wire [0:0] andOp_310_out;
	andOp #(.WIDTH(1)) andOp_310(.in0(andOp_310_in0), .in1(andOp_310_in1), .out(andOp_310_out));

	reg [0:0] notOp_311_in0;
	wire [0:0] notOp_311_out;
	notOp #(.WIDTH(1)) notOp_311(.in(notOp_311_in0), .out(notOp_311_out));

	reg [0:0] andOp_312_in0;
	reg [0:0] andOp_312_in1;
	wire [0:0] andOp_312_out;
	andOp #(.WIDTH(1)) andOp_312(.in0(andOp_312_in0), .in1(andOp_312_in1), .out(andOp_312_out));

	reg [0:0] notOp_313_in0;
	wire [0:0] notOp_313_out;
	notOp #(.WIDTH(1)) notOp_313(.in(notOp_313_in0), .out(notOp_313_out));

	reg [0:0] andOp_314_in0;
	reg [0:0] andOp_314_in1;
	wire [0:0] andOp_314_out;
	andOp #(.WIDTH(1)) andOp_314(.in0(andOp_314_in0), .in1(andOp_314_in1), .out(andOp_314_out));

	reg [0:0] notOp_315_in0;
	wire [0:0] notOp_315_out;
	notOp #(.WIDTH(1)) notOp_315(.in(notOp_315_in0), .out(notOp_315_out));

	reg [0:0] andOp_316_in0;
	reg [0:0] andOp_316_in1;
	wire [0:0] andOp_316_out;
	andOp #(.WIDTH(1)) andOp_316(.in0(andOp_316_in0), .in1(andOp_316_in1), .out(andOp_316_out));

	reg [0:0] andOp_317_in0;
	reg [0:0] andOp_317_in1;
	wire [0:0] andOp_317_out;
	andOp #(.WIDTH(1)) andOp_317(.in0(andOp_317_in0), .in1(andOp_317_in1), .out(andOp_317_out));

	reg [31:0] eq_318_in0;
	reg [31:0] eq_318_in1;
	wire [0:0] eq_318_out;
	eq #(.WIDTH(32)) eq_318(.in0(eq_318_in0), .in1(eq_318_in1), .out(eq_318_out));

	reg [0:0] andOp_319_in0;
	reg [0:0] andOp_319_in1;
	wire [0:0] andOp_319_out;
	andOp #(.WIDTH(1)) andOp_319(.in0(andOp_319_in0), .in1(andOp_319_in1), .out(andOp_319_out));

	reg [0:0] notOp_320_in0;
	wire [0:0] notOp_320_out;
	notOp #(.WIDTH(1)) notOp_320(.in(notOp_320_in0), .out(notOp_320_out));

	reg [0:0] andOp_321_in0;
	reg [0:0] andOp_321_in1;
	wire [0:0] andOp_321_out;
	andOp #(.WIDTH(1)) andOp_321(.in0(andOp_321_in0), .in1(andOp_321_in1), .out(andOp_321_out));

	reg [0:0] notOp_322_in0;
	wire [0:0] notOp_322_out;
	notOp #(.WIDTH(1)) notOp_322(.in(notOp_322_in0), .out(notOp_322_out));

	reg [0:0] andOp_323_in0;
	reg [0:0] andOp_323_in1;
	wire [0:0] andOp_323_out;
	andOp #(.WIDTH(1)) andOp_323(.in0(andOp_323_in0), .in1(andOp_323_in1), .out(andOp_323_out));

	reg [0:0] notOp_324_in0;
	wire [0:0] notOp_324_out;
	notOp #(.WIDTH(1)) notOp_324(.in(notOp_324_in0), .out(notOp_324_out));

	reg [0:0] andOp_325_in0;
	reg [0:0] andOp_325_in1;
	wire [0:0] andOp_325_out;
	andOp #(.WIDTH(1)) andOp_325(.in0(andOp_325_in0), .in1(andOp_325_in1), .out(andOp_325_out));

	reg [0:0] andOp_326_in0;
	reg [0:0] andOp_326_in1;
	wire [0:0] andOp_326_out;
	andOp #(.WIDTH(1)) andOp_326(.in0(andOp_326_in0), .in1(andOp_326_in1), .out(andOp_326_out));

	reg [31:0] eq_327_in0;
	reg [31:0] eq_327_in1;
	wire [0:0] eq_327_out;
	eq #(.WIDTH(32)) eq_327(.in0(eq_327_in0), .in1(eq_327_in1), .out(eq_327_out));

	reg [0:0] andOp_328_in0;
	reg [0:0] andOp_328_in1;
	wire [0:0] andOp_328_out;
	andOp #(.WIDTH(1)) andOp_328(.in0(andOp_328_in0), .in1(andOp_328_in1), .out(andOp_328_out));

	reg [0:0] notOp_329_in0;
	wire [0:0] notOp_329_out;
	notOp #(.WIDTH(1)) notOp_329(.in(notOp_329_in0), .out(notOp_329_out));

	reg [0:0] andOp_330_in0;
	reg [0:0] andOp_330_in1;
	wire [0:0] andOp_330_out;
	andOp #(.WIDTH(1)) andOp_330(.in0(andOp_330_in0), .in1(andOp_330_in1), .out(andOp_330_out));

	reg [0:0] notOp_331_in0;
	wire [0:0] notOp_331_out;
	notOp #(.WIDTH(1)) notOp_331(.in(notOp_331_in0), .out(notOp_331_out));

	reg [0:0] andOp_332_in0;
	reg [0:0] andOp_332_in1;
	wire [0:0] andOp_332_out;
	andOp #(.WIDTH(1)) andOp_332(.in0(andOp_332_in0), .in1(andOp_332_in1), .out(andOp_332_out));

	reg [0:0] notOp_333_in0;
	wire [0:0] notOp_333_out;
	notOp #(.WIDTH(1)) notOp_333(.in(notOp_333_in0), .out(notOp_333_out));

	reg [0:0] andOp_334_in0;
	reg [0:0] andOp_334_in1;
	wire [0:0] andOp_334_out;
	andOp #(.WIDTH(1)) andOp_334(.in0(andOp_334_in0), .in1(andOp_334_in1), .out(andOp_334_out));

	// End Functional Units

	reg [31:0] data_store_1_0;
	reg [31:0] data_store_1_2;
	reg [0:0] data_store_1_4;
	reg [31:0] data_store_1_6;
	reg [31:0] data_store_2_10;
	reg [0:0] data_store_2_12;
	reg [31:0] data_store_2_14;
	reg [31:0] data_store_2_8;
	reg [31:0] data_store_3_16;
	reg [31:0] data_store_3_18;
	reg [0:0] data_store_3_20;
	reg [31:0] data_store_3_22;
	reg [31:0] data_store_4_24;
	reg [31:0] data_store_4_26;
	reg [0:0] data_store_4_28;
	reg [31:0] data_store_4_30;
	reg [31:0] global_state;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_3_last_state;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;
	reg [31:0] state_4_last_state;

	// controller for add_add_12.add_in0_add_12
	// controller for add_add_12.add_in1_add_12
	// Insensitive connections
	always @(*) begin
		add_in0_add_12 = valid ? rdata_ram_0 : rdata_ram_0;
		add_in1_add_12 = valid ? tmp_output_152_out_data : tmp_output_152_out_data;
	end
	// controller for add_add_14.add_in0_add_14
	// controller for add_add_14.add_in1_add_14
	// Insensitive connections
	always @(*) begin
		add_in0_add_14 = valid ? data_in_3_17_out_data : data_in_3_17_out_data;
		add_in1_add_14 = valid ? 32'd1 : 32'd1;
	end
	// controller for andOp_110.andOp_110_in0
	// controller for andOp_110.andOp_110_in1
	// Insensitive connections
	always @(*) begin
		andOp_110_in0 = valid ? notOp_109_out : notOp_109_out;
		andOp_110_in1 = valid ? andOp_33_out : andOp_33_out;
	end
	// controller for andOp_113.andOp_113_in0
	// controller for andOp_113.andOp_113_in1
	// Insensitive connections
	always @(*) begin
		andOp_113_in0 = valid ? notOp_112_out : notOp_112_out;
		andOp_113_in1 = valid ? andOp_48_out : andOp_48_out;
	end
	// controller for andOp_116.andOp_116_in0
	// controller for andOp_116.andOp_116_in1
	// Insensitive connections
	always @(*) begin
		andOp_116_in0 = valid ? notOp_115_out : notOp_115_out;
		andOp_116_in1 = valid ? andOp_39_out : andOp_39_out;
	end
	// controller for andOp_121.andOp_121_in0
	// controller for andOp_121.andOp_121_in1
	// Insensitive connections
	always @(*) begin
		andOp_121_in0 = valid ? notOp_120_out : notOp_120_out;
		andOp_121_in1 = valid ? andOp_51_out : andOp_51_out;
	end
	// controller for andOp_124.andOp_124_in0
	// controller for andOp_124.andOp_124_in1
	// Insensitive connections
	always @(*) begin
		andOp_124_in0 = valid ? notOp_123_out : notOp_123_out;
		andOp_124_in1 = valid ? andOp_59_out : andOp_59_out;
	end
	// controller for andOp_127.andOp_127_in0
	// controller for andOp_127.andOp_127_in1
	// Insensitive connections
	always @(*) begin
		andOp_127_in0 = valid ? notOp_126_out : notOp_126_out;
		andOp_127_in1 = valid ? andOp_75_out : andOp_75_out;
	end
	// controller for andOp_130.andOp_130_in0
	// controller for andOp_130.andOp_130_in1
	// Insensitive connections
	always @(*) begin
		andOp_130_in0 = valid ? notOp_129_out : notOp_129_out;
		andOp_130_in1 = valid ? andOp_63_out : andOp_63_out;
	end
	// controller for andOp_133.andOp_133_in0
	// controller for andOp_133.andOp_133_in1
	// Insensitive connections
	always @(*) begin
		andOp_133_in0 = valid ? notOp_132_out : notOp_132_out;
		andOp_133_in1 = valid ? andOp_66_out : andOp_66_out;
	end
	// controller for andOp_136.andOp_136_in0
	// controller for andOp_136.andOp_136_in1
	// Insensitive connections
	always @(*) begin
		andOp_136_in0 = valid ? notOp_135_out : notOp_135_out;
		andOp_136_in1 = valid ? andOp_71_out : andOp_71_out;
	end
	// controller for andOp_138.andOp_138_in0
	// controller for andOp_138.andOp_138_in1
	// Insensitive connections
	always @(*) begin
		andOp_138_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_138_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_139.andOp_139_in0
	// controller for andOp_139.andOp_139_in1
	// Insensitive connections
	always @(*) begin
		andOp_139_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_139_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_140.andOp_140_in0
	// controller for andOp_140.andOp_140_in1
	// Insensitive connections
	always @(*) begin
		andOp_140_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_140_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_141.andOp_141_in0
	// controller for andOp_141.andOp_141_in1
	// Insensitive connections
	always @(*) begin
		andOp_141_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_141_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_142.andOp_142_in0
	// controller for andOp_142.andOp_142_in1
	// Insensitive connections
	always @(*) begin
		andOp_142_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_142_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_143.andOp_143_in0
	// controller for andOp_143.andOp_143_in1
	// Insensitive connections
	always @(*) begin
		andOp_143_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_143_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_144.andOp_144_in0
	// controller for andOp_144.andOp_144_in1
	// Insensitive connections
	always @(*) begin
		andOp_144_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_144_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_145.andOp_145_in0
	// controller for andOp_145.andOp_145_in1
	// Insensitive connections
	always @(*) begin
		andOp_145_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_145_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_148.andOp_148_in0
	// controller for andOp_148.andOp_148_in1
	// Insensitive connections
	always @(*) begin
		andOp_148_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
		andOp_148_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_149.andOp_149_in0
	// controller for andOp_149.andOp_149_in1
	// Insensitive connections
	always @(*) begin
		andOp_149_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_149_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_150.andOp_150_in0
	// controller for andOp_150.andOp_150_in1
	// Insensitive connections
	always @(*) begin
		andOp_150_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_150_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_151.andOp_151_in0
	// controller for andOp_151.andOp_151_in1
	// Insensitive connections
	always @(*) begin
		andOp_151_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_151_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_154.andOp_154_in0
	// controller for andOp_154.andOp_154_in1
	// Insensitive connections
	always @(*) begin
		andOp_154_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_154_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_155.andOp_155_in0
	// controller for andOp_155.andOp_155_in1
	// Insensitive connections
	always @(*) begin
		andOp_155_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_155_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_156.andOp_156_in0
	// controller for andOp_156.andOp_156_in1
	// Insensitive connections
	always @(*) begin
		andOp_156_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_156_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_157.andOp_157_in0
	// controller for andOp_157.andOp_157_in1
	// Insensitive connections
	always @(*) begin
		andOp_157_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_157_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_158.andOp_158_in0
	// controller for andOp_158.andOp_158_in1
	// Insensitive connections
	always @(*) begin
		andOp_158_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_158_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_159.andOp_159_in0
	// controller for andOp_159.andOp_159_in1
	// Insensitive connections
	always @(*) begin
		andOp_159_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_159_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_160.andOp_160_in0
	// controller for andOp_160.andOp_160_in1
	// Insensitive connections
	always @(*) begin
		andOp_160_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
		andOp_160_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_161.andOp_161_in0
	// controller for andOp_161.andOp_161_in1
	// Insensitive connections
	always @(*) begin
		andOp_161_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_161_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_162.andOp_162_in0
	// controller for andOp_162.andOp_162_in1
	// Insensitive connections
	always @(*) begin
		andOp_162_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_162_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_163.andOp_163_in0
	// controller for andOp_163.andOp_163_in1
	// Insensitive connections
	always @(*) begin
		andOp_163_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_163_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_164.andOp_164_in0
	// controller for andOp_164.andOp_164_in1
	// Insensitive connections
	always @(*) begin
		andOp_164_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_164_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_166.andOp_166_in0
	// controller for andOp_166.andOp_166_in1
	// Insensitive connections
	always @(*) begin
		andOp_166_in0 = valid ? notOp_165_out : notOp_165_out;
		andOp_166_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_168.andOp_168_in0
	// controller for andOp_168.andOp_168_in1
	// Insensitive connections
	always @(*) begin
		andOp_168_in0 = valid ? notOp_167_out : notOp_167_out;
		andOp_168_in1 = valid ? andOp_166_out : andOp_166_out;
	end
	// controller for andOp_170.andOp_170_in0
	// controller for andOp_170.andOp_170_in1
	// Insensitive connections
	always @(*) begin
		andOp_170_in0 = valid ? notOp_169_out : notOp_169_out;
		andOp_170_in1 = valid ? andOp_168_out : andOp_168_out;
	end
	// controller for andOp_172.andOp_172_in0
	// controller for andOp_172.andOp_172_in1
	// Insensitive connections
	always @(*) begin
		andOp_172_in0 = valid ? notOp_171_out : notOp_171_out;
		andOp_172_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_174.andOp_174_in0
	// controller for andOp_174.andOp_174_in1
	// Insensitive connections
	always @(*) begin
		andOp_174_in0 = valid ? notOp_173_out : notOp_173_out;
		andOp_174_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_176.andOp_176_in0
	// controller for andOp_176.andOp_176_in1
	// Insensitive connections
	always @(*) begin
		andOp_176_in0 = valid ? notOp_175_out : notOp_175_out;
		andOp_176_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_178.andOp_178_in0
	// controller for andOp_178.andOp_178_in1
	// Insensitive connections
	always @(*) begin
		andOp_178_in0 = valid ? notOp_177_out : notOp_177_out;
		andOp_178_in1 = valid ? andOp_176_out : andOp_176_out;
	end
	// controller for andOp_180.andOp_180_in0
	// controller for andOp_180.andOp_180_in1
	// Insensitive connections
	always @(*) begin
		andOp_180_in0 = valid ? notOp_179_out : notOp_179_out;
		andOp_180_in1 = valid ? andOp_178_out : andOp_178_out;
	end
	// controller for andOp_185.andOp_185_in0
	// controller for andOp_185.andOp_185_in1
	// Insensitive connections
	always @(*) begin
		andOp_185_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_185_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_187.andOp_187_in0
	// controller for andOp_187.andOp_187_in1
	// Insensitive connections
	always @(*) begin
		andOp_187_in0 = valid ? andOp_185_out : andOp_185_out;
		andOp_187_in1 = valid ? eq_186_out : eq_186_out;
	end
	// controller for andOp_189.andOp_189_in0
	// controller for andOp_189.andOp_189_in1
	// Insensitive connections
	always @(*) begin
		andOp_189_in0 = valid ? andOp_185_out : andOp_185_out;
		andOp_189_in1 = valid ? notOp_188_out : notOp_188_out;
	end
	// controller for andOp_191.andOp_191_in0
	// controller for andOp_191.andOp_191_in1
	// Insensitive connections
	always @(*) begin
		andOp_191_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_191_in1 = valid ? notOp_190_out : notOp_190_out;
	end
	// controller for andOp_193.andOp_193_in0
	// controller for andOp_193.andOp_193_in1
	// Insensitive connections
	always @(*) begin
		andOp_193_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_193_in1 = valid ? notOp_192_out : notOp_192_out;
	end
	// controller for andOp_194.andOp_194_in0
	// controller for andOp_194.andOp_194_in1
	// Insensitive connections
	always @(*) begin
		andOp_194_in0 = valid ? 1'd0 : 1'd0;
		andOp_194_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_196.andOp_196_in0
	// controller for andOp_196.andOp_196_in1
	// Insensitive connections
	always @(*) begin
		andOp_196_in0 = valid ? andOp_194_out : andOp_194_out;
		andOp_196_in1 = valid ? eq_195_out : eq_195_out;
	end
	// controller for andOp_198.andOp_198_in0
	// controller for andOp_198.andOp_198_in1
	// Insensitive connections
	always @(*) begin
		andOp_198_in0 = valid ? andOp_194_out : andOp_194_out;
		andOp_198_in1 = valid ? notOp_197_out : notOp_197_out;
	end
	// controller for andOp_200.andOp_200_in0
	// controller for andOp_200.andOp_200_in1
	// Insensitive connections
	always @(*) begin
		andOp_200_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_200_in1 = valid ? notOp_199_out : notOp_199_out;
	end
	// controller for andOp_202.andOp_202_in0
	// controller for andOp_202.andOp_202_in1
	// Insensitive connections
	always @(*) begin
		andOp_202_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_202_in1 = valid ? notOp_201_out : notOp_201_out;
	end
	// controller for andOp_203.andOp_203_in0
	// controller for andOp_203.andOp_203_in1
	// Insensitive connections
	always @(*) begin
		andOp_203_in0 = valid ? 1'd0 : 1'd0;
		andOp_203_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_205.andOp_205_in0
	// controller for andOp_205.andOp_205_in1
	// Insensitive connections
	always @(*) begin
		andOp_205_in0 = valid ? andOp_203_out : andOp_203_out;
		andOp_205_in1 = valid ? eq_204_out : eq_204_out;
	end
	// controller for andOp_207.andOp_207_in0
	// controller for andOp_207.andOp_207_in1
	// Insensitive connections
	always @(*) begin
		andOp_207_in0 = valid ? andOp_203_out : andOp_203_out;
		andOp_207_in1 = valid ? notOp_206_out : notOp_206_out;
	end
	// controller for andOp_209.andOp_209_in0
	// controller for andOp_209.andOp_209_in1
	// Insensitive connections
	always @(*) begin
		andOp_209_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_209_in1 = valid ? notOp_208_out : notOp_208_out;
	end
	// controller for andOp_211.andOp_211_in0
	// controller for andOp_211.andOp_211_in1
	// Insensitive connections
	always @(*) begin
		andOp_211_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_211_in1 = valid ? notOp_210_out : notOp_210_out;
	end
	// controller for andOp_212.andOp_212_in0
	// controller for andOp_212.andOp_212_in1
	// Insensitive connections
	always @(*) begin
		andOp_212_in0 = valid ? 1'd0 : 1'd0;
		andOp_212_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_214.andOp_214_in0
	// controller for andOp_214.andOp_214_in1
	// Insensitive connections
	always @(*) begin
		andOp_214_in0 = valid ? andOp_212_out : andOp_212_out;
		andOp_214_in1 = valid ? eq_213_out : eq_213_out;
	end
	// controller for andOp_216.andOp_216_in0
	// controller for andOp_216.andOp_216_in1
	// Insensitive connections
	always @(*) begin
		andOp_216_in0 = valid ? andOp_212_out : andOp_212_out;
		andOp_216_in1 = valid ? notOp_215_out : notOp_215_out;
	end
	// controller for andOp_218.andOp_218_in0
	// controller for andOp_218.andOp_218_in1
	// Insensitive connections
	always @(*) begin
		andOp_218_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_218_in1 = valid ? notOp_217_out : notOp_217_out;
	end
	// controller for andOp_220.andOp_220_in0
	// controller for andOp_220.andOp_220_in1
	// Insensitive connections
	always @(*) begin
		andOp_220_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_220_in1 = valid ? notOp_219_out : notOp_219_out;
	end
	// controller for andOp_223.andOp_223_in0
	// controller for andOp_223.andOp_223_in1
	// Insensitive connections
	always @(*) begin
		andOp_223_in0 = valid ? 1'd0 : 1'd0;
		andOp_223_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_225.andOp_225_in0
	// controller for andOp_225.andOp_225_in1
	// Insensitive connections
	always @(*) begin
		andOp_225_in0 = valid ? andOp_223_out : andOp_223_out;
		andOp_225_in1 = valid ? eq_224_out : eq_224_out;
	end
	// controller for andOp_227.andOp_227_in0
	// controller for andOp_227.andOp_227_in1
	// Insensitive connections
	always @(*) begin
		andOp_227_in0 = valid ? andOp_223_out : andOp_223_out;
		andOp_227_in1 = valid ? notOp_226_out : notOp_226_out;
	end
	// controller for andOp_229.andOp_229_in0
	// controller for andOp_229.andOp_229_in1
	// Insensitive connections
	always @(*) begin
		andOp_229_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_229_in1 = valid ? notOp_228_out : notOp_228_out;
	end
	// controller for andOp_231.andOp_231_in0
	// controller for andOp_231.andOp_231_in1
	// Insensitive connections
	always @(*) begin
		andOp_231_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_231_in1 = valid ? notOp_230_out : notOp_230_out;
	end
	// controller for andOp_232.andOp_232_in0
	// controller for andOp_232.andOp_232_in1
	// Insensitive connections
	always @(*) begin
		andOp_232_in0 = valid ? 1'd0 : 1'd0;
		andOp_232_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_234.andOp_234_in0
	// controller for andOp_234.andOp_234_in1
	// Insensitive connections
	always @(*) begin
		andOp_234_in0 = valid ? andOp_232_out : andOp_232_out;
		andOp_234_in1 = valid ? eq_233_out : eq_233_out;
	end
	// controller for andOp_236.andOp_236_in0
	// controller for andOp_236.andOp_236_in1
	// Insensitive connections
	always @(*) begin
		andOp_236_in0 = valid ? andOp_232_out : andOp_232_out;
		andOp_236_in1 = valid ? notOp_235_out : notOp_235_out;
	end
	// controller for andOp_238.andOp_238_in0
	// controller for andOp_238.andOp_238_in1
	// Insensitive connections
	always @(*) begin
		andOp_238_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_238_in1 = valid ? notOp_237_out : notOp_237_out;
	end
	// controller for andOp_240.andOp_240_in0
	// controller for andOp_240.andOp_240_in1
	// Insensitive connections
	always @(*) begin
		andOp_240_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_240_in1 = valid ? notOp_239_out : notOp_239_out;
	end
	// controller for andOp_241.andOp_241_in0
	// controller for andOp_241.andOp_241_in1
	// Insensitive connections
	always @(*) begin
		andOp_241_in0 = valid ? 1'd0 : 1'd0;
		andOp_241_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_243.andOp_243_in0
	// controller for andOp_243.andOp_243_in1
	// Insensitive connections
	always @(*) begin
		andOp_243_in0 = valid ? andOp_241_out : andOp_241_out;
		andOp_243_in1 = valid ? eq_242_out : eq_242_out;
	end
	// controller for andOp_245.andOp_245_in0
	// controller for andOp_245.andOp_245_in1
	// Insensitive connections
	always @(*) begin
		andOp_245_in0 = valid ? andOp_241_out : andOp_241_out;
		andOp_245_in1 = valid ? notOp_244_out : notOp_244_out;
	end
	// controller for andOp_247.andOp_247_in0
	// controller for andOp_247.andOp_247_in1
	// Insensitive connections
	always @(*) begin
		andOp_247_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_247_in1 = valid ? notOp_246_out : notOp_246_out;
	end
	// controller for andOp_249.andOp_249_in0
	// controller for andOp_249.andOp_249_in1
	// Insensitive connections
	always @(*) begin
		andOp_249_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_249_in1 = valid ? notOp_248_out : notOp_248_out;
	end
	// controller for andOp_250.andOp_250_in0
	// controller for andOp_250.andOp_250_in1
	// Insensitive connections
	always @(*) begin
		andOp_250_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_250_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_252.andOp_252_in0
	// controller for andOp_252.andOp_252_in1
	// Insensitive connections
	always @(*) begin
		andOp_252_in0 = valid ? andOp_250_out : andOp_250_out;
		andOp_252_in1 = valid ? eq_251_out : eq_251_out;
	end
	// controller for andOp_254.andOp_254_in0
	// controller for andOp_254.andOp_254_in1
	// Insensitive connections
	always @(*) begin
		andOp_254_in0 = valid ? andOp_250_out : andOp_250_out;
		andOp_254_in1 = valid ? notOp_253_out : notOp_253_out;
	end
	// controller for andOp_256.andOp_256_in0
	// controller for andOp_256.andOp_256_in1
	// Insensitive connections
	always @(*) begin
		andOp_256_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_256_in1 = valid ? notOp_255_out : notOp_255_out;
	end
	// controller for andOp_258.andOp_258_in0
	// controller for andOp_258.andOp_258_in1
	// Insensitive connections
	always @(*) begin
		andOp_258_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_258_in1 = valid ? notOp_257_out : notOp_257_out;
	end
	// controller for andOp_261.andOp_261_in0
	// controller for andOp_261.andOp_261_in1
	// Insensitive connections
	always @(*) begin
		andOp_261_in0 = valid ? 1'd0 : 1'd0;
		andOp_261_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_263.andOp_263_in0
	// controller for andOp_263.andOp_263_in1
	// Insensitive connections
	always @(*) begin
		andOp_263_in0 = valid ? andOp_261_out : andOp_261_out;
		andOp_263_in1 = valid ? eq_262_out : eq_262_out;
	end
	// controller for andOp_265.andOp_265_in0
	// controller for andOp_265.andOp_265_in1
	// Insensitive connections
	always @(*) begin
		andOp_265_in0 = valid ? andOp_261_out : andOp_261_out;
		andOp_265_in1 = valid ? notOp_264_out : notOp_264_out;
	end
	// controller for andOp_267.andOp_267_in0
	// controller for andOp_267.andOp_267_in1
	// Insensitive connections
	always @(*) begin
		andOp_267_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_267_in1 = valid ? notOp_266_out : notOp_266_out;
	end
	// controller for andOp_269.andOp_269_in0
	// controller for andOp_269.andOp_269_in1
	// Insensitive connections
	always @(*) begin
		andOp_269_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_269_in1 = valid ? notOp_268_out : notOp_268_out;
	end
	// controller for andOp_270.andOp_270_in0
	// controller for andOp_270.andOp_270_in1
	// Insensitive connections
	always @(*) begin
		andOp_270_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_270_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_272.andOp_272_in0
	// controller for andOp_272.andOp_272_in1
	// Insensitive connections
	always @(*) begin
		andOp_272_in0 = valid ? andOp_270_out : andOp_270_out;
		andOp_272_in1 = valid ? eq_271_out : eq_271_out;
	end
	// controller for andOp_274.andOp_274_in0
	// controller for andOp_274.andOp_274_in1
	// Insensitive connections
	always @(*) begin
		andOp_274_in0 = valid ? andOp_270_out : andOp_270_out;
		andOp_274_in1 = valid ? notOp_273_out : notOp_273_out;
	end
	// controller for andOp_276.andOp_276_in0
	// controller for andOp_276.andOp_276_in1
	// Insensitive connections
	always @(*) begin
		andOp_276_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_276_in1 = valid ? notOp_275_out : notOp_275_out;
	end
	// controller for andOp_278.andOp_278_in0
	// controller for andOp_278.andOp_278_in1
	// Insensitive connections
	always @(*) begin
		andOp_278_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_278_in1 = valid ? notOp_277_out : notOp_277_out;
	end
	// controller for andOp_279.andOp_279_in0
	// controller for andOp_279.andOp_279_in1
	// Insensitive connections
	always @(*) begin
		andOp_279_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_279_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_281.andOp_281_in0
	// controller for andOp_281.andOp_281_in1
	// Insensitive connections
	always @(*) begin
		andOp_281_in0 = valid ? andOp_279_out : andOp_279_out;
		andOp_281_in1 = valid ? eq_280_out : eq_280_out;
	end
	// controller for andOp_283.andOp_283_in0
	// controller for andOp_283.andOp_283_in1
	// Insensitive connections
	always @(*) begin
		andOp_283_in0 = valid ? andOp_279_out : andOp_279_out;
		andOp_283_in1 = valid ? notOp_282_out : notOp_282_out;
	end
	// controller for andOp_285.andOp_285_in0
	// controller for andOp_285.andOp_285_in1
	// Insensitive connections
	always @(*) begin
		andOp_285_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_285_in1 = valid ? notOp_284_out : notOp_284_out;
	end
	// controller for andOp_287.andOp_287_in0
	// controller for andOp_287.andOp_287_in1
	// Insensitive connections
	always @(*) begin
		andOp_287_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_287_in1 = valid ? notOp_286_out : notOp_286_out;
	end
	// controller for andOp_288.andOp_288_in0
	// controller for andOp_288.andOp_288_in1
	// Insensitive connections
	always @(*) begin
		andOp_288_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_288_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_290.andOp_290_in0
	// controller for andOp_290.andOp_290_in1
	// Insensitive connections
	always @(*) begin
		andOp_290_in0 = valid ? andOp_288_out : andOp_288_out;
		andOp_290_in1 = valid ? eq_289_out : eq_289_out;
	end
	// controller for andOp_292.andOp_292_in0
	// controller for andOp_292.andOp_292_in1
	// Insensitive connections
	always @(*) begin
		andOp_292_in0 = valid ? andOp_288_out : andOp_288_out;
		andOp_292_in1 = valid ? notOp_291_out : notOp_291_out;
	end
	// controller for andOp_294.andOp_294_in0
	// controller for andOp_294.andOp_294_in1
	// Insensitive connections
	always @(*) begin
		andOp_294_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_294_in1 = valid ? notOp_293_out : notOp_293_out;
	end
	// controller for andOp_296.andOp_296_in0
	// controller for andOp_296.andOp_296_in1
	// Insensitive connections
	always @(*) begin
		andOp_296_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_296_in1 = valid ? notOp_295_out : notOp_295_out;
	end
	// controller for andOp_299.andOp_299_in0
	// controller for andOp_299.andOp_299_in1
	// Insensitive connections
	always @(*) begin
		andOp_299_in0 = valid ? 1'd0 : 1'd0;
		andOp_299_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_301.andOp_301_in0
	// controller for andOp_301.andOp_301_in1
	// Insensitive connections
	always @(*) begin
		andOp_301_in0 = valid ? andOp_299_out : andOp_299_out;
		andOp_301_in1 = valid ? eq_300_out : eq_300_out;
	end
	// controller for andOp_303.andOp_303_in0
	// controller for andOp_303.andOp_303_in1
	// Insensitive connections
	always @(*) begin
		andOp_303_in0 = valid ? andOp_299_out : andOp_299_out;
		andOp_303_in1 = valid ? notOp_302_out : notOp_302_out;
	end
	// controller for andOp_305.andOp_305_in0
	// controller for andOp_305.andOp_305_in1
	// Insensitive connections
	always @(*) begin
		andOp_305_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_305_in1 = valid ? notOp_304_out : notOp_304_out;
	end
	// controller for andOp_307.andOp_307_in0
	// controller for andOp_307.andOp_307_in1
	// Insensitive connections
	always @(*) begin
		andOp_307_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_307_in1 = valid ? notOp_306_out : notOp_306_out;
	end
	// controller for andOp_308.andOp_308_in0
	// controller for andOp_308.andOp_308_in1
	// Insensitive connections
	always @(*) begin
		andOp_308_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_308_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_310.andOp_310_in0
	// controller for andOp_310.andOp_310_in1
	// Insensitive connections
	always @(*) begin
		andOp_310_in0 = valid ? andOp_308_out : andOp_308_out;
		andOp_310_in1 = valid ? eq_309_out : eq_309_out;
	end
	// controller for andOp_312.andOp_312_in0
	// controller for andOp_312.andOp_312_in1
	// Insensitive connections
	always @(*) begin
		andOp_312_in0 = valid ? andOp_308_out : andOp_308_out;
		andOp_312_in1 = valid ? notOp_311_out : notOp_311_out;
	end
	// controller for andOp_314.andOp_314_in0
	// controller for andOp_314.andOp_314_in1
	// Insensitive connections
	always @(*) begin
		andOp_314_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_314_in1 = valid ? notOp_313_out : notOp_313_out;
	end
	// controller for andOp_316.andOp_316_in0
	// controller for andOp_316.andOp_316_in1
	// Insensitive connections
	always @(*) begin
		andOp_316_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_316_in1 = valid ? notOp_315_out : notOp_315_out;
	end
	// controller for andOp_317.andOp_317_in0
	// controller for andOp_317.andOp_317_in1
	// Insensitive connections
	always @(*) begin
		andOp_317_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_317_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_319.andOp_319_in0
	// controller for andOp_319.andOp_319_in1
	// Insensitive connections
	always @(*) begin
		andOp_319_in0 = valid ? andOp_317_out : andOp_317_out;
		andOp_319_in1 = valid ? eq_318_out : eq_318_out;
	end
	// controller for andOp_32.andOp_32_in0
	// controller for andOp_32.andOp_32_in1
	// Insensitive connections
	always @(*) begin
		andOp_32_in0 = valid ? bb_0_active_in_state_1_out_data : bb_0_active_in_state_1_out_data;
		andOp_32_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_321.andOp_321_in0
	// controller for andOp_321.andOp_321_in1
	// Insensitive connections
	always @(*) begin
		andOp_321_in0 = valid ? andOp_317_out : andOp_317_out;
		andOp_321_in1 = valid ? notOp_320_out : notOp_320_out;
	end
	// controller for andOp_323.andOp_323_in0
	// controller for andOp_323.andOp_323_in1
	// Insensitive connections
	always @(*) begin
		andOp_323_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_323_in1 = valid ? notOp_322_out : notOp_322_out;
	end
	// controller for andOp_325.andOp_325_in0
	// controller for andOp_325.andOp_325_in1
	// Insensitive connections
	always @(*) begin
		andOp_325_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_325_in1 = valid ? notOp_324_out : notOp_324_out;
	end
	// controller for andOp_326.andOp_326_in0
	// controller for andOp_326.andOp_326_in1
	// Insensitive connections
	always @(*) begin
		andOp_326_in0 = valid ? 1'd0 : 1'd0;
		andOp_326_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_328.andOp_328_in0
	// controller for andOp_328.andOp_328_in1
	// Insensitive connections
	always @(*) begin
		andOp_328_in0 = valid ? andOp_326_out : andOp_326_out;
		andOp_328_in1 = valid ? eq_327_out : eq_327_out;
	end
	// controller for andOp_33.andOp_33_in0
	// controller for andOp_33.andOp_33_in1
	// Insensitive connections
	always @(*) begin
		andOp_33_in0 = valid ? andOp_32_out : andOp_32_out;
		andOp_33_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_330.andOp_330_in0
	// controller for andOp_330.andOp_330_in1
	// Insensitive connections
	always @(*) begin
		andOp_330_in0 = valid ? andOp_326_out : andOp_326_out;
		andOp_330_in1 = valid ? notOp_329_out : notOp_329_out;
	end
	// controller for andOp_332.andOp_332_in0
	// controller for andOp_332.andOp_332_in1
	// Insensitive connections
	always @(*) begin
		andOp_332_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_332_in1 = valid ? notOp_331_out : notOp_331_out;
	end
	// controller for andOp_334.andOp_334_in0
	// controller for andOp_334.andOp_334_in1
	// Insensitive connections
	always @(*) begin
		andOp_334_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_334_in1 = valid ? notOp_333_out : notOp_333_out;
	end
	// controller for andOp_35.andOp_35_in0
	// controller for andOp_35.andOp_35_in1
	// Insensitive connections
	always @(*) begin
		andOp_35_in0 = valid ? bb_0_active_in_state_1_out_data : bb_0_active_in_state_1_out_data;
		andOp_35_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_36.andOp_36_in0
	// controller for andOp_36.andOp_36_in1
	// Insensitive connections
	always @(*) begin
		andOp_36_in0 = valid ? andOp_35_out : andOp_35_out;
		andOp_36_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_38.andOp_38_in0
	// controller for andOp_38.andOp_38_in1
	// Insensitive connections
	always @(*) begin
		andOp_38_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_38_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_39.andOp_39_in0
	// controller for andOp_39.andOp_39_in1
	// Insensitive connections
	always @(*) begin
		andOp_39_in0 = valid ? andOp_38_out : andOp_38_out;
		andOp_39_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_41.andOp_41_in0
	// controller for andOp_41.andOp_41_in1
	// Insensitive connections
	always @(*) begin
		andOp_41_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
		andOp_41_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_42.andOp_42_in0
	// controller for andOp_42.andOp_42_in1
	// Insensitive connections
	always @(*) begin
		andOp_42_in0 = valid ? andOp_41_out : andOp_41_out;
		andOp_42_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_44.andOp_44_in0
	// controller for andOp_44.andOp_44_in1
	// Insensitive connections
	always @(*) begin
		andOp_44_in0 = valid ? andOp_42_out : andOp_42_out;
		andOp_44_in1 = valid ? in_read_ready : in_read_ready;
	end
	// controller for andOp_46.andOp_46_in0
	// controller for andOp_46.andOp_46_in1
	// Insensitive connections
	always @(*) begin
		andOp_46_in0 = valid ? andOp_42_out : andOp_42_out;
		andOp_46_in1 = valid ? notOp_45_out : notOp_45_out;
	end
	// controller for andOp_47.andOp_47_in0
	// controller for andOp_47.andOp_47_in1
	// Insensitive connections
	always @(*) begin
		andOp_47_in0 = valid ? bb_8_active_in_state_1_out_data : bb_8_active_in_state_1_out_data;
		andOp_47_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_48.andOp_48_in0
	// controller for andOp_48.andOp_48_in1
	// Insensitive connections
	always @(*) begin
		andOp_48_in0 = valid ? andOp_47_out : andOp_47_out;
		andOp_48_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_50.andOp_50_in0
	// controller for andOp_50.andOp_50_in1
	// Insensitive connections
	always @(*) begin
		andOp_50_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_50_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_51.andOp_51_in0
	// controller for andOp_51.andOp_51_in1
	// Insensitive connections
	always @(*) begin
		andOp_51_in0 = valid ? andOp_50_out : andOp_50_out;
		andOp_51_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_53.andOp_53_in0
	// controller for andOp_53.andOp_53_in1
	// Insensitive connections
	always @(*) begin
		andOp_53_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_53_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_54.andOp_54_in0
	// controller for andOp_54.andOp_54_in1
	// Insensitive connections
	always @(*) begin
		andOp_54_in0 = valid ? andOp_53_out : andOp_53_out;
		andOp_54_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_56.andOp_56_in0
	// controller for andOp_56.andOp_56_in1
	// Insensitive connections
	always @(*) begin
		andOp_56_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_56_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_57.andOp_57_in0
	// controller for andOp_57.andOp_57_in1
	// Insensitive connections
	always @(*) begin
		andOp_57_in0 = valid ? andOp_56_out : andOp_56_out;
		andOp_57_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_59.andOp_59_in0
	// controller for andOp_59.andOp_59_in1
	// Insensitive connections
	always @(*) begin
		andOp_59_in0 = valid ? andOp_57_out : andOp_57_out;
		andOp_59_in1 = valid ? data_in_4_29_out_data : data_in_4_29_out_data;
	end
	// controller for andOp_61.andOp_61_in0
	// controller for andOp_61.andOp_61_in1
	// Insensitive connections
	always @(*) begin
		andOp_61_in0 = valid ? andOp_57_out : andOp_57_out;
		andOp_61_in1 = valid ? notOp_60_out : notOp_60_out;
	end
	// controller for andOp_62.andOp_62_in0
	// controller for andOp_62.andOp_62_in1
	// Insensitive connections
	always @(*) begin
		andOp_62_in0 = valid ? bb_1_active_in_state_4_out_data : bb_1_active_in_state_4_out_data;
		andOp_62_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_63.andOp_63_in0
	// controller for andOp_63.andOp_63_in1
	// Insensitive connections
	always @(*) begin
		andOp_63_in0 = valid ? andOp_62_out : andOp_62_out;
		andOp_63_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_65.andOp_65_in0
	// controller for andOp_65.andOp_65_in1
	// Insensitive connections
	always @(*) begin
		andOp_65_in0 = valid ? bb_5_active_in_state_4_out_data : bb_5_active_in_state_4_out_data;
		andOp_65_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_66.andOp_66_in0
	// controller for andOp_66.andOp_66_in1
	// Insensitive connections
	always @(*) begin
		andOp_66_in0 = valid ? andOp_65_out : andOp_65_out;
		andOp_66_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_68.andOp_68_in0
	// controller for andOp_68.andOp_68_in1
	// Insensitive connections
	always @(*) begin
		andOp_68_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
		andOp_68_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_69.andOp_69_in0
	// controller for andOp_69.andOp_69_in1
	// Insensitive connections
	always @(*) begin
		andOp_69_in0 = valid ? andOp_68_out : andOp_68_out;
		andOp_69_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_71.andOp_71_in0
	// controller for andOp_71.andOp_71_in1
	// Insensitive connections
	always @(*) begin
		andOp_71_in0 = valid ? andOp_69_out : andOp_69_out;
		andOp_71_in1 = valid ? out_write_ready : out_write_ready;
	end
	// controller for andOp_73.andOp_73_in0
	// controller for andOp_73.andOp_73_in1
	// Insensitive connections
	always @(*) begin
		andOp_73_in0 = valid ? andOp_69_out : andOp_69_out;
		andOp_73_in1 = valid ? notOp_72_out : notOp_72_out;
	end
	// controller for andOp_74.andOp_74_in0
	// controller for andOp_74.andOp_74_in1
	// Insensitive connections
	always @(*) begin
		andOp_74_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_74_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_75.andOp_75_in0
	// controller for andOp_75.andOp_75_in1
	// Insensitive connections
	always @(*) begin
		andOp_75_in0 = valid ? andOp_74_out : andOp_74_out;
		andOp_75_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_77.andOp_77_in0
	// controller for andOp_77.andOp_77_in1
	// Insensitive connections
	always @(*) begin
		andOp_77_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_77_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_78.andOp_78_in0
	// controller for andOp_78.andOp_78_in1
	// Insensitive connections
	always @(*) begin
		andOp_78_in0 = valid ? andOp_77_out : andOp_77_out;
		andOp_78_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_80.andOp_80_in0
	// controller for andOp_80.andOp_80_in1
	// Insensitive connections
	always @(*) begin
		andOp_80_in0 = valid ? andOp_78_out : andOp_78_out;
		andOp_80_in1 = valid ? data_in_4_29_out_data : data_in_4_29_out_data;
	end
	// controller for andOp_82.andOp_82_in0
	// controller for andOp_82.andOp_82_in1
	// Insensitive connections
	always @(*) begin
		andOp_82_in0 = valid ? andOp_78_out : andOp_78_out;
		andOp_82_in1 = valid ? notOp_81_out : notOp_81_out;
	end
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_83_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_active_in_state_1.bb_0_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_1_in_data = eq_84_out;
		end else begin
			bb_0_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_106_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_1.bb_0_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_107_out) begin 
			bb_0_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_2.bb_10_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_2_in_data = eq_91_out;
		end else begin
			bb_10_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_3.bb_10_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_3_in_data = eq_92_out;
		end else begin
			bb_10_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_2.bb_10_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_117_out) begin 
			bb_10_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_3.bb_10_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_118_out) begin 
			bb_10_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_4.bb_1_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_4_in_data = orOp_96_out;
		end else begin
			bb_1_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_4.bb_1_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_124_out) begin 
			bb_1_predecessor_in_state_4_in_data = 32'd4;
		end else if (eq_122_out) begin 
			bb_1_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_4.bb_2_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_4_in_data = orOp_98_out;
		end else begin
			bb_2_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_4.bb_2_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_127_out) begin 
			bb_2_predecessor_in_state_4_in_data = 32'd7;
		end else if (eq_125_out) begin 
			bb_2_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_1.bb_3_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_1_in_data = orOp_86_out;
		end else begin
			bb_3_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_1.bb_3_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_110_out) begin 
			bb_3_predecessor_in_state_1_in_data = 32'd0;
		end else if (eq_108_out) begin 
			bb_3_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_3.bb_4_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_3_in_data = orOp_94_out;
		end else begin
			bb_4_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_4.bb_4_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_4_in_data = eq_105_out;
		end else begin
			bb_4_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_3.bb_4_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_121_out) begin 
			bb_4_predecessor_in_state_3_in_data = 32'd10;
		end else if (eq_119_out) begin 
			bb_4_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_4.bb_4_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_137_out) begin 
			bb_4_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_5_active_in_state_4.bb_5_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_5_active_in_state_4_in_data = orOp_100_out;
		end else begin
			bb_5_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_5_predecessor_in_state_4.bb_5_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_130_out) begin 
			bb_5_predecessor_in_state_4_in_data = 32'd1;
		end else if (eq_128_out) begin 
			bb_5_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_5_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_6_active_in_state_4.bb_6_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_6_active_in_state_4_in_data = orOp_102_out;
		end else begin
			bb_6_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_6_predecessor_in_state_4.bb_6_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_133_out) begin 
			bb_6_predecessor_in_state_4_in_data = 32'd5;
		end else if (eq_131_out) begin 
			bb_6_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_6_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_7_active_in_state_4.bb_7_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_7_active_in_state_4_in_data = orOp_104_out;
		end else begin
			bb_7_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_7_predecessor_in_state_4.bb_7_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_136_out) begin 
			bb_7_predecessor_in_state_4_in_data = 32'd6;
		end else if (eq_134_out) begin 
			bb_7_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_7_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_8_active_in_state_1.bb_8_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_state_1_in_data = orOp_90_out;
		end else begin
			bb_8_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_8_predecessor_in_state_1.bb_8_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_116_out) begin 
			bb_8_predecessor_in_state_1_in_data = 32'd3;
		end else if (eq_114_out) begin 
			bb_8_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_8_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_9_active_in_state_1.bb_9_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_9_active_in_state_1_in_data = orOp_88_out;
		end else begin
			bb_9_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_9_predecessor_in_state_1.bb_9_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_113_out) begin 
			bb_9_predecessor_in_state_1_in_data = 32'd8;
		end else if (eq_111_out) begin 
			bb_9_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_9_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_33_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_34_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_1.br_0_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_36_out) begin 
			br_0_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_37_out) begin 
			br_0_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_2.br_10_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_51_out) begin 
			br_10_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_52_out) begin 
			br_10_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_3.br_10_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_54_out) begin 
			br_10_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_55_out) begin 
			br_10_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_1_happened_in_state_4.br_1_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_63_out) begin 
			br_1_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_64_out) begin 
			br_1_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_1_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_1.br_3_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_39_out) begin 
			br_3_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_40_out) begin 
			br_3_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_3.br_4_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_57_out) begin 
			br_4_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_58_out) begin 
			br_4_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_4.br_4_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_78_out) begin 
			br_4_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_79_out) begin 
			br_4_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_5_happened_in_state_4.br_5_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_66_out) begin 
			br_5_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_67_out) begin 
			br_5_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_5_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_6_happened_in_state_4.br_6_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_69_out) begin 
			br_6_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_70_out) begin 
			br_6_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_6_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_7_happened_in_state_4.br_7_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_75_out) begin 
			br_7_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_76_out) begin 
			br_7_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_7_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_8_happened_in_state_1.br_8_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_48_out) begin 
			br_8_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_49_out) begin 
			br_8_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_8_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_9_happened_in_state_1.br_9_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_42_out) begin 
			br_9_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_43_out) begin 
			br_9_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_9_happened_in_state_1_in_data = 0;
		end
	end
	// controller for concat_146.concat_146_in0
	// controller for concat_146.concat_146_in1
	// Insensitive connections
	always @(*) begin
		concat_146_in0 = valid ? data_in_1_3_out_data : data_in_1_3_out_data;
		concat_146_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for concat_147.concat_147_in0
	// controller for concat_147.concat_147_in1
	// Insensitive connections
	always @(*) begin
		concat_147_in0 = valid ? 32'd4 : 32'd4;
		concat_147_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for data_in_1_1.data_in_1_1_in_data
	always @(*) begin
		if (eq_182_out) begin 
			data_in_1_1_in_data = 32'd0;
		end else if (eq_183_out) begin 
			data_in_1_1_in_data = data_store_1_0;
		end else if (eq_184_out) begin 
			data_in_1_1_in_data = data_store_4_24;
		end else begin
			data_in_1_1_in_data = 0;
		end
	end
	// controller for data_in_1_3.data_in_1_3_in_data
	always @(*) begin
		if (eq_182_out) begin 
			data_in_1_3_in_data = 32'd0;
		end else if (eq_183_out) begin 
			data_in_1_3_in_data = data_store_1_2;
		end else if (eq_184_out) begin 
			data_in_1_3_in_data = data_store_4_26;
		end else begin
			data_in_1_3_in_data = 0;
		end
	end
	// controller for data_in_1_5.data_in_1_5_in_data
	always @(*) begin
		if (eq_182_out) begin 
			data_in_1_5_in_data = 1'd0;
		end else if (eq_183_out) begin 
			data_in_1_5_in_data = data_store_1_4;
		end else if (eq_184_out) begin 
			data_in_1_5_in_data = data_store_4_28;
		end else begin
			data_in_1_5_in_data = 0;
		end
	end
	// controller for data_in_1_7.data_in_1_7_in_data
	always @(*) begin
		if (eq_182_out) begin 
			data_in_1_7_in_data = 32'd0;
		end else if (eq_183_out) begin 
			data_in_1_7_in_data = data_store_1_6;
		end else if (eq_184_out) begin 
			data_in_1_7_in_data = data_store_4_30;
		end else begin
			data_in_1_7_in_data = 0;
		end
	end
	// controller for data_in_2_11.data_in_2_11_in_data
	always @(*) begin
		if (eq_221_out) begin 
			data_in_2_11_in_data = data_store_1_2;
		end else if (eq_222_out) begin 
			data_in_2_11_in_data = data_store_2_10;
		end else begin
			data_in_2_11_in_data = 0;
		end
	end
	// controller for data_in_2_13.data_in_2_13_in_data
	always @(*) begin
		if (eq_221_out) begin 
			data_in_2_13_in_data = data_store_1_4;
		end else if (eq_222_out) begin 
			data_in_2_13_in_data = data_store_2_12;
		end else begin
			data_in_2_13_in_data = 0;
		end
	end
	// controller for data_in_2_15.data_in_2_15_in_data
	always @(*) begin
		if (eq_221_out) begin 
			data_in_2_15_in_data = data_store_1_6;
		end else if (eq_222_out) begin 
			data_in_2_15_in_data = data_store_2_14;
		end else begin
			data_in_2_15_in_data = 0;
		end
	end
	// controller for data_in_2_9.data_in_2_9_in_data
	always @(*) begin
		if (eq_221_out) begin 
			data_in_2_9_in_data = data_store_1_0;
		end else if (eq_222_out) begin 
			data_in_2_9_in_data = data_store_2_8;
		end else begin
			data_in_2_9_in_data = 0;
		end
	end
	// controller for data_in_3_17.data_in_3_17_in_data
	always @(*) begin
		if (eq_259_out) begin 
			data_in_3_17_in_data = data_store_2_8;
		end else if (eq_260_out) begin 
			data_in_3_17_in_data = data_store_3_16;
		end else begin
			data_in_3_17_in_data = 0;
		end
	end
	// controller for data_in_3_19.data_in_3_19_in_data
	always @(*) begin
		if (eq_259_out) begin 
			data_in_3_19_in_data = data_store_2_10;
		end else if (eq_260_out) begin 
			data_in_3_19_in_data = data_store_3_18;
		end else begin
			data_in_3_19_in_data = 0;
		end
	end
	// controller for data_in_3_21.data_in_3_21_in_data
	always @(*) begin
		if (eq_259_out) begin 
			data_in_3_21_in_data = data_store_2_12;
		end else if (eq_260_out) begin 
			data_in_3_21_in_data = data_store_3_20;
		end else begin
			data_in_3_21_in_data = 0;
		end
	end
	// controller for data_in_3_23.data_in_3_23_in_data
	always @(*) begin
		if (eq_259_out) begin 
			data_in_3_23_in_data = data_store_2_14;
		end else if (eq_260_out) begin 
			data_in_3_23_in_data = data_store_3_22;
		end else begin
			data_in_3_23_in_data = 0;
		end
	end
	// controller for data_in_4_25.data_in_4_25_in_data
	always @(*) begin
		if (eq_297_out) begin 
			data_in_4_25_in_data = data_store_3_16;
		end else if (eq_298_out) begin 
			data_in_4_25_in_data = data_store_4_24;
		end else begin
			data_in_4_25_in_data = 0;
		end
	end
	// controller for data_in_4_27.data_in_4_27_in_data
	always @(*) begin
		if (eq_297_out) begin 
			data_in_4_27_in_data = data_store_3_18;
		end else if (eq_298_out) begin 
			data_in_4_27_in_data = data_store_4_26;
		end else begin
			data_in_4_27_in_data = 0;
		end
	end
	// controller for data_in_4_29.data_in_4_29_in_data
	always @(*) begin
		if (eq_297_out) begin 
			data_in_4_29_in_data = data_store_3_20;
		end else if (eq_298_out) begin 
			data_in_4_29_in_data = data_store_4_28;
		end else begin
			data_in_4_29_in_data = 0;
		end
	end
	// controller for data_in_4_31.data_in_4_31_in_data
	always @(*) begin
		if (eq_297_out) begin 
			data_in_4_31_in_data = data_store_3_22;
		end else if (eq_298_out) begin 
			data_in_4_31_in_data = data_store_4_30;
		end else begin
			data_in_4_31_in_data = 0;
		end
	end
	// controller for eq_101.eq_101_in0
	// controller for eq_101.eq_101_in1
	// Insensitive connections
	always @(*) begin
		eq_101_in0 = valid ? 32'd6 : 32'd6;
		eq_101_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_103.eq_103_in0
	// controller for eq_103.eq_103_in1
	// Insensitive connections
	always @(*) begin
		eq_103_in0 = valid ? 32'd7 : 32'd7;
		eq_103_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_105.eq_105_in0
	// controller for eq_105.eq_105_in1
	// Insensitive connections
	always @(*) begin
		eq_105_in0 = valid ? 32'd4 : 32'd4;
		eq_105_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_106.eq_106_in0
	// controller for eq_106.eq_106_in1
	// Insensitive connections
	always @(*) begin
		eq_106_in0 = valid ? 32'd0 : 32'd0;
		eq_106_in1 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
	end
	// controller for eq_107.eq_107_in0
	// controller for eq_107.eq_107_in1
	// Insensitive connections
	always @(*) begin
		eq_107_in0 = valid ? 32'd0 : 32'd0;
		eq_107_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_108.eq_108_in0
	// controller for eq_108.eq_108_in1
	// Insensitive connections
	always @(*) begin
		eq_108_in0 = valid ? 32'd3 : 32'd3;
		eq_108_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_111.eq_111_in0
	// controller for eq_111.eq_111_in1
	// Insensitive connections
	always @(*) begin
		eq_111_in0 = valid ? 32'd9 : 32'd9;
		eq_111_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_114.eq_114_in0
	// controller for eq_114.eq_114_in1
	// Insensitive connections
	always @(*) begin
		eq_114_in0 = valid ? 32'd8 : 32'd8;
		eq_114_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_117.eq_117_in0
	// controller for eq_117.eq_117_in1
	// Insensitive connections
	always @(*) begin
		eq_117_in0 = valid ? 32'd10 : 32'd10;
		eq_117_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_118.eq_118_in0
	// controller for eq_118.eq_118_in1
	// Insensitive connections
	always @(*) begin
		eq_118_in0 = valid ? 32'd10 : 32'd10;
		eq_118_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_119.eq_119_in0
	// controller for eq_119.eq_119_in1
	// Insensitive connections
	always @(*) begin
		eq_119_in0 = valid ? 32'd4 : 32'd4;
		eq_119_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_122.eq_122_in0
	// controller for eq_122.eq_122_in1
	// Insensitive connections
	always @(*) begin
		eq_122_in0 = valid ? 32'd1 : 32'd1;
		eq_122_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_125.eq_125_in0
	// controller for eq_125.eq_125_in1
	// Insensitive connections
	always @(*) begin
		eq_125_in0 = valid ? 32'd2 : 32'd2;
		eq_125_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_128.eq_128_in0
	// controller for eq_128.eq_128_in1
	// Insensitive connections
	always @(*) begin
		eq_128_in0 = valid ? 32'd5 : 32'd5;
		eq_128_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_131.eq_131_in0
	// controller for eq_131.eq_131_in1
	// Insensitive connections
	always @(*) begin
		eq_131_in0 = valid ? 32'd6 : 32'd6;
		eq_131_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_134.eq_134_in0
	// controller for eq_134.eq_134_in1
	// Insensitive connections
	always @(*) begin
		eq_134_in0 = valid ? 32'd7 : 32'd7;
		eq_134_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_137.eq_137_in0
	// controller for eq_137.eq_137_in1
	// Insensitive connections
	always @(*) begin
		eq_137_in0 = valid ? 32'd4 : 32'd4;
		eq_137_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_153.eq_153_in0
	// controller for eq_153.eq_153_in1
	// Insensitive connections
	always @(*) begin
		eq_153_in0 = valid ? 32'd10 : 32'd10;
		eq_153_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_181.eq_181_in0
	// controller for eq_181.eq_181_in1
	// Insensitive connections
	always @(*) begin
		eq_181_in0 = valid ? 32'd0 : 32'd0;
		eq_181_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_182.eq_182_in0
	// controller for eq_182.eq_182_in1
	// Insensitive connections
	always @(*) begin
		eq_182_in0 = valid ? 32'd0 : 32'd0;
		eq_182_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_183.eq_183_in0
	// controller for eq_183.eq_183_in1
	// Insensitive connections
	always @(*) begin
		eq_183_in0 = valid ? 32'd1 : 32'd1;
		eq_183_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_184.eq_184_in0
	// controller for eq_184.eq_184_in1
	// Insensitive connections
	always @(*) begin
		eq_184_in0 = valid ? 32'd4 : 32'd4;
		eq_184_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_186.eq_186_in0
	// controller for eq_186.eq_186_in1
	// Insensitive connections
	always @(*) begin
		eq_186_in0 = valid ? 32'd1 : 32'd1;
		eq_186_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_195.eq_195_in0
	// controller for eq_195.eq_195_in1
	// Insensitive connections
	always @(*) begin
		eq_195_in0 = valid ? 32'd3 : 32'd3;
		eq_195_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_204.eq_204_in0
	// controller for eq_204.eq_204_in1
	// Insensitive connections
	always @(*) begin
		eq_204_in0 = valid ? 32'd3 : 32'd3;
		eq_204_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_213.eq_213_in0
	// controller for eq_213.eq_213_in1
	// Insensitive connections
	always @(*) begin
		eq_213_in0 = valid ? 32'd3 : 32'd3;
		eq_213_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_221.eq_221_in0
	// controller for eq_221.eq_221_in1
	// Insensitive connections
	always @(*) begin
		eq_221_in0 = valid ? 32'd1 : 32'd1;
		eq_221_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_222.eq_222_in0
	// controller for eq_222.eq_222_in1
	// Insensitive connections
	always @(*) begin
		eq_222_in0 = valid ? 32'd2 : 32'd2;
		eq_222_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_224.eq_224_in0
	// controller for eq_224.eq_224_in1
	// Insensitive connections
	always @(*) begin
		eq_224_in0 = valid ? 32'd1 : 32'd1;
		eq_224_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_233.eq_233_in0
	// controller for eq_233.eq_233_in1
	// Insensitive connections
	always @(*) begin
		eq_233_in0 = valid ? 32'd3 : 32'd3;
		eq_233_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_242.eq_242_in0
	// controller for eq_242.eq_242_in1
	// Insensitive connections
	always @(*) begin
		eq_242_in0 = valid ? 32'd3 : 32'd3;
		eq_242_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_251.eq_251_in0
	// controller for eq_251.eq_251_in1
	// Insensitive connections
	always @(*) begin
		eq_251_in0 = valid ? 32'd3 : 32'd3;
		eq_251_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_259.eq_259_in0
	// controller for eq_259.eq_259_in1
	// Insensitive connections
	always @(*) begin
		eq_259_in0 = valid ? 32'd2 : 32'd2;
		eq_259_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_260.eq_260_in0
	// controller for eq_260.eq_260_in1
	// Insensitive connections
	always @(*) begin
		eq_260_in0 = valid ? 32'd3 : 32'd3;
		eq_260_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_262.eq_262_in0
	// controller for eq_262.eq_262_in1
	// Insensitive connections
	always @(*) begin
		eq_262_in0 = valid ? 32'd1 : 32'd1;
		eq_262_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_271.eq_271_in0
	// controller for eq_271.eq_271_in1
	// Insensitive connections
	always @(*) begin
		eq_271_in0 = valid ? 32'd3 : 32'd3;
		eq_271_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_280.eq_280_in0
	// controller for eq_280.eq_280_in1
	// Insensitive connections
	always @(*) begin
		eq_280_in0 = valid ? 32'd3 : 32'd3;
		eq_280_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_289.eq_289_in0
	// controller for eq_289.eq_289_in1
	// Insensitive connections
	always @(*) begin
		eq_289_in0 = valid ? 32'd3 : 32'd3;
		eq_289_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_297.eq_297_in0
	// controller for eq_297.eq_297_in1
	// Insensitive connections
	always @(*) begin
		eq_297_in0 = valid ? 32'd3 : 32'd3;
		eq_297_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_298.eq_298_in0
	// controller for eq_298.eq_298_in1
	// Insensitive connections
	always @(*) begin
		eq_298_in0 = valid ? 32'd4 : 32'd4;
		eq_298_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_300.eq_300_in0
	// controller for eq_300.eq_300_in1
	// Insensitive connections
	always @(*) begin
		eq_300_in0 = valid ? 32'd1 : 32'd1;
		eq_300_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_309.eq_309_in0
	// controller for eq_309.eq_309_in1
	// Insensitive connections
	always @(*) begin
		eq_309_in0 = valid ? 32'd3 : 32'd3;
		eq_309_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_318.eq_318_in0
	// controller for eq_318.eq_318_in1
	// Insensitive connections
	always @(*) begin
		eq_318_in0 = valid ? 32'd3 : 32'd3;
		eq_318_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_327.eq_327_in0
	// controller for eq_327.eq_327_in1
	// Insensitive connections
	always @(*) begin
		eq_327_in0 = valid ? 32'd3 : 32'd3;
		eq_327_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_83.eq_83_in0
	// controller for eq_83.eq_83_in1
	// Insensitive connections
	always @(*) begin
		eq_83_in0 = valid ? 32'd0 : 32'd0;
		eq_83_in1 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
	end
	// controller for eq_84.eq_84_in0
	// controller for eq_84.eq_84_in1
	// Insensitive connections
	always @(*) begin
		eq_84_in0 = valid ? 32'd0 : 32'd0;
		eq_84_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_85.eq_85_in0
	// controller for eq_85.eq_85_in1
	// Insensitive connections
	always @(*) begin
		eq_85_in0 = valid ? 32'd3 : 32'd3;
		eq_85_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_87.eq_87_in0
	// controller for eq_87.eq_87_in1
	// Insensitive connections
	always @(*) begin
		eq_87_in0 = valid ? 32'd9 : 32'd9;
		eq_87_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_89.eq_89_in0
	// controller for eq_89.eq_89_in1
	// Insensitive connections
	always @(*) begin
		eq_89_in0 = valid ? 32'd8 : 32'd8;
		eq_89_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_91.eq_91_in0
	// controller for eq_91.eq_91_in1
	// Insensitive connections
	always @(*) begin
		eq_91_in0 = valid ? 32'd10 : 32'd10;
		eq_91_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_92.eq_92_in0
	// controller for eq_92.eq_92_in1
	// Insensitive connections
	always @(*) begin
		eq_92_in0 = valid ? 32'd10 : 32'd10;
		eq_92_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_93.eq_93_in0
	// controller for eq_93.eq_93_in1
	// Insensitive connections
	always @(*) begin
		eq_93_in0 = valid ? 32'd4 : 32'd4;
		eq_93_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_95.eq_95_in0
	// controller for eq_95.eq_95_in1
	// Insensitive connections
	always @(*) begin
		eq_95_in0 = valid ? 32'd1 : 32'd1;
		eq_95_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_97.eq_97_in0
	// controller for eq_97.eq_97_in1
	// Insensitive connections
	always @(*) begin
		eq_97_in0 = valid ? 32'd2 : 32'd2;
		eq_97_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_99.eq_99_in0
	// controller for eq_99.eq_99_in1
	// Insensitive connections
	always @(*) begin
		eq_99_in0 = valid ? 32'd5 : 32'd5;
		eq_99_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for icmp_15.cmp_in0_icmp_15
	// controller for icmp_15.cmp_in1_icmp_15
	// Insensitive connections
	always @(*) begin
		cmp_in0_icmp_15 = valid ? add_out_add_14 : add_out_add_14;
		cmp_in1_icmp_15 = valid ? 32'd4 : 32'd4;
	end
	// controller for in.in_read_valid_reg
	always @(*) begin
		if (andOp_149_out) begin 
			in_read_valid_reg = -(1'd1);
		end else begin
			in_read_valid_reg = 0;
		end
	end
	// controller for notOp_109.notOp_109_in0
	// Insensitive connections
	always @(*) begin
		notOp_109_in0 = valid ? eq_108_out : eq_108_out;
	end
	// controller for notOp_112.notOp_112_in0
	// Insensitive connections
	always @(*) begin
		notOp_112_in0 = valid ? eq_111_out : eq_111_out;
	end
	// controller for notOp_115.notOp_115_in0
	// Insensitive connections
	always @(*) begin
		notOp_115_in0 = valid ? eq_114_out : eq_114_out;
	end
	// controller for notOp_120.notOp_120_in0
	// Insensitive connections
	always @(*) begin
		notOp_120_in0 = valid ? eq_119_out : eq_119_out;
	end
	// controller for notOp_123.notOp_123_in0
	// Insensitive connections
	always @(*) begin
		notOp_123_in0 = valid ? eq_122_out : eq_122_out;
	end
	// controller for notOp_126.notOp_126_in0
	// Insensitive connections
	always @(*) begin
		notOp_126_in0 = valid ? eq_125_out : eq_125_out;
	end
	// controller for notOp_129.notOp_129_in0
	// Insensitive connections
	always @(*) begin
		notOp_129_in0 = valid ? eq_128_out : eq_128_out;
	end
	// controller for notOp_132.notOp_132_in0
	// Insensitive connections
	always @(*) begin
		notOp_132_in0 = valid ? eq_131_out : eq_131_out;
	end
	// controller for notOp_135.notOp_135_in0
	// Insensitive connections
	always @(*) begin
		notOp_135_in0 = valid ? eq_134_out : eq_134_out;
	end
	// controller for notOp_165.notOp_165_in0
	// Insensitive connections
	always @(*) begin
		notOp_165_in0 = valid ? andOp_161_out : andOp_161_out;
	end
	// controller for notOp_167.notOp_167_in0
	// Insensitive connections
	always @(*) begin
		notOp_167_in0 = valid ? andOp_46_out : andOp_46_out;
	end
	// controller for notOp_169.notOp_169_in0
	// Insensitive connections
	always @(*) begin
		notOp_169_in0 = valid ? andOp_61_out : andOp_61_out;
	end
	// controller for notOp_171.notOp_171_in0
	// Insensitive connections
	always @(*) begin
		notOp_171_in0 = valid ? andOp_44_out : andOp_44_out;
	end
	// controller for notOp_173.notOp_173_in0
	// Insensitive connections
	always @(*) begin
		notOp_173_in0 = valid ? andOp_162_out : andOp_162_out;
	end
	// controller for notOp_175.notOp_175_in0
	// Insensitive connections
	always @(*) begin
		notOp_175_in0 = valid ? andOp_163_out : andOp_163_out;
	end
	// controller for notOp_177.notOp_177_in0
	// Insensitive connections
	always @(*) begin
		notOp_177_in0 = valid ? andOp_164_out : andOp_164_out;
	end
	// controller for notOp_179.notOp_179_in0
	// Insensitive connections
	always @(*) begin
		notOp_179_in0 = valid ? andOp_73_out : andOp_73_out;
	end
	// controller for notOp_188.notOp_188_in0
	// Insensitive connections
	always @(*) begin
		notOp_188_in0 = valid ? eq_186_out : eq_186_out;
	end
	// controller for notOp_190.notOp_190_in0
	// Insensitive connections
	always @(*) begin
		notOp_190_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
	end
	// controller for notOp_192.notOp_192_in0
	// Insensitive connections
	always @(*) begin
		notOp_192_in0 = valid ? andOp_187_out : andOp_187_out;
	end
	// controller for notOp_197.notOp_197_in0
	// Insensitive connections
	always @(*) begin
		notOp_197_in0 = valid ? eq_195_out : eq_195_out;
	end
	// controller for notOp_199.notOp_199_in0
	// Insensitive connections
	always @(*) begin
		notOp_199_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_201.notOp_201_in0
	// Insensitive connections
	always @(*) begin
		notOp_201_in0 = valid ? andOp_196_out : andOp_196_out;
	end
	// controller for notOp_206.notOp_206_in0
	// Insensitive connections
	always @(*) begin
		notOp_206_in0 = valid ? eq_204_out : eq_204_out;
	end
	// controller for notOp_208.notOp_208_in0
	// Insensitive connections
	always @(*) begin
		notOp_208_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_210.notOp_210_in0
	// Insensitive connections
	always @(*) begin
		notOp_210_in0 = valid ? andOp_205_out : andOp_205_out;
	end
	// controller for notOp_215.notOp_215_in0
	// Insensitive connections
	always @(*) begin
		notOp_215_in0 = valid ? eq_213_out : eq_213_out;
	end
	// controller for notOp_217.notOp_217_in0
	// Insensitive connections
	always @(*) begin
		notOp_217_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_219.notOp_219_in0
	// Insensitive connections
	always @(*) begin
		notOp_219_in0 = valid ? andOp_214_out : andOp_214_out;
	end
	// controller for notOp_226.notOp_226_in0
	// Insensitive connections
	always @(*) begin
		notOp_226_in0 = valid ? eq_224_out : eq_224_out;
	end
	// controller for notOp_228.notOp_228_in0
	// Insensitive connections
	always @(*) begin
		notOp_228_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_230.notOp_230_in0
	// Insensitive connections
	always @(*) begin
		notOp_230_in0 = valid ? andOp_225_out : andOp_225_out;
	end
	// controller for notOp_235.notOp_235_in0
	// Insensitive connections
	always @(*) begin
		notOp_235_in0 = valid ? eq_233_out : eq_233_out;
	end
	// controller for notOp_237.notOp_237_in0
	// Insensitive connections
	always @(*) begin
		notOp_237_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_239.notOp_239_in0
	// Insensitive connections
	always @(*) begin
		notOp_239_in0 = valid ? andOp_234_out : andOp_234_out;
	end
	// controller for notOp_244.notOp_244_in0
	// Insensitive connections
	always @(*) begin
		notOp_244_in0 = valid ? eq_242_out : eq_242_out;
	end
	// controller for notOp_246.notOp_246_in0
	// Insensitive connections
	always @(*) begin
		notOp_246_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_248.notOp_248_in0
	// Insensitive connections
	always @(*) begin
		notOp_248_in0 = valid ? andOp_243_out : andOp_243_out;
	end
	// controller for notOp_253.notOp_253_in0
	// Insensitive connections
	always @(*) begin
		notOp_253_in0 = valid ? eq_251_out : eq_251_out;
	end
	// controller for notOp_255.notOp_255_in0
	// Insensitive connections
	always @(*) begin
		notOp_255_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
	end
	// controller for notOp_257.notOp_257_in0
	// Insensitive connections
	always @(*) begin
		notOp_257_in0 = valid ? andOp_252_out : andOp_252_out;
	end
	// controller for notOp_264.notOp_264_in0
	// Insensitive connections
	always @(*) begin
		notOp_264_in0 = valid ? eq_262_out : eq_262_out;
	end
	// controller for notOp_266.notOp_266_in0
	// Insensitive connections
	always @(*) begin
		notOp_266_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_268.notOp_268_in0
	// Insensitive connections
	always @(*) begin
		notOp_268_in0 = valid ? andOp_263_out : andOp_263_out;
	end
	// controller for notOp_273.notOp_273_in0
	// Insensitive connections
	always @(*) begin
		notOp_273_in0 = valid ? eq_271_out : eq_271_out;
	end
	// controller for notOp_275.notOp_275_in0
	// Insensitive connections
	always @(*) begin
		notOp_275_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
	end
	// controller for notOp_277.notOp_277_in0
	// Insensitive connections
	always @(*) begin
		notOp_277_in0 = valid ? andOp_272_out : andOp_272_out;
	end
	// controller for notOp_282.notOp_282_in0
	// Insensitive connections
	always @(*) begin
		notOp_282_in0 = valid ? eq_280_out : eq_280_out;
	end
	// controller for notOp_284.notOp_284_in0
	// Insensitive connections
	always @(*) begin
		notOp_284_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
	end
	// controller for notOp_286.notOp_286_in0
	// Insensitive connections
	always @(*) begin
		notOp_286_in0 = valid ? andOp_281_out : andOp_281_out;
	end
	// controller for notOp_291.notOp_291_in0
	// Insensitive connections
	always @(*) begin
		notOp_291_in0 = valid ? eq_289_out : eq_289_out;
	end
	// controller for notOp_293.notOp_293_in0
	// Insensitive connections
	always @(*) begin
		notOp_293_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
	end
	// controller for notOp_295.notOp_295_in0
	// Insensitive connections
	always @(*) begin
		notOp_295_in0 = valid ? andOp_290_out : andOp_290_out;
	end
	// controller for notOp_302.notOp_302_in0
	// Insensitive connections
	always @(*) begin
		notOp_302_in0 = valid ? eq_300_out : eq_300_out;
	end
	// controller for notOp_304.notOp_304_in0
	// Insensitive connections
	always @(*) begin
		notOp_304_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_306.notOp_306_in0
	// Insensitive connections
	always @(*) begin
		notOp_306_in0 = valid ? andOp_301_out : andOp_301_out;
	end
	// controller for notOp_311.notOp_311_in0
	// Insensitive connections
	always @(*) begin
		notOp_311_in0 = valid ? eq_309_out : eq_309_out;
	end
	// controller for notOp_313.notOp_313_in0
	// Insensitive connections
	always @(*) begin
		notOp_313_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
	end
	// controller for notOp_315.notOp_315_in0
	// Insensitive connections
	always @(*) begin
		notOp_315_in0 = valid ? andOp_310_out : andOp_310_out;
	end
	// controller for notOp_320.notOp_320_in0
	// Insensitive connections
	always @(*) begin
		notOp_320_in0 = valid ? eq_318_out : eq_318_out;
	end
	// controller for notOp_322.notOp_322_in0
	// Insensitive connections
	always @(*) begin
		notOp_322_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
	end
	// controller for notOp_324.notOp_324_in0
	// Insensitive connections
	always @(*) begin
		notOp_324_in0 = valid ? andOp_319_out : andOp_319_out;
	end
	// controller for notOp_329.notOp_329_in0
	// Insensitive connections
	always @(*) begin
		notOp_329_in0 = valid ? eq_327_out : eq_327_out;
	end
	// controller for notOp_331.notOp_331_in0
	// Insensitive connections
	always @(*) begin
		notOp_331_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_333.notOp_333_in0
	// Insensitive connections
	always @(*) begin
		notOp_333_in0 = valid ? andOp_328_out : andOp_328_out;
	end
	// controller for notOp_34.notOp_34_in0
	// Insensitive connections
	always @(*) begin
		notOp_34_in0 = valid ? andOp_33_out : andOp_33_out;
	end
	// controller for notOp_37.notOp_37_in0
	// Insensitive connections
	always @(*) begin
		notOp_37_in0 = valid ? andOp_36_out : andOp_36_out;
	end
	// controller for notOp_40.notOp_40_in0
	// Insensitive connections
	always @(*) begin
		notOp_40_in0 = valid ? andOp_39_out : andOp_39_out;
	end
	// controller for notOp_43.notOp_43_in0
	// Insensitive connections
	always @(*) begin
		notOp_43_in0 = valid ? andOp_42_out : andOp_42_out;
	end
	// controller for notOp_45.notOp_45_in0
	// Insensitive connections
	always @(*) begin
		notOp_45_in0 = valid ? in_read_ready : in_read_ready;
	end
	// controller for notOp_49.notOp_49_in0
	// Insensitive connections
	always @(*) begin
		notOp_49_in0 = valid ? andOp_48_out : andOp_48_out;
	end
	// controller for notOp_52.notOp_52_in0
	// Insensitive connections
	always @(*) begin
		notOp_52_in0 = valid ? andOp_51_out : andOp_51_out;
	end
	// controller for notOp_55.notOp_55_in0
	// Insensitive connections
	always @(*) begin
		notOp_55_in0 = valid ? andOp_54_out : andOp_54_out;
	end
	// controller for notOp_58.notOp_58_in0
	// Insensitive connections
	always @(*) begin
		notOp_58_in0 = valid ? andOp_57_out : andOp_57_out;
	end
	// controller for notOp_60.notOp_60_in0
	// Insensitive connections
	always @(*) begin
		notOp_60_in0 = valid ? data_in_4_29_out_data : data_in_4_29_out_data;
	end
	// controller for notOp_64.notOp_64_in0
	// Insensitive connections
	always @(*) begin
		notOp_64_in0 = valid ? andOp_63_out : andOp_63_out;
	end
	// controller for notOp_67.notOp_67_in0
	// Insensitive connections
	always @(*) begin
		notOp_67_in0 = valid ? andOp_66_out : andOp_66_out;
	end
	// controller for notOp_70.notOp_70_in0
	// Insensitive connections
	always @(*) begin
		notOp_70_in0 = valid ? andOp_69_out : andOp_69_out;
	end
	// controller for notOp_72.notOp_72_in0
	// Insensitive connections
	always @(*) begin
		notOp_72_in0 = valid ? out_write_ready : out_write_ready;
	end
	// controller for notOp_76.notOp_76_in0
	// Insensitive connections
	always @(*) begin
		notOp_76_in0 = valid ? andOp_75_out : andOp_75_out;
	end
	// controller for notOp_79.notOp_79_in0
	// Insensitive connections
	always @(*) begin
		notOp_79_in0 = valid ? andOp_78_out : andOp_78_out;
	end
	// controller for notOp_81.notOp_81_in0
	// Insensitive connections
	always @(*) begin
		notOp_81_in0 = valid ? data_in_4_29_out_data : data_in_4_29_out_data;
	end
	// controller for orOp_100.orOp_100_in0
	// controller for orOp_100.orOp_100_in1
	// Insensitive connections
	always @(*) begin
		orOp_100_in0 = valid ? eq_99_out : eq_99_out;
		orOp_100_in1 = valid ? andOp_63_out : andOp_63_out;
	end
	// controller for orOp_102.orOp_102_in0
	// controller for orOp_102.orOp_102_in1
	// Insensitive connections
	always @(*) begin
		orOp_102_in0 = valid ? eq_101_out : eq_101_out;
		orOp_102_in1 = valid ? andOp_66_out : andOp_66_out;
	end
	// controller for orOp_104.orOp_104_in0
	// controller for orOp_104.orOp_104_in1
	// Insensitive connections
	always @(*) begin
		orOp_104_in0 = valid ? eq_103_out : eq_103_out;
		orOp_104_in1 = valid ? andOp_71_out : andOp_71_out;
	end
	// controller for orOp_86.orOp_86_in0
	// controller for orOp_86.orOp_86_in1
	// Insensitive connections
	always @(*) begin
		orOp_86_in0 = valid ? eq_85_out : eq_85_out;
		orOp_86_in1 = valid ? andOp_33_out : andOp_33_out;
	end
	// controller for orOp_88.orOp_88_in0
	// controller for orOp_88.orOp_88_in1
	// Insensitive connections
	always @(*) begin
		orOp_88_in0 = valid ? eq_87_out : eq_87_out;
		orOp_88_in1 = valid ? andOp_48_out : andOp_48_out;
	end
	// controller for orOp_90.orOp_90_in0
	// controller for orOp_90.orOp_90_in1
	// Insensitive connections
	always @(*) begin
		orOp_90_in0 = valid ? eq_89_out : eq_89_out;
		orOp_90_in1 = valid ? andOp_39_out : andOp_39_out;
	end
	// controller for orOp_94.orOp_94_in0
	// controller for orOp_94.orOp_94_in1
	// Insensitive connections
	always @(*) begin
		orOp_94_in0 = valid ? eq_93_out : eq_93_out;
		orOp_94_in1 = valid ? andOp_51_out : andOp_51_out;
	end
	// controller for orOp_96.orOp_96_in0
	// controller for orOp_96.orOp_96_in1
	// Insensitive connections
	always @(*) begin
		orOp_96_in0 = valid ? eq_95_out : eq_95_out;
		orOp_96_in1 = valid ? andOp_59_out : andOp_59_out;
	end
	// controller for orOp_98.orOp_98_in0
	// controller for orOp_98.orOp_98_in1
	// Insensitive connections
	always @(*) begin
		orOp_98_in0 = valid ? eq_97_out : eq_97_out;
		orOp_98_in1 = valid ? andOp_75_out : andOp_75_out;
	end
	// controller for out.out_in_data_reg
	always @(*) begin
		if (andOp_159_out) begin 
			out_in_data_reg = rdata_ram_0;
		end else begin
			out_in_data_reg = 0;
		end
	end
	// controller for out.out_write_valid_reg
	always @(*) begin
		if (andOp_158_out) begin 
			out_write_valid_reg = -(1'd1);
		end else begin
			out_write_valid_reg = 0;
		end
	end
	// controller for phi_5.phi_in_phi_5
	// controller for phi_5.phi_last_block_phi_5
	// controller for phi_5.phi_s_phi_5
	// Insensitive connections
	always @(*) begin
		phi_in_phi_5 = valid ? concat_146_out : concat_146_out;
		phi_last_block_phi_5 = valid ? bb_3_predecessor_in_state_1_out_data : bb_3_predecessor_in_state_1_out_data;
		phi_s_phi_5 = valid ? concat_147_out : concat_147_out;
	end
	// controller for ram_0.raddr_ram_0_reg
	always @(*) begin
		if (andOp_142_out) begin 
			raddr_ram_0_reg = 32'd0;
		end else if (andOp_144_out) begin 
			raddr_ram_0_reg = 32'd0;
		end else begin
			raddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.waddr_ram_0_reg
	always @(*) begin
		if (andOp_141_out) begin 
			waddr_ram_0_reg = 32'd0;
		end else if (andOp_143_out) begin 
			waddr_ram_0_reg = 32'd0;
		end else begin
			waddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wdata_ram_0_reg
	always @(*) begin
		if (andOp_141_out) begin 
			wdata_ram_0_reg = 32'd0;
		end else if (andOp_143_out) begin 
			wdata_ram_0_reg = add_out_add_12;
		end else begin
			wdata_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wen_ram_0_reg
	always @(*) begin
		if (andOp_141_out) begin 
			wen_ram_0_reg = 1'd1;
		end else if (andOp_143_out) begin 
			wen_ram_0_reg = 1'd1;
		end else begin
			wen_ram_0_reg = 0;
		end
	end
	// controller for ret_19.valid_reg
	always @(*) begin
		if (andOp_157_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// controller for tmp_output_152.tmp_output_152_in_data
	always @(*) begin
		if (eq_153_out) begin 
			tmp_output_152_in_data = in_out_data;
		end else begin
			tmp_output_152_in_data = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			data_store_1_0 <= 0;
		end else begin
			if (andOp_187_out) begin
				data_store_1_0 <= phi_out_phi_5;
			end
			if (andOp_193_out) begin
				data_store_1_0 <= data_in_1_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_2 <= 0;
		end else begin
			if (andOp_196_out) begin
				data_store_1_2 <= add_out_add_14;
			end
			if (andOp_202_out) begin
				data_store_1_2 <= data_in_1_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_4 <= 0;
		end else begin
			if (andOp_205_out) begin
				data_store_1_4 <= cmp_out_icmp_15;
			end
			if (andOp_211_out) begin
				data_store_1_4 <= data_in_1_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_6 <= 0;
		end else begin
			if (andOp_214_out) begin
				data_store_1_6 <= in_out_data;
			end
			if (andOp_220_out) begin
				data_store_1_6 <= data_in_1_7_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_10 <= 0;
		end else begin
			if (andOp_234_out) begin
				data_store_2_10 <= add_out_add_14;
			end
			if (andOp_240_out) begin
				data_store_2_10 <= data_in_2_11_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_12 <= 0;
		end else begin
			if (andOp_243_out) begin
				data_store_2_12 <= cmp_out_icmp_15;
			end
			if (andOp_249_out) begin
				data_store_2_12 <= data_in_2_13_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_14 <= 0;
		end else begin
			if (andOp_252_out) begin
				data_store_2_14 <= in_out_data;
			end
			if (andOp_258_out) begin
				data_store_2_14 <= data_in_2_15_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_8 <= 0;
		end else begin
			if (andOp_225_out) begin
				data_store_2_8 <= phi_out_phi_5;
			end
			if (andOp_231_out) begin
				data_store_2_8 <= data_in_2_9_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_16 <= 0;
		end else begin
			if (andOp_263_out) begin
				data_store_3_16 <= phi_out_phi_5;
			end
			if (andOp_269_out) begin
				data_store_3_16 <= data_in_3_17_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_18 <= 0;
		end else begin
			if (andOp_272_out) begin
				data_store_3_18 <= add_out_add_14;
			end
			if (andOp_278_out) begin
				data_store_3_18 <= data_in_3_19_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_20 <= 0;
		end else begin
			if (andOp_281_out) begin
				data_store_3_20 <= cmp_out_icmp_15;
			end
			if (andOp_287_out) begin
				data_store_3_20 <= data_in_3_21_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_22 <= 0;
		end else begin
			if (andOp_290_out) begin
				data_store_3_22 <= in_out_data;
			end
			if (andOp_296_out) begin
				data_store_3_22 <= data_in_3_23_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_24 <= 0;
		end else begin
			if (andOp_301_out) begin
				data_store_4_24 <= phi_out_phi_5;
			end
			if (andOp_307_out) begin
				data_store_4_24 <= data_in_4_25_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_26 <= 0;
		end else begin
			if (andOp_310_out) begin
				data_store_4_26 <= add_out_add_14;
			end
			if (andOp_316_out) begin
				data_store_4_26 <= data_in_4_27_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_28 <= 0;
		end else begin
			if (andOp_319_out) begin
				data_store_4_28 <= cmp_out_icmp_15;
			end
			if (andOp_325_out) begin
				data_store_4_28 <= data_in_4_29_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_30 <= 0;
		end else begin
			if (andOp_328_out) begin
				data_store_4_30 <= in_out_data;
			end
			if (andOp_334_out) begin
				data_store_4_30 <= data_in_4_31_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_161_out) begin
				global_state <= 32'd1;
			end
			if (andOp_162_out) begin
				global_state <= 32'd3;
			end
			if (andOp_163_out) begin
				global_state <= 32'd4;
			end
			if (andOp_164_out) begin
				global_state <= 32'd4;
			end
			if (andOp_44_out) begin
				global_state <= 32'd2;
			end
			if (andOp_46_out) begin
				global_state <= 32'd1;
			end
			if (andOp_61_out) begin
				global_state <= 32'd1;
			end
			if (andOp_73_out) begin
				global_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (1'd1) begin
				state_0_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_161_out) begin
				state_1_entry_BB_reg <= 32'd0;
			end
			if (andOp_46_out) begin
				state_1_entry_BB_reg <= 32'd9;
			end
			if (andOp_61_out) begin
				state_1_entry_BB_reg <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_161_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_170_out) begin
				state_1_is_active <= 1'd0;
			end
			if (andOp_46_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_61_out) begin
				state_1_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_161_out) begin
				state_1_last_BB_reg <= bb_0_predecessor_in_state_0_out_data;
			end
			if (andOp_46_out) begin
				state_1_last_BB_reg <= 32'd9;
			end
			if (andOp_61_out) begin
				state_1_last_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_161_out) begin
				state_1_last_state <= 32'd0;
			end
			if (andOp_46_out) begin
				state_1_last_state <= 32'd1;
			end
			if (andOp_61_out) begin
				state_1_last_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_44_out) begin
				state_2_entry_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_172_out) begin
				state_2_is_active <= 1'd0;
			end
			if (andOp_44_out) begin
				state_2_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_44_out) begin
				state_2_last_BB_reg <= 32'd9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_44_out) begin
				state_2_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_162_out) begin
				state_3_entry_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_162_out) begin
				state_3_is_active <= 1'd1;
			end
			if (andOp_174_out) begin
				state_3_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_162_out) begin
				state_3_last_BB_reg <= bb_10_predecessor_in_state_2_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_state <= 0;
		end else begin
			if (andOp_162_out) begin
				state_3_last_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_163_out) begin
				state_4_entry_BB_reg <= 32'd4;
			end
			if (andOp_164_out) begin
				state_4_entry_BB_reg <= 32'd2;
			end
			if (andOp_73_out) begin
				state_4_entry_BB_reg <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_163_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_164_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_180_out) begin
				state_4_is_active <= 1'd0;
			end
			if (andOp_73_out) begin
				state_4_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_163_out) begin
				state_4_last_BB_reg <= bb_4_predecessor_in_state_3_out_data;
			end
			if (andOp_164_out) begin
				state_4_last_BB_reg <= bb_2_predecessor_in_state_4_out_data;
			end
			if (andOp_73_out) begin
				state_4_last_BB_reg <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_state <= 0;
		end else begin
			if (andOp_163_out) begin
				state_4_last_state <= 32'd3;
			end
			if (andOp_164_out) begin
				state_4_last_state <= 32'd4;
			end
			if (andOp_73_out) begin
				state_4_last_state <= 32'd4;
			end
		end
	end

endmodule

