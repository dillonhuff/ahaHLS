module channel_reduce_4(input [0:0] clk, input [0:0] rst, output [31:0] out_in_data, output [0:0] out_read_valid, output [0:0] out_rst, output [0:0] out_write_valid, input [31:0] out_out_data, input [0:0] out_read_ready, input [0:0] out_write_ready, output [31:0] in_in_data, output [0:0] in_read_valid, output [0:0] in_rst, output [0:0] in_write_valid, input [31:0] in_out_data, input [0:0] in_read_ready, input [0:0] in_write_ready, output [0:0] valid);

	reg [31:0] out_in_data_reg;
	reg [0:0] out_read_valid_reg;
	reg [0:0] out_rst_reg;
	reg [0:0] out_write_valid_reg;
	reg [31:0] in_in_data_reg;
	reg [0:0] in_read_valid_reg;
	reg [0:0] in_rst_reg;
	reg [0:0] in_write_valid_reg;
	reg [0:0] valid_reg;

	assign out_in_data = out_in_data_reg;
	assign out_read_valid = out_read_valid_reg;
	assign out_rst = out_rst_reg;
	assign out_write_valid = out_write_valid_reg;
	assign in_in_data = in_in_data_reg;
	assign in_read_valid = in_read_valid_reg;
	assign in_rst = in_rst_reg;
	assign in_write_valid = in_write_valid_reg;
	assign valid = valid_reg;

	// Start debug wires and ports

	initial begin
	end





	// End debug wires and ports

	// Start Functional Units
	br_dummy br_unit();

	reg [31:0] raddr_ram_0_reg;
	reg [31:0] waddr_ram_0_reg;
	reg [31:0] wdata_ram_0_reg;
	reg [0:0] wen_ram_0_reg;
	wire [31:0] rdata_ram_0;
	register #(.WIDTH(32)) ram_0(.clk(clk), .raddr(raddr_ram_0_reg), .rdata(rdata_ram_0), .rst(rst), .waddr(waddr_ram_0_reg), .wdata(wdata_ram_0_reg), .wen(wen_ram_0_reg));

	add alloca_0();

	add bitcast_1();

	add call_2();

	add call_26();

	reg [63:0] phi_in_phi_9;
	reg [31:0] phi_last_block_phi_9;
	reg [63:0] phi_s_phi_9;
	wire [31:0] phi_out_phi_9;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_9(.in(phi_in_phi_9), .last_block(phi_last_block_phi_9), .out(phi_out_phi_9), .s(phi_s_phi_9));

	reg [31:0] add_in0_add_14;
	reg [31:0] add_in1_add_14;
	wire [31:0] add_out_add_14;
	add #(.WIDTH(32)) add_add_14(.in0(add_in0_add_14), .in1(add_in1_add_14), .out(add_out_add_14));

	reg [31:0] add_in0_add_16;
	reg [31:0] add_in1_add_16;
	wire [31:0] add_out_add_16;
	add #(.WIDTH(32)) add_add_16(.in0(add_in0_add_16), .in1(add_in1_add_16), .out(add_out_add_16));

	reg [31:0] cmp_in0_icmp_17;
	reg [31:0] cmp_in1_icmp_17;
	wire [0:0] cmp_out_icmp_17;
	eq #(.WIDTH(32)) icmp_17(.in0(cmp_in0_icmp_17), .in1(cmp_in1_icmp_17), .out(cmp_out_icmp_17));

	reg [31:0] data_in_0_1_in_data;
	wire [31:0] data_in_0_1_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_1(.in_data(data_in_0_1_in_data), .out_data(data_in_0_1_out_data));

	reg [31:0] data_in_0_3_in_data;
	wire [31:0] data_in_0_3_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_3(.in_data(data_in_0_3_in_data), .out_data(data_in_0_3_out_data));

	reg [31:0] data_in_0_5_in_data;
	wire [31:0] data_in_0_5_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_5(.in_data(data_in_0_5_in_data), .out_data(data_in_0_5_out_data));

	reg [0:0] data_in_0_7_in_data;
	wire [0:0] data_in_0_7_out_data;
	hls_wire #(.WIDTH(1)) data_in_0_7(.in_data(data_in_0_7_in_data), .out_data(data_in_0_7_out_data));

	reg [31:0] data_in_1_9_in_data;
	wire [31:0] data_in_1_9_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_9(.in_data(data_in_1_9_in_data), .out_data(data_in_1_9_out_data));

	reg [31:0] data_in_1_11_in_data;
	wire [31:0] data_in_1_11_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_11(.in_data(data_in_1_11_in_data), .out_data(data_in_1_11_out_data));

	reg [31:0] data_in_1_13_in_data;
	wire [31:0] data_in_1_13_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_13(.in_data(data_in_1_13_in_data), .out_data(data_in_1_13_out_data));

	reg [0:0] data_in_1_15_in_data;
	wire [0:0] data_in_1_15_out_data;
	hls_wire #(.WIDTH(1)) data_in_1_15(.in_data(data_in_1_15_in_data), .out_data(data_in_1_15_out_data));

	reg [31:0] data_in_2_17_in_data;
	wire [31:0] data_in_2_17_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_17(.in_data(data_in_2_17_in_data), .out_data(data_in_2_17_out_data));

	reg [31:0] data_in_2_19_in_data;
	wire [31:0] data_in_2_19_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_19(.in_data(data_in_2_19_in_data), .out_data(data_in_2_19_out_data));

	reg [31:0] data_in_2_21_in_data;
	wire [31:0] data_in_2_21_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_21(.in_data(data_in_2_21_in_data), .out_data(data_in_2_21_out_data));

	reg [0:0] data_in_2_23_in_data;
	wire [0:0] data_in_2_23_out_data;
	hls_wire #(.WIDTH(1)) data_in_2_23(.in_data(data_in_2_23_in_data), .out_data(data_in_2_23_out_data));

	reg [31:0] data_in_3_25_in_data;
	wire [31:0] data_in_3_25_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_25(.in_data(data_in_3_25_in_data), .out_data(data_in_3_25_out_data));

	reg [31:0] data_in_3_27_in_data;
	wire [31:0] data_in_3_27_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_27(.in_data(data_in_3_27_in_data), .out_data(data_in_3_27_out_data));

	reg [31:0] data_in_3_29_in_data;
	wire [31:0] data_in_3_29_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_29(.in_data(data_in_3_29_in_data), .out_data(data_in_3_29_out_data));

	reg [0:0] data_in_3_31_in_data;
	wire [0:0] data_in_3_31_out_data;
	hls_wire #(.WIDTH(1)) data_in_3_31(.in_data(data_in_3_31_in_data), .out_data(data_in_3_31_out_data));

	reg [31:0] data_in_4_33_in_data;
	wire [31:0] data_in_4_33_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_33(.in_data(data_in_4_33_in_data), .out_data(data_in_4_33_out_data));

	reg [31:0] data_in_4_35_in_data;
	wire [31:0] data_in_4_35_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_35(.in_data(data_in_4_35_in_data), .out_data(data_in_4_35_out_data));

	reg [31:0] data_in_4_37_in_data;
	wire [31:0] data_in_4_37_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_37(.in_data(data_in_4_37_in_data), .out_data(data_in_4_37_out_data));

	reg [0:0] data_in_4_39_in_data;
	wire [0:0] data_in_4_39_out_data;
	hls_wire #(.WIDTH(1)) data_in_4_39(.in_data(data_in_4_39_in_data), .out_data(data_in_4_39_out_data));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] bb_8_active_in_state_1_in_data;
	wire [0:0] bb_8_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active_in_state_1(.in_data(bb_8_active_in_state_1_in_data), .out_data(bb_8_active_in_state_1_out_data));

	reg [31:0] bb_8_predecessor_in_state_1_in_data;
	wire [31:0] bb_8_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor_in_state_1(.in_data(bb_8_predecessor_in_state_1_in_data), .out_data(bb_8_predecessor_in_state_1_out_data));

	reg [0:0] bb_9_active_in_state_1_in_data;
	wire [0:0] bb_9_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_9_active_in_state_1(.in_data(bb_9_active_in_state_1_in_data), .out_data(bb_9_active_in_state_1_out_data));

	reg [31:0] bb_9_predecessor_in_state_1_in_data;
	wire [31:0] bb_9_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_9_predecessor_in_state_1(.in_data(bb_9_predecessor_in_state_1_in_data), .out_data(bb_9_predecessor_in_state_1_out_data));

	reg [0:0] bb_0_active_in_state_1_in_data;
	wire [0:0] bb_0_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_1(.in_data(bb_0_active_in_state_1_in_data), .out_data(bb_0_active_in_state_1_out_data));

	reg [31:0] bb_0_predecessor_in_state_1_in_data;
	wire [31:0] bb_0_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_1(.in_data(bb_0_predecessor_in_state_1_in_data), .out_data(bb_0_predecessor_in_state_1_out_data));

	reg [0:0] bb_3_active_in_state_1_in_data;
	wire [0:0] bb_3_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_1(.in_data(bb_3_active_in_state_1_in_data), .out_data(bb_3_active_in_state_1_out_data));

	reg [31:0] bb_3_predecessor_in_state_1_in_data;
	wire [31:0] bb_3_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_1(.in_data(bb_3_predecessor_in_state_1_in_data), .out_data(bb_3_predecessor_in_state_1_out_data));

	reg [0:0] bb_10_active_in_state_2_in_data;
	wire [0:0] bb_10_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_2(.in_data(bb_10_active_in_state_2_in_data), .out_data(bb_10_active_in_state_2_out_data));

	reg [31:0] bb_10_predecessor_in_state_2_in_data;
	wire [31:0] bb_10_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_2(.in_data(bb_10_predecessor_in_state_2_in_data), .out_data(bb_10_predecessor_in_state_2_out_data));

	reg [0:0] bb_4_active_in_state_3_in_data;
	wire [0:0] bb_4_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_3(.in_data(bb_4_active_in_state_3_in_data), .out_data(bb_4_active_in_state_3_out_data));

	reg [31:0] bb_4_predecessor_in_state_3_in_data;
	wire [31:0] bb_4_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_3(.in_data(bb_4_predecessor_in_state_3_in_data), .out_data(bb_4_predecessor_in_state_3_out_data));

	reg [0:0] bb_10_active_in_state_3_in_data;
	wire [0:0] bb_10_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_3(.in_data(bb_10_active_in_state_3_in_data), .out_data(bb_10_active_in_state_3_out_data));

	reg [31:0] bb_10_predecessor_in_state_3_in_data;
	wire [31:0] bb_10_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_3(.in_data(bb_10_predecessor_in_state_3_in_data), .out_data(bb_10_predecessor_in_state_3_out_data));

	reg [0:0] bb_2_active_in_state_4_in_data;
	wire [0:0] bb_2_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_4(.in_data(bb_2_active_in_state_4_in_data), .out_data(bb_2_active_in_state_4_out_data));

	reg [31:0] bb_2_predecessor_in_state_4_in_data;
	wire [31:0] bb_2_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_4(.in_data(bb_2_predecessor_in_state_4_in_data), .out_data(bb_2_predecessor_in_state_4_out_data));

	reg [0:0] bb_5_active_in_state_4_in_data;
	wire [0:0] bb_5_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_5_active_in_state_4(.in_data(bb_5_active_in_state_4_in_data), .out_data(bb_5_active_in_state_4_out_data));

	reg [31:0] bb_5_predecessor_in_state_4_in_data;
	wire [31:0] bb_5_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_5_predecessor_in_state_4(.in_data(bb_5_predecessor_in_state_4_in_data), .out_data(bb_5_predecessor_in_state_4_out_data));

	reg [0:0] bb_7_active_in_state_4_in_data;
	wire [0:0] bb_7_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_7_active_in_state_4(.in_data(bb_7_active_in_state_4_in_data), .out_data(bb_7_active_in_state_4_out_data));

	reg [31:0] bb_7_predecessor_in_state_4_in_data;
	wire [31:0] bb_7_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_7_predecessor_in_state_4(.in_data(bb_7_predecessor_in_state_4_in_data), .out_data(bb_7_predecessor_in_state_4_out_data));

	reg [0:0] bb_6_active_in_state_4_in_data;
	wire [0:0] bb_6_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_6_active_in_state_4(.in_data(bb_6_active_in_state_4_in_data), .out_data(bb_6_active_in_state_4_out_data));

	reg [31:0] bb_6_predecessor_in_state_4_in_data;
	wire [31:0] bb_6_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_6_predecessor_in_state_4(.in_data(bb_6_predecessor_in_state_4_in_data), .out_data(bb_6_predecessor_in_state_4_out_data));

	reg [0:0] bb_4_active_in_state_4_in_data;
	wire [0:0] bb_4_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_4(.in_data(bb_4_active_in_state_4_in_data), .out_data(bb_4_active_in_state_4_out_data));

	reg [31:0] bb_4_predecessor_in_state_4_in_data;
	wire [31:0] bb_4_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_4(.in_data(bb_4_predecessor_in_state_4_in_data), .out_data(bb_4_predecessor_in_state_4_out_data));

	reg [0:0] bb_1_active_in_state_4_in_data;
	wire [0:0] bb_1_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_4(.in_data(bb_1_active_in_state_4_in_data), .out_data(bb_1_active_in_state_4_out_data));

	reg [31:0] bb_1_predecessor_in_state_4_in_data;
	wire [31:0] bb_1_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_4(.in_data(bb_1_predecessor_in_state_4_in_data), .out_data(bb_1_predecessor_in_state_4_out_data));

	reg [0:0] andOp_40_in0;
	reg [0:0] andOp_40_in1;
	wire [0:0] andOp_40_out;
	andOp #(.WIDTH(1)) andOp_40(.in0(andOp_40_in0), .in1(andOp_40_in1), .out(andOp_40_out));

	reg [0:0] andOp_41_in0;
	reg [0:0] andOp_41_in1;
	wire [0:0] andOp_41_out;
	andOp #(.WIDTH(1)) andOp_41(.in0(andOp_41_in0), .in1(andOp_41_in1), .out(andOp_41_out));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] notOp_42_in0;
	wire [0:0] notOp_42_out;
	notOp #(.WIDTH(1)) notOp_42(.in(notOp_42_in0), .out(notOp_42_out));

	reg [0:0] andOp_43_in0;
	reg [0:0] andOp_43_in1;
	wire [0:0] andOp_43_out;
	andOp #(.WIDTH(1)) andOp_43(.in0(andOp_43_in0), .in1(andOp_43_in1), .out(andOp_43_out));

	reg [0:0] andOp_44_in0;
	reg [0:0] andOp_44_in1;
	wire [0:0] andOp_44_out;
	andOp #(.WIDTH(1)) andOp_44(.in0(andOp_44_in0), .in1(andOp_44_in1), .out(andOp_44_out));

	reg [0:0] br_8_happened_in_state_1_in_data;
	wire [0:0] br_8_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_8_happened_in_state_1(.in_data(br_8_happened_in_state_1_in_data), .out_data(br_8_happened_in_state_1_out_data));

	reg [0:0] notOp_45_in0;
	wire [0:0] notOp_45_out;
	notOp #(.WIDTH(1)) notOp_45(.in(notOp_45_in0), .out(notOp_45_out));

	reg [0:0] andOp_46_in0;
	reg [0:0] andOp_46_in1;
	wire [0:0] andOp_46_out;
	andOp #(.WIDTH(1)) andOp_46(.in0(andOp_46_in0), .in1(andOp_46_in1), .out(andOp_46_out));

	reg [0:0] andOp_47_in0;
	reg [0:0] andOp_47_in1;
	wire [0:0] andOp_47_out;
	andOp #(.WIDTH(1)) andOp_47(.in0(andOp_47_in0), .in1(andOp_47_in1), .out(andOp_47_out));

	reg [0:0] br_9_happened_in_state_1_in_data;
	wire [0:0] br_9_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_9_happened_in_state_1(.in_data(br_9_happened_in_state_1_in_data), .out_data(br_9_happened_in_state_1_out_data));

	reg [0:0] notOp_48_in0;
	wire [0:0] notOp_48_out;
	notOp #(.WIDTH(1)) notOp_48(.in(notOp_48_in0), .out(notOp_48_out));

	reg [0:0] andOp_49_in0;
	reg [0:0] andOp_49_in1;
	wire [0:0] andOp_49_out;
	andOp #(.WIDTH(1)) andOp_49(.in0(andOp_49_in0), .in1(andOp_49_in1), .out(andOp_49_out));

	reg [0:0] notOp_50_in0;
	wire [0:0] notOp_50_out;
	notOp #(.WIDTH(1)) notOp_50(.in(notOp_50_in0), .out(notOp_50_out));

	reg [0:0] andOp_51_in0;
	reg [0:0] andOp_51_in1;
	wire [0:0] andOp_51_out;
	andOp #(.WIDTH(1)) andOp_51(.in0(andOp_51_in0), .in1(andOp_51_in1), .out(andOp_51_out));

	reg [0:0] andOp_52_in0;
	reg [0:0] andOp_52_in1;
	wire [0:0] andOp_52_out;
	andOp #(.WIDTH(1)) andOp_52(.in0(andOp_52_in0), .in1(andOp_52_in1), .out(andOp_52_out));

	reg [0:0] andOp_53_in0;
	reg [0:0] andOp_53_in1;
	wire [0:0] andOp_53_out;
	andOp #(.WIDTH(1)) andOp_53(.in0(andOp_53_in0), .in1(andOp_53_in1), .out(andOp_53_out));

	reg [0:0] br_0_happened_in_state_1_in_data;
	wire [0:0] br_0_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_1(.in_data(br_0_happened_in_state_1_in_data), .out_data(br_0_happened_in_state_1_out_data));

	reg [0:0] notOp_54_in0;
	wire [0:0] notOp_54_out;
	notOp #(.WIDTH(1)) notOp_54(.in(notOp_54_in0), .out(notOp_54_out));

	reg [0:0] andOp_55_in0;
	reg [0:0] andOp_55_in1;
	wire [0:0] andOp_55_out;
	andOp #(.WIDTH(1)) andOp_55(.in0(andOp_55_in0), .in1(andOp_55_in1), .out(andOp_55_out));

	reg [0:0] andOp_56_in0;
	reg [0:0] andOp_56_in1;
	wire [0:0] andOp_56_out;
	andOp #(.WIDTH(1)) andOp_56(.in0(andOp_56_in0), .in1(andOp_56_in1), .out(andOp_56_out));

	reg [0:0] br_3_happened_in_state_1_in_data;
	wire [0:0] br_3_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_1(.in_data(br_3_happened_in_state_1_in_data), .out_data(br_3_happened_in_state_1_out_data));

	reg [0:0] notOp_57_in0;
	wire [0:0] notOp_57_out;
	notOp #(.WIDTH(1)) notOp_57(.in(notOp_57_in0), .out(notOp_57_out));

	reg [0:0] andOp_58_in0;
	reg [0:0] andOp_58_in1;
	wire [0:0] andOp_58_out;
	andOp #(.WIDTH(1)) andOp_58(.in0(andOp_58_in0), .in1(andOp_58_in1), .out(andOp_58_out));

	reg [0:0] andOp_59_in0;
	reg [0:0] andOp_59_in1;
	wire [0:0] andOp_59_out;
	andOp #(.WIDTH(1)) andOp_59(.in0(andOp_59_in0), .in1(andOp_59_in1), .out(andOp_59_out));

	reg [0:0] br_10_happened_in_state_2_in_data;
	wire [0:0] br_10_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_2(.in_data(br_10_happened_in_state_2_in_data), .out_data(br_10_happened_in_state_2_out_data));

	reg [0:0] notOp_60_in0;
	wire [0:0] notOp_60_out;
	notOp #(.WIDTH(1)) notOp_60(.in(notOp_60_in0), .out(notOp_60_out));

	reg [0:0] andOp_61_in0;
	reg [0:0] andOp_61_in1;
	wire [0:0] andOp_61_out;
	andOp #(.WIDTH(1)) andOp_61(.in0(andOp_61_in0), .in1(andOp_61_in1), .out(andOp_61_out));

	reg [0:0] andOp_62_in0;
	reg [0:0] andOp_62_in1;
	wire [0:0] andOp_62_out;
	andOp #(.WIDTH(1)) andOp_62(.in0(andOp_62_in0), .in1(andOp_62_in1), .out(andOp_62_out));

	reg [0:0] br_4_happened_in_state_3_in_data;
	wire [0:0] br_4_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_3(.in_data(br_4_happened_in_state_3_in_data), .out_data(br_4_happened_in_state_3_out_data));

	reg [0:0] notOp_63_in0;
	wire [0:0] notOp_63_out;
	notOp #(.WIDTH(1)) notOp_63(.in(notOp_63_in0), .out(notOp_63_out));

	reg [0:0] andOp_64_in0;
	reg [0:0] andOp_64_in1;
	wire [0:0] andOp_64_out;
	andOp #(.WIDTH(1)) andOp_64(.in0(andOp_64_in0), .in1(andOp_64_in1), .out(andOp_64_out));

	reg [0:0] notOp_65_in0;
	wire [0:0] notOp_65_out;
	notOp #(.WIDTH(1)) notOp_65(.in(notOp_65_in0), .out(notOp_65_out));

	reg [0:0] andOp_66_in0;
	reg [0:0] andOp_66_in1;
	wire [0:0] andOp_66_out;
	andOp #(.WIDTH(1)) andOp_66(.in0(andOp_66_in0), .in1(andOp_66_in1), .out(andOp_66_out));

	reg [0:0] andOp_67_in0;
	reg [0:0] andOp_67_in1;
	wire [0:0] andOp_67_out;
	andOp #(.WIDTH(1)) andOp_67(.in0(andOp_67_in0), .in1(andOp_67_in1), .out(andOp_67_out));

	reg [0:0] andOp_68_in0;
	reg [0:0] andOp_68_in1;
	wire [0:0] andOp_68_out;
	andOp #(.WIDTH(1)) andOp_68(.in0(andOp_68_in0), .in1(andOp_68_in1), .out(andOp_68_out));

	reg [0:0] br_10_happened_in_state_3_in_data;
	wire [0:0] br_10_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_3(.in_data(br_10_happened_in_state_3_in_data), .out_data(br_10_happened_in_state_3_out_data));

	reg [0:0] notOp_69_in0;
	wire [0:0] notOp_69_out;
	notOp #(.WIDTH(1)) notOp_69(.in(notOp_69_in0), .out(notOp_69_out));

	reg [0:0] andOp_70_in0;
	reg [0:0] andOp_70_in1;
	wire [0:0] andOp_70_out;
	andOp #(.WIDTH(1)) andOp_70(.in0(andOp_70_in0), .in1(andOp_70_in1), .out(andOp_70_out));

	reg [0:0] andOp_71_in0;
	reg [0:0] andOp_71_in1;
	wire [0:0] andOp_71_out;
	andOp #(.WIDTH(1)) andOp_71(.in0(andOp_71_in0), .in1(andOp_71_in1), .out(andOp_71_out));

	reg [0:0] br_5_happened_in_state_4_in_data;
	wire [0:0] br_5_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_5_happened_in_state_4(.in_data(br_5_happened_in_state_4_in_data), .out_data(br_5_happened_in_state_4_out_data));

	reg [0:0] notOp_72_in0;
	wire [0:0] notOp_72_out;
	notOp #(.WIDTH(1)) notOp_72(.in(notOp_72_in0), .out(notOp_72_out));

	reg [0:0] andOp_73_in0;
	reg [0:0] andOp_73_in1;
	wire [0:0] andOp_73_out;
	andOp #(.WIDTH(1)) andOp_73(.in0(andOp_73_in0), .in1(andOp_73_in1), .out(andOp_73_out));

	reg [0:0] andOp_74_in0;
	reg [0:0] andOp_74_in1;
	wire [0:0] andOp_74_out;
	andOp #(.WIDTH(1)) andOp_74(.in0(andOp_74_in0), .in1(andOp_74_in1), .out(andOp_74_out));

	reg [0:0] br_7_happened_in_state_4_in_data;
	wire [0:0] br_7_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_7_happened_in_state_4(.in_data(br_7_happened_in_state_4_in_data), .out_data(br_7_happened_in_state_4_out_data));

	reg [0:0] notOp_75_in0;
	wire [0:0] notOp_75_out;
	notOp #(.WIDTH(1)) notOp_75(.in(notOp_75_in0), .out(notOp_75_out));

	reg [0:0] andOp_76_in0;
	reg [0:0] andOp_76_in1;
	wire [0:0] andOp_76_out;
	andOp #(.WIDTH(1)) andOp_76(.in0(andOp_76_in0), .in1(andOp_76_in1), .out(andOp_76_out));

	reg [0:0] andOp_77_in0;
	reg [0:0] andOp_77_in1;
	wire [0:0] andOp_77_out;
	andOp #(.WIDTH(1)) andOp_77(.in0(andOp_77_in0), .in1(andOp_77_in1), .out(andOp_77_out));

	reg [0:0] br_6_happened_in_state_4_in_data;
	wire [0:0] br_6_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_6_happened_in_state_4(.in_data(br_6_happened_in_state_4_in_data), .out_data(br_6_happened_in_state_4_out_data));

	reg [0:0] notOp_78_in0;
	wire [0:0] notOp_78_out;
	notOp #(.WIDTH(1)) notOp_78(.in(notOp_78_in0), .out(notOp_78_out));

	reg [0:0] andOp_79_in0;
	reg [0:0] andOp_79_in1;
	wire [0:0] andOp_79_out;
	andOp #(.WIDTH(1)) andOp_79(.in0(andOp_79_in0), .in1(andOp_79_in1), .out(andOp_79_out));

	reg [0:0] notOp_80_in0;
	wire [0:0] notOp_80_out;
	notOp #(.WIDTH(1)) notOp_80(.in(notOp_80_in0), .out(notOp_80_out));

	reg [0:0] andOp_81_in0;
	reg [0:0] andOp_81_in1;
	wire [0:0] andOp_81_out;
	andOp #(.WIDTH(1)) andOp_81(.in0(andOp_81_in0), .in1(andOp_81_in1), .out(andOp_81_out));

	reg [0:0] andOp_82_in0;
	reg [0:0] andOp_82_in1;
	wire [0:0] andOp_82_out;
	andOp #(.WIDTH(1)) andOp_82(.in0(andOp_82_in0), .in1(andOp_82_in1), .out(andOp_82_out));

	reg [0:0] andOp_83_in0;
	reg [0:0] andOp_83_in1;
	wire [0:0] andOp_83_out;
	andOp #(.WIDTH(1)) andOp_83(.in0(andOp_83_in0), .in1(andOp_83_in1), .out(andOp_83_out));

	reg [0:0] br_4_happened_in_state_4_in_data;
	wire [0:0] br_4_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_4(.in_data(br_4_happened_in_state_4_in_data), .out_data(br_4_happened_in_state_4_out_data));

	reg [0:0] notOp_84_in0;
	wire [0:0] notOp_84_out;
	notOp #(.WIDTH(1)) notOp_84(.in(notOp_84_in0), .out(notOp_84_out));

	reg [0:0] andOp_85_in0;
	reg [0:0] andOp_85_in1;
	wire [0:0] andOp_85_out;
	andOp #(.WIDTH(1)) andOp_85(.in0(andOp_85_in0), .in1(andOp_85_in1), .out(andOp_85_out));

	reg [0:0] notOp_86_in0;
	wire [0:0] notOp_86_out;
	notOp #(.WIDTH(1)) notOp_86(.in(notOp_86_in0), .out(notOp_86_out));

	reg [0:0] andOp_87_in0;
	reg [0:0] andOp_87_in1;
	wire [0:0] andOp_87_out;
	andOp #(.WIDTH(1)) andOp_87(.in0(andOp_87_in0), .in1(andOp_87_in1), .out(andOp_87_out));

	reg [0:0] andOp_88_in0;
	reg [0:0] andOp_88_in1;
	wire [0:0] andOp_88_out;
	andOp #(.WIDTH(1)) andOp_88(.in0(andOp_88_in0), .in1(andOp_88_in1), .out(andOp_88_out));

	reg [0:0] andOp_89_in0;
	reg [0:0] andOp_89_in1;
	wire [0:0] andOp_89_out;
	andOp #(.WIDTH(1)) andOp_89(.in0(andOp_89_in0), .in1(andOp_89_in1), .out(andOp_89_out));

	reg [0:0] br_1_happened_in_state_4_in_data;
	wire [0:0] br_1_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened_in_state_4(.in_data(br_1_happened_in_state_4_in_data), .out_data(br_1_happened_in_state_4_out_data));

	reg [0:0] notOp_90_in0;
	wire [0:0] notOp_90_out;
	notOp #(.WIDTH(1)) notOp_90(.in(notOp_90_in0), .out(notOp_90_out));

	reg [31:0] eq_91_in0;
	reg [31:0] eq_91_in1;
	wire [0:0] eq_91_out;
	eq #(.WIDTH(32)) eq_91(.in0(eq_91_in0), .in1(eq_91_in1), .out(eq_91_out));

	reg [31:0] eq_92_in0;
	reg [31:0] eq_92_in1;
	wire [0:0] eq_92_out;
	eq #(.WIDTH(32)) eq_92(.in0(eq_92_in0), .in1(eq_92_in1), .out(eq_92_out));

	reg [0:0] orOp_93_in0;
	reg [0:0] orOp_93_in1;
	wire [0:0] orOp_93_out;
	orOp #(.WIDTH(1)) orOp_93(.in0(orOp_93_in0), .in1(orOp_93_in1), .out(orOp_93_out));

	reg [31:0] eq_94_in0;
	reg [31:0] eq_94_in1;
	wire [0:0] eq_94_out;
	eq #(.WIDTH(32)) eq_94(.in0(eq_94_in0), .in1(eq_94_in1), .out(eq_94_out));

	reg [0:0] orOp_95_in0;
	reg [0:0] orOp_95_in1;
	wire [0:0] orOp_95_out;
	orOp #(.WIDTH(1)) orOp_95(.in0(orOp_95_in0), .in1(orOp_95_in1), .out(orOp_95_out));

	reg [31:0] eq_96_in0;
	reg [31:0] eq_96_in1;
	wire [0:0] eq_96_out;
	eq #(.WIDTH(32)) eq_96(.in0(eq_96_in0), .in1(eq_96_in1), .out(eq_96_out));

	reg [31:0] eq_97_in0;
	reg [31:0] eq_97_in1;
	wire [0:0] eq_97_out;
	eq #(.WIDTH(32)) eq_97(.in0(eq_97_in0), .in1(eq_97_in1), .out(eq_97_out));

	reg [0:0] orOp_98_in0;
	reg [0:0] orOp_98_in1;
	wire [0:0] orOp_98_out;
	orOp #(.WIDTH(1)) orOp_98(.in0(orOp_98_in0), .in1(orOp_98_in1), .out(orOp_98_out));

	reg [31:0] eq_99_in0;
	reg [31:0] eq_99_in1;
	wire [0:0] eq_99_out;
	eq #(.WIDTH(32)) eq_99(.in0(eq_99_in0), .in1(eq_99_in1), .out(eq_99_out));

	reg [31:0] eq_100_in0;
	reg [31:0] eq_100_in1;
	wire [0:0] eq_100_out;
	eq #(.WIDTH(32)) eq_100(.in0(eq_100_in0), .in1(eq_100_in1), .out(eq_100_out));

	reg [0:0] orOp_101_in0;
	reg [0:0] orOp_101_in1;
	wire [0:0] orOp_101_out;
	orOp #(.WIDTH(1)) orOp_101(.in0(orOp_101_in0), .in1(orOp_101_in1), .out(orOp_101_out));

	reg [31:0] eq_102_in0;
	reg [31:0] eq_102_in1;
	wire [0:0] eq_102_out;
	eq #(.WIDTH(32)) eq_102(.in0(eq_102_in0), .in1(eq_102_in1), .out(eq_102_out));

	reg [31:0] eq_103_in0;
	reg [31:0] eq_103_in1;
	wire [0:0] eq_103_out;
	eq #(.WIDTH(32)) eq_103(.in0(eq_103_in0), .in1(eq_103_in1), .out(eq_103_out));

	reg [0:0] orOp_104_in0;
	reg [0:0] orOp_104_in1;
	wire [0:0] orOp_104_out;
	orOp #(.WIDTH(1)) orOp_104(.in0(orOp_104_in0), .in1(orOp_104_in1), .out(orOp_104_out));

	reg [31:0] eq_105_in0;
	reg [31:0] eq_105_in1;
	wire [0:0] eq_105_out;
	eq #(.WIDTH(32)) eq_105(.in0(eq_105_in0), .in1(eq_105_in1), .out(eq_105_out));

	reg [0:0] orOp_106_in0;
	reg [0:0] orOp_106_in1;
	wire [0:0] orOp_106_out;
	orOp #(.WIDTH(1)) orOp_106(.in0(orOp_106_in0), .in1(orOp_106_in1), .out(orOp_106_out));

	reg [31:0] eq_107_in0;
	reg [31:0] eq_107_in1;
	wire [0:0] eq_107_out;
	eq #(.WIDTH(32)) eq_107(.in0(eq_107_in0), .in1(eq_107_in1), .out(eq_107_out));

	reg [0:0] orOp_108_in0;
	reg [0:0] orOp_108_in1;
	wire [0:0] orOp_108_out;
	orOp #(.WIDTH(1)) orOp_108(.in0(orOp_108_in0), .in1(orOp_108_in1), .out(orOp_108_out));

	reg [31:0] eq_109_in0;
	reg [31:0] eq_109_in1;
	wire [0:0] eq_109_out;
	eq #(.WIDTH(32)) eq_109(.in0(eq_109_in0), .in1(eq_109_in1), .out(eq_109_out));

	reg [0:0] orOp_110_in0;
	reg [0:0] orOp_110_in1;
	wire [0:0] orOp_110_out;
	orOp #(.WIDTH(1)) orOp_110(.in0(orOp_110_in0), .in1(orOp_110_in1), .out(orOp_110_out));

	reg [31:0] eq_111_in0;
	reg [31:0] eq_111_in1;
	wire [0:0] eq_111_out;
	eq #(.WIDTH(32)) eq_111(.in0(eq_111_in0), .in1(eq_111_in1), .out(eq_111_out));

	reg [31:0] eq_112_in0;
	reg [31:0] eq_112_in1;
	wire [0:0] eq_112_out;
	eq #(.WIDTH(32)) eq_112(.in0(eq_112_in0), .in1(eq_112_in1), .out(eq_112_out));

	reg [0:0] orOp_113_in0;
	reg [0:0] orOp_113_in1;
	wire [0:0] orOp_113_out;
	orOp #(.WIDTH(1)) orOp_113(.in0(orOp_113_in0), .in1(orOp_113_in1), .out(orOp_113_out));

	reg [31:0] eq_114_in0;
	reg [31:0] eq_114_in1;
	wire [0:0] eq_114_out;
	eq #(.WIDTH(32)) eq_114(.in0(eq_114_in0), .in1(eq_114_in1), .out(eq_114_out));

	reg [31:0] eq_115_in0;
	reg [31:0] eq_115_in1;
	wire [0:0] eq_115_out;
	eq #(.WIDTH(32)) eq_115(.in0(eq_115_in0), .in1(eq_115_in1), .out(eq_115_out));

	reg [0:0] notOp_116_in0;
	wire [0:0] notOp_116_out;
	notOp #(.WIDTH(1)) notOp_116(.in(notOp_116_in0), .out(notOp_116_out));

	reg [0:0] andOp_117_in0;
	reg [0:0] andOp_117_in1;
	wire [0:0] andOp_117_out;
	andOp #(.WIDTH(1)) andOp_117(.in0(andOp_117_in0), .in1(andOp_117_in1), .out(andOp_117_out));

	reg [31:0] eq_118_in0;
	reg [31:0] eq_118_in1;
	wire [0:0] eq_118_out;
	eq #(.WIDTH(32)) eq_118(.in0(eq_118_in0), .in1(eq_118_in1), .out(eq_118_out));

	reg [0:0] notOp_119_in0;
	wire [0:0] notOp_119_out;
	notOp #(.WIDTH(1)) notOp_119(.in(notOp_119_in0), .out(notOp_119_out));

	reg [0:0] andOp_120_in0;
	reg [0:0] andOp_120_in1;
	wire [0:0] andOp_120_out;
	andOp #(.WIDTH(1)) andOp_120(.in0(andOp_120_in0), .in1(andOp_120_in1), .out(andOp_120_out));

	reg [31:0] eq_121_in0;
	reg [31:0] eq_121_in1;
	wire [0:0] eq_121_out;
	eq #(.WIDTH(32)) eq_121(.in0(eq_121_in0), .in1(eq_121_in1), .out(eq_121_out));

	reg [31:0] eq_122_in0;
	reg [31:0] eq_122_in1;
	wire [0:0] eq_122_out;
	eq #(.WIDTH(32)) eq_122(.in0(eq_122_in0), .in1(eq_122_in1), .out(eq_122_out));

	reg [0:0] notOp_123_in0;
	wire [0:0] notOp_123_out;
	notOp #(.WIDTH(1)) notOp_123(.in(notOp_123_in0), .out(notOp_123_out));

	reg [0:0] andOp_124_in0;
	reg [0:0] andOp_124_in1;
	wire [0:0] andOp_124_out;
	andOp #(.WIDTH(1)) andOp_124(.in0(andOp_124_in0), .in1(andOp_124_in1), .out(andOp_124_out));

	reg [31:0] eq_125_in0;
	reg [31:0] eq_125_in1;
	wire [0:0] eq_125_out;
	eq #(.WIDTH(32)) eq_125(.in0(eq_125_in0), .in1(eq_125_in1), .out(eq_125_out));

	reg [31:0] eq_126_in0;
	reg [31:0] eq_126_in1;
	wire [0:0] eq_126_out;
	eq #(.WIDTH(32)) eq_126(.in0(eq_126_in0), .in1(eq_126_in1), .out(eq_126_out));

	reg [0:0] notOp_127_in0;
	wire [0:0] notOp_127_out;
	notOp #(.WIDTH(1)) notOp_127(.in(notOp_127_in0), .out(notOp_127_out));

	reg [0:0] andOp_128_in0;
	reg [0:0] andOp_128_in1;
	wire [0:0] andOp_128_out;
	andOp #(.WIDTH(1)) andOp_128(.in0(andOp_128_in0), .in1(andOp_128_in1), .out(andOp_128_out));

	reg [31:0] eq_129_in0;
	reg [31:0] eq_129_in1;
	wire [0:0] eq_129_out;
	eq #(.WIDTH(32)) eq_129(.in0(eq_129_in0), .in1(eq_129_in1), .out(eq_129_out));

	reg [31:0] eq_130_in0;
	reg [31:0] eq_130_in1;
	wire [0:0] eq_130_out;
	eq #(.WIDTH(32)) eq_130(.in0(eq_130_in0), .in1(eq_130_in1), .out(eq_130_out));

	reg [0:0] notOp_131_in0;
	wire [0:0] notOp_131_out;
	notOp #(.WIDTH(1)) notOp_131(.in(notOp_131_in0), .out(notOp_131_out));

	reg [0:0] andOp_132_in0;
	reg [0:0] andOp_132_in1;
	wire [0:0] andOp_132_out;
	andOp #(.WIDTH(1)) andOp_132(.in0(andOp_132_in0), .in1(andOp_132_in1), .out(andOp_132_out));

	reg [31:0] eq_133_in0;
	reg [31:0] eq_133_in1;
	wire [0:0] eq_133_out;
	eq #(.WIDTH(32)) eq_133(.in0(eq_133_in0), .in1(eq_133_in1), .out(eq_133_out));

	reg [0:0] notOp_134_in0;
	wire [0:0] notOp_134_out;
	notOp #(.WIDTH(1)) notOp_134(.in(notOp_134_in0), .out(notOp_134_out));

	reg [0:0] andOp_135_in0;
	reg [0:0] andOp_135_in1;
	wire [0:0] andOp_135_out;
	andOp #(.WIDTH(1)) andOp_135(.in0(andOp_135_in0), .in1(andOp_135_in1), .out(andOp_135_out));

	reg [31:0] eq_136_in0;
	reg [31:0] eq_136_in1;
	wire [0:0] eq_136_out;
	eq #(.WIDTH(32)) eq_136(.in0(eq_136_in0), .in1(eq_136_in1), .out(eq_136_out));

	reg [0:0] notOp_137_in0;
	wire [0:0] notOp_137_out;
	notOp #(.WIDTH(1)) notOp_137(.in(notOp_137_in0), .out(notOp_137_out));

	reg [0:0] andOp_138_in0;
	reg [0:0] andOp_138_in1;
	wire [0:0] andOp_138_out;
	andOp #(.WIDTH(1)) andOp_138(.in0(andOp_138_in0), .in1(andOp_138_in1), .out(andOp_138_out));

	reg [31:0] eq_139_in0;
	reg [31:0] eq_139_in1;
	wire [0:0] eq_139_out;
	eq #(.WIDTH(32)) eq_139(.in0(eq_139_in0), .in1(eq_139_in1), .out(eq_139_out));

	reg [0:0] notOp_140_in0;
	wire [0:0] notOp_140_out;
	notOp #(.WIDTH(1)) notOp_140(.in(notOp_140_in0), .out(notOp_140_out));

	reg [0:0] andOp_141_in0;
	reg [0:0] andOp_141_in1;
	wire [0:0] andOp_141_out;
	andOp #(.WIDTH(1)) andOp_141(.in0(andOp_141_in0), .in1(andOp_141_in1), .out(andOp_141_out));

	reg [31:0] eq_142_in0;
	reg [31:0] eq_142_in1;
	wire [0:0] eq_142_out;
	eq #(.WIDTH(32)) eq_142(.in0(eq_142_in0), .in1(eq_142_in1), .out(eq_142_out));

	reg [31:0] eq_143_in0;
	reg [31:0] eq_143_in1;
	wire [0:0] eq_143_out;
	eq #(.WIDTH(32)) eq_143(.in0(eq_143_in0), .in1(eq_143_in1), .out(eq_143_out));

	reg [0:0] notOp_144_in0;
	wire [0:0] notOp_144_out;
	notOp #(.WIDTH(1)) notOp_144(.in(notOp_144_in0), .out(notOp_144_out));

	reg [0:0] andOp_145_in0;
	reg [0:0] andOp_145_in1;
	wire [0:0] andOp_145_out;
	andOp #(.WIDTH(1)) andOp_145(.in0(andOp_145_in0), .in1(andOp_145_in1), .out(andOp_145_out));

	reg [0:0] andOp_146_in0;
	reg [0:0] andOp_146_in1;
	wire [0:0] andOp_146_out;
	andOp #(.WIDTH(1)) andOp_146(.in0(andOp_146_in0), .in1(andOp_146_in1), .out(andOp_146_out));

	reg [0:0] andOp_147_in0;
	reg [0:0] andOp_147_in1;
	wire [0:0] andOp_147_out;
	andOp #(.WIDTH(1)) andOp_147(.in0(andOp_147_in0), .in1(andOp_147_in1), .out(andOp_147_out));

	reg [0:0] andOp_148_in0;
	reg [0:0] andOp_148_in1;
	wire [0:0] andOp_148_out;
	andOp #(.WIDTH(1)) andOp_148(.in0(andOp_148_in0), .in1(andOp_148_in1), .out(andOp_148_out));

	reg [0:0] andOp_149_in0;
	reg [0:0] andOp_149_in1;
	wire [0:0] andOp_149_out;
	andOp #(.WIDTH(1)) andOp_149(.in0(andOp_149_in0), .in1(andOp_149_in1), .out(andOp_149_out));

	reg [0:0] andOp_150_in0;
	reg [0:0] andOp_150_in1;
	wire [0:0] andOp_150_out;
	andOp #(.WIDTH(1)) andOp_150(.in0(andOp_150_in0), .in1(andOp_150_in1), .out(andOp_150_out));

	reg [0:0] andOp_151_in0;
	reg [0:0] andOp_151_in1;
	wire [0:0] andOp_151_out;
	andOp #(.WIDTH(1)) andOp_151(.in0(andOp_151_in0), .in1(andOp_151_in1), .out(andOp_151_out));

	reg [0:0] andOp_152_in0;
	reg [0:0] andOp_152_in1;
	wire [0:0] andOp_152_out;
	andOp #(.WIDTH(1)) andOp_152(.in0(andOp_152_in0), .in1(andOp_152_in1), .out(andOp_152_out));

	reg [0:0] andOp_153_in0;
	reg [0:0] andOp_153_in1;
	wire [0:0] andOp_153_out;
	andOp #(.WIDTH(1)) andOp_153(.in0(andOp_153_in0), .in1(andOp_153_in1), .out(andOp_153_out));

	reg [0:0] andOp_154_in0;
	reg [0:0] andOp_154_in1;
	wire [0:0] andOp_154_out;
	andOp #(.WIDTH(1)) andOp_154(.in0(andOp_154_in0), .in1(andOp_154_in1), .out(andOp_154_out));

	reg [0:0] andOp_155_in0;
	reg [0:0] andOp_155_in1;
	wire [0:0] andOp_155_out;
	andOp #(.WIDTH(1)) andOp_155(.in0(andOp_155_in0), .in1(andOp_155_in1), .out(andOp_155_out));

	reg [0:0] andOp_156_in0;
	reg [0:0] andOp_156_in1;
	wire [0:0] andOp_156_out;
	andOp #(.WIDTH(1)) andOp_156(.in0(andOp_156_in0), .in1(andOp_156_in1), .out(andOp_156_out));

	reg [31:0] concat_157_in0;
	reg [31:0] concat_157_in1;
	wire [63:0] concat_157_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_157(.in0(concat_157_in0), .in1(concat_157_in1), .out(concat_157_out));

	reg [31:0] concat_158_in0;
	reg [31:0] concat_158_in1;
	wire [63:0] concat_158_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_158(.in0(concat_158_in0), .in1(concat_158_in1), .out(concat_158_out));

	reg [0:0] andOp_159_in0;
	reg [0:0] andOp_159_in1;
	wire [0:0] andOp_159_out;
	andOp #(.WIDTH(1)) andOp_159(.in0(andOp_159_in0), .in1(andOp_159_in1), .out(andOp_159_out));

	reg [31:0] tmp_output_160_in_data;
	wire [31:0] tmp_output_160_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_160(.in_data(tmp_output_160_in_data), .out_data(tmp_output_160_out_data));

	reg [31:0] eq_161_in0;
	reg [31:0] eq_161_in1;
	wire [0:0] eq_161_out;
	eq #(.WIDTH(32)) eq_161(.in0(eq_161_in0), .in1(eq_161_in1), .out(eq_161_out));

	reg [0:0] andOp_162_in0;
	reg [0:0] andOp_162_in1;
	wire [0:0] andOp_162_out;
	andOp #(.WIDTH(1)) andOp_162(.in0(andOp_162_in0), .in1(andOp_162_in1), .out(andOp_162_out));

	reg [0:0] andOp_163_in0;
	reg [0:0] andOp_163_in1;
	wire [0:0] andOp_163_out;
	andOp #(.WIDTH(1)) andOp_163(.in0(andOp_163_in0), .in1(andOp_163_in1), .out(andOp_163_out));

	reg [0:0] andOp_164_in0;
	reg [0:0] andOp_164_in1;
	wire [0:0] andOp_164_out;
	andOp #(.WIDTH(1)) andOp_164(.in0(andOp_164_in0), .in1(andOp_164_in1), .out(andOp_164_out));

	reg [0:0] andOp_165_in0;
	reg [0:0] andOp_165_in1;
	wire [0:0] andOp_165_out;
	andOp #(.WIDTH(1)) andOp_165(.in0(andOp_165_in0), .in1(andOp_165_in1), .out(andOp_165_out));

	reg [0:0] andOp_166_in0;
	reg [0:0] andOp_166_in1;
	wire [0:0] andOp_166_out;
	andOp #(.WIDTH(1)) andOp_166(.in0(andOp_166_in0), .in1(andOp_166_in1), .out(andOp_166_out));

	reg [0:0] andOp_167_in0;
	reg [0:0] andOp_167_in1;
	wire [0:0] andOp_167_out;
	andOp #(.WIDTH(1)) andOp_167(.in0(andOp_167_in0), .in1(andOp_167_in1), .out(andOp_167_out));

	reg [0:0] andOp_168_in0;
	reg [0:0] andOp_168_in1;
	wire [0:0] andOp_168_out;
	andOp #(.WIDTH(1)) andOp_168(.in0(andOp_168_in0), .in1(andOp_168_in1), .out(andOp_168_out));

	reg [0:0] andOp_169_in0;
	reg [0:0] andOp_169_in1;
	wire [0:0] andOp_169_out;
	andOp #(.WIDTH(1)) andOp_169(.in0(andOp_169_in0), .in1(andOp_169_in1), .out(andOp_169_out));

	reg [0:0] andOp_170_in0;
	reg [0:0] andOp_170_in1;
	wire [0:0] andOp_170_out;
	andOp #(.WIDTH(1)) andOp_170(.in0(andOp_170_in0), .in1(andOp_170_in1), .out(andOp_170_out));

	reg [0:0] andOp_171_in0;
	reg [0:0] andOp_171_in1;
	wire [0:0] andOp_171_out;
	andOp #(.WIDTH(1)) andOp_171(.in0(andOp_171_in0), .in1(andOp_171_in1), .out(andOp_171_out));

	reg [0:0] andOp_172_in0;
	reg [0:0] andOp_172_in1;
	wire [0:0] andOp_172_out;
	andOp #(.WIDTH(1)) andOp_172(.in0(andOp_172_in0), .in1(andOp_172_in1), .out(andOp_172_out));

	reg [0:0] notOp_173_in0;
	wire [0:0] notOp_173_out;
	notOp #(.WIDTH(1)) notOp_173(.in(notOp_173_in0), .out(notOp_173_out));

	reg [0:0] andOp_174_in0;
	reg [0:0] andOp_174_in1;
	wire [0:0] andOp_174_out;
	andOp #(.WIDTH(1)) andOp_174(.in0(andOp_174_in0), .in1(andOp_174_in1), .out(andOp_174_out));

	reg [0:0] notOp_175_in0;
	wire [0:0] notOp_175_out;
	notOp #(.WIDTH(1)) notOp_175(.in(notOp_175_in0), .out(notOp_175_out));

	reg [0:0] andOp_176_in0;
	reg [0:0] andOp_176_in1;
	wire [0:0] andOp_176_out;
	andOp #(.WIDTH(1)) andOp_176(.in0(andOp_176_in0), .in1(andOp_176_in1), .out(andOp_176_out));

	reg [0:0] notOp_177_in0;
	wire [0:0] notOp_177_out;
	notOp #(.WIDTH(1)) notOp_177(.in(notOp_177_in0), .out(notOp_177_out));

	reg [0:0] andOp_178_in0;
	reg [0:0] andOp_178_in1;
	wire [0:0] andOp_178_out;
	andOp #(.WIDTH(1)) andOp_178(.in0(andOp_178_in0), .in1(andOp_178_in1), .out(andOp_178_out));

	reg [0:0] notOp_179_in0;
	wire [0:0] notOp_179_out;
	notOp #(.WIDTH(1)) notOp_179(.in(notOp_179_in0), .out(notOp_179_out));

	reg [0:0] andOp_180_in0;
	reg [0:0] andOp_180_in1;
	wire [0:0] andOp_180_out;
	andOp #(.WIDTH(1)) andOp_180(.in0(andOp_180_in0), .in1(andOp_180_in1), .out(andOp_180_out));

	reg [0:0] notOp_181_in0;
	wire [0:0] notOp_181_out;
	notOp #(.WIDTH(1)) notOp_181(.in(notOp_181_in0), .out(notOp_181_out));

	reg [0:0] andOp_182_in0;
	reg [0:0] andOp_182_in1;
	wire [0:0] andOp_182_out;
	andOp #(.WIDTH(1)) andOp_182(.in0(andOp_182_in0), .in1(andOp_182_in1), .out(andOp_182_out));

	reg [0:0] notOp_183_in0;
	wire [0:0] notOp_183_out;
	notOp #(.WIDTH(1)) notOp_183(.in(notOp_183_in0), .out(notOp_183_out));

	reg [0:0] andOp_184_in0;
	reg [0:0] andOp_184_in1;
	wire [0:0] andOp_184_out;
	andOp #(.WIDTH(1)) andOp_184(.in0(andOp_184_in0), .in1(andOp_184_in1), .out(andOp_184_out));

	reg [0:0] notOp_185_in0;
	wire [0:0] notOp_185_out;
	notOp #(.WIDTH(1)) notOp_185(.in(notOp_185_in0), .out(notOp_185_out));

	reg [0:0] andOp_186_in0;
	reg [0:0] andOp_186_in1;
	wire [0:0] andOp_186_out;
	andOp #(.WIDTH(1)) andOp_186(.in0(andOp_186_in0), .in1(andOp_186_in1), .out(andOp_186_out));

	reg [0:0] notOp_187_in0;
	wire [0:0] notOp_187_out;
	notOp #(.WIDTH(1)) notOp_187(.in(notOp_187_in0), .out(notOp_187_out));

	reg [0:0] andOp_188_in0;
	reg [0:0] andOp_188_in1;
	wire [0:0] andOp_188_out;
	andOp #(.WIDTH(1)) andOp_188(.in0(andOp_188_in0), .in1(andOp_188_in1), .out(andOp_188_out));

	reg [31:0] eq_189_in0;
	reg [31:0] eq_189_in1;
	wire [0:0] eq_189_out;
	eq #(.WIDTH(32)) eq_189(.in0(eq_189_in0), .in1(eq_189_in1), .out(eq_189_out));

	reg [0:0] andOp_190_in0;
	reg [0:0] andOp_190_in1;
	wire [0:0] andOp_190_out;
	andOp #(.WIDTH(1)) andOp_190(.in0(andOp_190_in0), .in1(andOp_190_in1), .out(andOp_190_out));

	reg [31:0] eq_191_in0;
	reg [31:0] eq_191_in1;
	wire [0:0] eq_191_out;
	eq #(.WIDTH(32)) eq_191(.in0(eq_191_in0), .in1(eq_191_in1), .out(eq_191_out));

	reg [0:0] andOp_192_in0;
	reg [0:0] andOp_192_in1;
	wire [0:0] andOp_192_out;
	andOp #(.WIDTH(1)) andOp_192(.in0(andOp_192_in0), .in1(andOp_192_in1), .out(andOp_192_out));

	reg [0:0] notOp_193_in0;
	wire [0:0] notOp_193_out;
	notOp #(.WIDTH(1)) notOp_193(.in(notOp_193_in0), .out(notOp_193_out));

	reg [0:0] andOp_194_in0;
	reg [0:0] andOp_194_in1;
	wire [0:0] andOp_194_out;
	andOp #(.WIDTH(1)) andOp_194(.in0(andOp_194_in0), .in1(andOp_194_in1), .out(andOp_194_out));

	reg [0:0] notOp_195_in0;
	wire [0:0] notOp_195_out;
	notOp #(.WIDTH(1)) notOp_195(.in(notOp_195_in0), .out(notOp_195_out));

	reg [0:0] andOp_196_in0;
	reg [0:0] andOp_196_in1;
	wire [0:0] andOp_196_out;
	andOp #(.WIDTH(1)) andOp_196(.in0(andOp_196_in0), .in1(andOp_196_in1), .out(andOp_196_out));

	reg [0:0] notOp_197_in0;
	wire [0:0] notOp_197_out;
	notOp #(.WIDTH(1)) notOp_197(.in(notOp_197_in0), .out(notOp_197_out));

	reg [0:0] andOp_198_in0;
	reg [0:0] andOp_198_in1;
	wire [0:0] andOp_198_out;
	andOp #(.WIDTH(1)) andOp_198(.in0(andOp_198_in0), .in1(andOp_198_in1), .out(andOp_198_out));

	reg [0:0] andOp_199_in0;
	reg [0:0] andOp_199_in1;
	wire [0:0] andOp_199_out;
	andOp #(.WIDTH(1)) andOp_199(.in0(andOp_199_in0), .in1(andOp_199_in1), .out(andOp_199_out));

	reg [31:0] eq_200_in0;
	reg [31:0] eq_200_in1;
	wire [0:0] eq_200_out;
	eq #(.WIDTH(32)) eq_200(.in0(eq_200_in0), .in1(eq_200_in1), .out(eq_200_out));

	reg [0:0] andOp_201_in0;
	reg [0:0] andOp_201_in1;
	wire [0:0] andOp_201_out;
	andOp #(.WIDTH(1)) andOp_201(.in0(andOp_201_in0), .in1(andOp_201_in1), .out(andOp_201_out));

	reg [0:0] notOp_202_in0;
	wire [0:0] notOp_202_out;
	notOp #(.WIDTH(1)) notOp_202(.in(notOp_202_in0), .out(notOp_202_out));

	reg [0:0] andOp_203_in0;
	reg [0:0] andOp_203_in1;
	wire [0:0] andOp_203_out;
	andOp #(.WIDTH(1)) andOp_203(.in0(andOp_203_in0), .in1(andOp_203_in1), .out(andOp_203_out));

	reg [0:0] notOp_204_in0;
	wire [0:0] notOp_204_out;
	notOp #(.WIDTH(1)) notOp_204(.in(notOp_204_in0), .out(notOp_204_out));

	reg [0:0] andOp_205_in0;
	reg [0:0] andOp_205_in1;
	wire [0:0] andOp_205_out;
	andOp #(.WIDTH(1)) andOp_205(.in0(andOp_205_in0), .in1(andOp_205_in1), .out(andOp_205_out));

	reg [0:0] notOp_206_in0;
	wire [0:0] notOp_206_out;
	notOp #(.WIDTH(1)) notOp_206(.in(notOp_206_in0), .out(notOp_206_out));

	reg [0:0] andOp_207_in0;
	reg [0:0] andOp_207_in1;
	wire [0:0] andOp_207_out;
	andOp #(.WIDTH(1)) andOp_207(.in0(andOp_207_in0), .in1(andOp_207_in1), .out(andOp_207_out));

	reg [0:0] andOp_208_in0;
	reg [0:0] andOp_208_in1;
	wire [0:0] andOp_208_out;
	andOp #(.WIDTH(1)) andOp_208(.in0(andOp_208_in0), .in1(andOp_208_in1), .out(andOp_208_out));

	reg [31:0] eq_209_in0;
	reg [31:0] eq_209_in1;
	wire [0:0] eq_209_out;
	eq #(.WIDTH(32)) eq_209(.in0(eq_209_in0), .in1(eq_209_in1), .out(eq_209_out));

	reg [0:0] andOp_210_in0;
	reg [0:0] andOp_210_in1;
	wire [0:0] andOp_210_out;
	andOp #(.WIDTH(1)) andOp_210(.in0(andOp_210_in0), .in1(andOp_210_in1), .out(andOp_210_out));

	reg [0:0] notOp_211_in0;
	wire [0:0] notOp_211_out;
	notOp #(.WIDTH(1)) notOp_211(.in(notOp_211_in0), .out(notOp_211_out));

	reg [0:0] andOp_212_in0;
	reg [0:0] andOp_212_in1;
	wire [0:0] andOp_212_out;
	andOp #(.WIDTH(1)) andOp_212(.in0(andOp_212_in0), .in1(andOp_212_in1), .out(andOp_212_out));

	reg [0:0] notOp_213_in0;
	wire [0:0] notOp_213_out;
	notOp #(.WIDTH(1)) notOp_213(.in(notOp_213_in0), .out(notOp_213_out));

	reg [0:0] andOp_214_in0;
	reg [0:0] andOp_214_in1;
	wire [0:0] andOp_214_out;
	andOp #(.WIDTH(1)) andOp_214(.in0(andOp_214_in0), .in1(andOp_214_in1), .out(andOp_214_out));

	reg [0:0] notOp_215_in0;
	wire [0:0] notOp_215_out;
	notOp #(.WIDTH(1)) notOp_215(.in(notOp_215_in0), .out(notOp_215_out));

	reg [0:0] andOp_216_in0;
	reg [0:0] andOp_216_in1;
	wire [0:0] andOp_216_out;
	andOp #(.WIDTH(1)) andOp_216(.in0(andOp_216_in0), .in1(andOp_216_in1), .out(andOp_216_out));

	reg [0:0] andOp_217_in0;
	reg [0:0] andOp_217_in1;
	wire [0:0] andOp_217_out;
	andOp #(.WIDTH(1)) andOp_217(.in0(andOp_217_in0), .in1(andOp_217_in1), .out(andOp_217_out));

	reg [31:0] eq_218_in0;
	reg [31:0] eq_218_in1;
	wire [0:0] eq_218_out;
	eq #(.WIDTH(32)) eq_218(.in0(eq_218_in0), .in1(eq_218_in1), .out(eq_218_out));

	reg [0:0] andOp_219_in0;
	reg [0:0] andOp_219_in1;
	wire [0:0] andOp_219_out;
	andOp #(.WIDTH(1)) andOp_219(.in0(andOp_219_in0), .in1(andOp_219_in1), .out(andOp_219_out));

	reg [0:0] notOp_220_in0;
	wire [0:0] notOp_220_out;
	notOp #(.WIDTH(1)) notOp_220(.in(notOp_220_in0), .out(notOp_220_out));

	reg [0:0] andOp_221_in0;
	reg [0:0] andOp_221_in1;
	wire [0:0] andOp_221_out;
	andOp #(.WIDTH(1)) andOp_221(.in0(andOp_221_in0), .in1(andOp_221_in1), .out(andOp_221_out));

	reg [0:0] notOp_222_in0;
	wire [0:0] notOp_222_out;
	notOp #(.WIDTH(1)) notOp_222(.in(notOp_222_in0), .out(notOp_222_out));

	reg [0:0] andOp_223_in0;
	reg [0:0] andOp_223_in1;
	wire [0:0] andOp_223_out;
	andOp #(.WIDTH(1)) andOp_223(.in0(andOp_223_in0), .in1(andOp_223_in1), .out(andOp_223_out));

	reg [0:0] notOp_224_in0;
	wire [0:0] notOp_224_out;
	notOp #(.WIDTH(1)) notOp_224(.in(notOp_224_in0), .out(notOp_224_out));

	reg [0:0] andOp_225_in0;
	reg [0:0] andOp_225_in1;
	wire [0:0] andOp_225_out;
	andOp #(.WIDTH(1)) andOp_225(.in0(andOp_225_in0), .in1(andOp_225_in1), .out(andOp_225_out));

	reg [31:0] eq_226_in0;
	reg [31:0] eq_226_in1;
	wire [0:0] eq_226_out;
	eq #(.WIDTH(32)) eq_226(.in0(eq_226_in0), .in1(eq_226_in1), .out(eq_226_out));

	reg [31:0] eq_227_in0;
	reg [31:0] eq_227_in1;
	wire [0:0] eq_227_out;
	eq #(.WIDTH(32)) eq_227(.in0(eq_227_in0), .in1(eq_227_in1), .out(eq_227_out));

	reg [31:0] eq_228_in0;
	reg [31:0] eq_228_in1;
	wire [0:0] eq_228_out;
	eq #(.WIDTH(32)) eq_228(.in0(eq_228_in0), .in1(eq_228_in1), .out(eq_228_out));

	reg [0:0] andOp_229_in0;
	reg [0:0] andOp_229_in1;
	wire [0:0] andOp_229_out;
	andOp #(.WIDTH(1)) andOp_229(.in0(andOp_229_in0), .in1(andOp_229_in1), .out(andOp_229_out));

	reg [31:0] eq_230_in0;
	reg [31:0] eq_230_in1;
	wire [0:0] eq_230_out;
	eq #(.WIDTH(32)) eq_230(.in0(eq_230_in0), .in1(eq_230_in1), .out(eq_230_out));

	reg [0:0] andOp_231_in0;
	reg [0:0] andOp_231_in1;
	wire [0:0] andOp_231_out;
	andOp #(.WIDTH(1)) andOp_231(.in0(andOp_231_in0), .in1(andOp_231_in1), .out(andOp_231_out));

	reg [0:0] notOp_232_in0;
	wire [0:0] notOp_232_out;
	notOp #(.WIDTH(1)) notOp_232(.in(notOp_232_in0), .out(notOp_232_out));

	reg [0:0] andOp_233_in0;
	reg [0:0] andOp_233_in1;
	wire [0:0] andOp_233_out;
	andOp #(.WIDTH(1)) andOp_233(.in0(andOp_233_in0), .in1(andOp_233_in1), .out(andOp_233_out));

	reg [0:0] notOp_234_in0;
	wire [0:0] notOp_234_out;
	notOp #(.WIDTH(1)) notOp_234(.in(notOp_234_in0), .out(notOp_234_out));

	reg [0:0] andOp_235_in0;
	reg [0:0] andOp_235_in1;
	wire [0:0] andOp_235_out;
	andOp #(.WIDTH(1)) andOp_235(.in0(andOp_235_in0), .in1(andOp_235_in1), .out(andOp_235_out));

	reg [0:0] notOp_236_in0;
	wire [0:0] notOp_236_out;
	notOp #(.WIDTH(1)) notOp_236(.in(notOp_236_in0), .out(notOp_236_out));

	reg [0:0] andOp_237_in0;
	reg [0:0] andOp_237_in1;
	wire [0:0] andOp_237_out;
	andOp #(.WIDTH(1)) andOp_237(.in0(andOp_237_in0), .in1(andOp_237_in1), .out(andOp_237_out));

	reg [0:0] andOp_238_in0;
	reg [0:0] andOp_238_in1;
	wire [0:0] andOp_238_out;
	andOp #(.WIDTH(1)) andOp_238(.in0(andOp_238_in0), .in1(andOp_238_in1), .out(andOp_238_out));

	reg [31:0] eq_239_in0;
	reg [31:0] eq_239_in1;
	wire [0:0] eq_239_out;
	eq #(.WIDTH(32)) eq_239(.in0(eq_239_in0), .in1(eq_239_in1), .out(eq_239_out));

	reg [0:0] andOp_240_in0;
	reg [0:0] andOp_240_in1;
	wire [0:0] andOp_240_out;
	andOp #(.WIDTH(1)) andOp_240(.in0(andOp_240_in0), .in1(andOp_240_in1), .out(andOp_240_out));

	reg [0:0] notOp_241_in0;
	wire [0:0] notOp_241_out;
	notOp #(.WIDTH(1)) notOp_241(.in(notOp_241_in0), .out(notOp_241_out));

	reg [0:0] andOp_242_in0;
	reg [0:0] andOp_242_in1;
	wire [0:0] andOp_242_out;
	andOp #(.WIDTH(1)) andOp_242(.in0(andOp_242_in0), .in1(andOp_242_in1), .out(andOp_242_out));

	reg [0:0] notOp_243_in0;
	wire [0:0] notOp_243_out;
	notOp #(.WIDTH(1)) notOp_243(.in(notOp_243_in0), .out(notOp_243_out));

	reg [0:0] andOp_244_in0;
	reg [0:0] andOp_244_in1;
	wire [0:0] andOp_244_out;
	andOp #(.WIDTH(1)) andOp_244(.in0(andOp_244_in0), .in1(andOp_244_in1), .out(andOp_244_out));

	reg [0:0] notOp_245_in0;
	wire [0:0] notOp_245_out;
	notOp #(.WIDTH(1)) notOp_245(.in(notOp_245_in0), .out(notOp_245_out));

	reg [0:0] andOp_246_in0;
	reg [0:0] andOp_246_in1;
	wire [0:0] andOp_246_out;
	andOp #(.WIDTH(1)) andOp_246(.in0(andOp_246_in0), .in1(andOp_246_in1), .out(andOp_246_out));

	reg [0:0] andOp_247_in0;
	reg [0:0] andOp_247_in1;
	wire [0:0] andOp_247_out;
	andOp #(.WIDTH(1)) andOp_247(.in0(andOp_247_in0), .in1(andOp_247_in1), .out(andOp_247_out));

	reg [31:0] eq_248_in0;
	reg [31:0] eq_248_in1;
	wire [0:0] eq_248_out;
	eq #(.WIDTH(32)) eq_248(.in0(eq_248_in0), .in1(eq_248_in1), .out(eq_248_out));

	reg [0:0] andOp_249_in0;
	reg [0:0] andOp_249_in1;
	wire [0:0] andOp_249_out;
	andOp #(.WIDTH(1)) andOp_249(.in0(andOp_249_in0), .in1(andOp_249_in1), .out(andOp_249_out));

	reg [0:0] notOp_250_in0;
	wire [0:0] notOp_250_out;
	notOp #(.WIDTH(1)) notOp_250(.in(notOp_250_in0), .out(notOp_250_out));

	reg [0:0] andOp_251_in0;
	reg [0:0] andOp_251_in1;
	wire [0:0] andOp_251_out;
	andOp #(.WIDTH(1)) andOp_251(.in0(andOp_251_in0), .in1(andOp_251_in1), .out(andOp_251_out));

	reg [0:0] notOp_252_in0;
	wire [0:0] notOp_252_out;
	notOp #(.WIDTH(1)) notOp_252(.in(notOp_252_in0), .out(notOp_252_out));

	reg [0:0] andOp_253_in0;
	reg [0:0] andOp_253_in1;
	wire [0:0] andOp_253_out;
	andOp #(.WIDTH(1)) andOp_253(.in0(andOp_253_in0), .in1(andOp_253_in1), .out(andOp_253_out));

	reg [0:0] notOp_254_in0;
	wire [0:0] notOp_254_out;
	notOp #(.WIDTH(1)) notOp_254(.in(notOp_254_in0), .out(notOp_254_out));

	reg [0:0] andOp_255_in0;
	reg [0:0] andOp_255_in1;
	wire [0:0] andOp_255_out;
	andOp #(.WIDTH(1)) andOp_255(.in0(andOp_255_in0), .in1(andOp_255_in1), .out(andOp_255_out));

	reg [0:0] andOp_256_in0;
	reg [0:0] andOp_256_in1;
	wire [0:0] andOp_256_out;
	andOp #(.WIDTH(1)) andOp_256(.in0(andOp_256_in0), .in1(andOp_256_in1), .out(andOp_256_out));

	reg [31:0] eq_257_in0;
	reg [31:0] eq_257_in1;
	wire [0:0] eq_257_out;
	eq #(.WIDTH(32)) eq_257(.in0(eq_257_in0), .in1(eq_257_in1), .out(eq_257_out));

	reg [0:0] andOp_258_in0;
	reg [0:0] andOp_258_in1;
	wire [0:0] andOp_258_out;
	andOp #(.WIDTH(1)) andOp_258(.in0(andOp_258_in0), .in1(andOp_258_in1), .out(andOp_258_out));

	reg [0:0] notOp_259_in0;
	wire [0:0] notOp_259_out;
	notOp #(.WIDTH(1)) notOp_259(.in(notOp_259_in0), .out(notOp_259_out));

	reg [0:0] andOp_260_in0;
	reg [0:0] andOp_260_in1;
	wire [0:0] andOp_260_out;
	andOp #(.WIDTH(1)) andOp_260(.in0(andOp_260_in0), .in1(andOp_260_in1), .out(andOp_260_out));

	reg [0:0] notOp_261_in0;
	wire [0:0] notOp_261_out;
	notOp #(.WIDTH(1)) notOp_261(.in(notOp_261_in0), .out(notOp_261_out));

	reg [0:0] andOp_262_in0;
	reg [0:0] andOp_262_in1;
	wire [0:0] andOp_262_out;
	andOp #(.WIDTH(1)) andOp_262(.in0(andOp_262_in0), .in1(andOp_262_in1), .out(andOp_262_out));

	reg [0:0] notOp_263_in0;
	wire [0:0] notOp_263_out;
	notOp #(.WIDTH(1)) notOp_263(.in(notOp_263_in0), .out(notOp_263_out));

	reg [0:0] andOp_264_in0;
	reg [0:0] andOp_264_in1;
	wire [0:0] andOp_264_out;
	andOp #(.WIDTH(1)) andOp_264(.in0(andOp_264_in0), .in1(andOp_264_in1), .out(andOp_264_out));

	reg [31:0] eq_265_in0;
	reg [31:0] eq_265_in1;
	wire [0:0] eq_265_out;
	eq #(.WIDTH(32)) eq_265(.in0(eq_265_in0), .in1(eq_265_in1), .out(eq_265_out));

	reg [31:0] eq_266_in0;
	reg [31:0] eq_266_in1;
	wire [0:0] eq_266_out;
	eq #(.WIDTH(32)) eq_266(.in0(eq_266_in0), .in1(eq_266_in1), .out(eq_266_out));

	reg [0:0] andOp_267_in0;
	reg [0:0] andOp_267_in1;
	wire [0:0] andOp_267_out;
	andOp #(.WIDTH(1)) andOp_267(.in0(andOp_267_in0), .in1(andOp_267_in1), .out(andOp_267_out));

	reg [31:0] eq_268_in0;
	reg [31:0] eq_268_in1;
	wire [0:0] eq_268_out;
	eq #(.WIDTH(32)) eq_268(.in0(eq_268_in0), .in1(eq_268_in1), .out(eq_268_out));

	reg [0:0] andOp_269_in0;
	reg [0:0] andOp_269_in1;
	wire [0:0] andOp_269_out;
	andOp #(.WIDTH(1)) andOp_269(.in0(andOp_269_in0), .in1(andOp_269_in1), .out(andOp_269_out));

	reg [0:0] notOp_270_in0;
	wire [0:0] notOp_270_out;
	notOp #(.WIDTH(1)) notOp_270(.in(notOp_270_in0), .out(notOp_270_out));

	reg [0:0] andOp_271_in0;
	reg [0:0] andOp_271_in1;
	wire [0:0] andOp_271_out;
	andOp #(.WIDTH(1)) andOp_271(.in0(andOp_271_in0), .in1(andOp_271_in1), .out(andOp_271_out));

	reg [0:0] notOp_272_in0;
	wire [0:0] notOp_272_out;
	notOp #(.WIDTH(1)) notOp_272(.in(notOp_272_in0), .out(notOp_272_out));

	reg [0:0] andOp_273_in0;
	reg [0:0] andOp_273_in1;
	wire [0:0] andOp_273_out;
	andOp #(.WIDTH(1)) andOp_273(.in0(andOp_273_in0), .in1(andOp_273_in1), .out(andOp_273_out));

	reg [0:0] notOp_274_in0;
	wire [0:0] notOp_274_out;
	notOp #(.WIDTH(1)) notOp_274(.in(notOp_274_in0), .out(notOp_274_out));

	reg [0:0] andOp_275_in0;
	reg [0:0] andOp_275_in1;
	wire [0:0] andOp_275_out;
	andOp #(.WIDTH(1)) andOp_275(.in0(andOp_275_in0), .in1(andOp_275_in1), .out(andOp_275_out));

	reg [0:0] andOp_276_in0;
	reg [0:0] andOp_276_in1;
	wire [0:0] andOp_276_out;
	andOp #(.WIDTH(1)) andOp_276(.in0(andOp_276_in0), .in1(andOp_276_in1), .out(andOp_276_out));

	reg [31:0] eq_277_in0;
	reg [31:0] eq_277_in1;
	wire [0:0] eq_277_out;
	eq #(.WIDTH(32)) eq_277(.in0(eq_277_in0), .in1(eq_277_in1), .out(eq_277_out));

	reg [0:0] andOp_278_in0;
	reg [0:0] andOp_278_in1;
	wire [0:0] andOp_278_out;
	andOp #(.WIDTH(1)) andOp_278(.in0(andOp_278_in0), .in1(andOp_278_in1), .out(andOp_278_out));

	reg [0:0] notOp_279_in0;
	wire [0:0] notOp_279_out;
	notOp #(.WIDTH(1)) notOp_279(.in(notOp_279_in0), .out(notOp_279_out));

	reg [0:0] andOp_280_in0;
	reg [0:0] andOp_280_in1;
	wire [0:0] andOp_280_out;
	andOp #(.WIDTH(1)) andOp_280(.in0(andOp_280_in0), .in1(andOp_280_in1), .out(andOp_280_out));

	reg [0:0] notOp_281_in0;
	wire [0:0] notOp_281_out;
	notOp #(.WIDTH(1)) notOp_281(.in(notOp_281_in0), .out(notOp_281_out));

	reg [0:0] andOp_282_in0;
	reg [0:0] andOp_282_in1;
	wire [0:0] andOp_282_out;
	andOp #(.WIDTH(1)) andOp_282(.in0(andOp_282_in0), .in1(andOp_282_in1), .out(andOp_282_out));

	reg [0:0] notOp_283_in0;
	wire [0:0] notOp_283_out;
	notOp #(.WIDTH(1)) notOp_283(.in(notOp_283_in0), .out(notOp_283_out));

	reg [0:0] andOp_284_in0;
	reg [0:0] andOp_284_in1;
	wire [0:0] andOp_284_out;
	andOp #(.WIDTH(1)) andOp_284(.in0(andOp_284_in0), .in1(andOp_284_in1), .out(andOp_284_out));

	reg [0:0] andOp_285_in0;
	reg [0:0] andOp_285_in1;
	wire [0:0] andOp_285_out;
	andOp #(.WIDTH(1)) andOp_285(.in0(andOp_285_in0), .in1(andOp_285_in1), .out(andOp_285_out));

	reg [31:0] eq_286_in0;
	reg [31:0] eq_286_in1;
	wire [0:0] eq_286_out;
	eq #(.WIDTH(32)) eq_286(.in0(eq_286_in0), .in1(eq_286_in1), .out(eq_286_out));

	reg [0:0] andOp_287_in0;
	reg [0:0] andOp_287_in1;
	wire [0:0] andOp_287_out;
	andOp #(.WIDTH(1)) andOp_287(.in0(andOp_287_in0), .in1(andOp_287_in1), .out(andOp_287_out));

	reg [0:0] notOp_288_in0;
	wire [0:0] notOp_288_out;
	notOp #(.WIDTH(1)) notOp_288(.in(notOp_288_in0), .out(notOp_288_out));

	reg [0:0] andOp_289_in0;
	reg [0:0] andOp_289_in1;
	wire [0:0] andOp_289_out;
	andOp #(.WIDTH(1)) andOp_289(.in0(andOp_289_in0), .in1(andOp_289_in1), .out(andOp_289_out));

	reg [0:0] notOp_290_in0;
	wire [0:0] notOp_290_out;
	notOp #(.WIDTH(1)) notOp_290(.in(notOp_290_in0), .out(notOp_290_out));

	reg [0:0] andOp_291_in0;
	reg [0:0] andOp_291_in1;
	wire [0:0] andOp_291_out;
	andOp #(.WIDTH(1)) andOp_291(.in0(andOp_291_in0), .in1(andOp_291_in1), .out(andOp_291_out));

	reg [0:0] notOp_292_in0;
	wire [0:0] notOp_292_out;
	notOp #(.WIDTH(1)) notOp_292(.in(notOp_292_in0), .out(notOp_292_out));

	reg [0:0] andOp_293_in0;
	reg [0:0] andOp_293_in1;
	wire [0:0] andOp_293_out;
	andOp #(.WIDTH(1)) andOp_293(.in0(andOp_293_in0), .in1(andOp_293_in1), .out(andOp_293_out));

	reg [0:0] andOp_294_in0;
	reg [0:0] andOp_294_in1;
	wire [0:0] andOp_294_out;
	andOp #(.WIDTH(1)) andOp_294(.in0(andOp_294_in0), .in1(andOp_294_in1), .out(andOp_294_out));

	reg [31:0] eq_295_in0;
	reg [31:0] eq_295_in1;
	wire [0:0] eq_295_out;
	eq #(.WIDTH(32)) eq_295(.in0(eq_295_in0), .in1(eq_295_in1), .out(eq_295_out));

	reg [0:0] andOp_296_in0;
	reg [0:0] andOp_296_in1;
	wire [0:0] andOp_296_out;
	andOp #(.WIDTH(1)) andOp_296(.in0(andOp_296_in0), .in1(andOp_296_in1), .out(andOp_296_out));

	reg [0:0] notOp_297_in0;
	wire [0:0] notOp_297_out;
	notOp #(.WIDTH(1)) notOp_297(.in(notOp_297_in0), .out(notOp_297_out));

	reg [0:0] andOp_298_in0;
	reg [0:0] andOp_298_in1;
	wire [0:0] andOp_298_out;
	andOp #(.WIDTH(1)) andOp_298(.in0(andOp_298_in0), .in1(andOp_298_in1), .out(andOp_298_out));

	reg [0:0] notOp_299_in0;
	wire [0:0] notOp_299_out;
	notOp #(.WIDTH(1)) notOp_299(.in(notOp_299_in0), .out(notOp_299_out));

	reg [0:0] andOp_300_in0;
	reg [0:0] andOp_300_in1;
	wire [0:0] andOp_300_out;
	andOp #(.WIDTH(1)) andOp_300(.in0(andOp_300_in0), .in1(andOp_300_in1), .out(andOp_300_out));

	reg [0:0] notOp_301_in0;
	wire [0:0] notOp_301_out;
	notOp #(.WIDTH(1)) notOp_301(.in(notOp_301_in0), .out(notOp_301_out));

	reg [0:0] andOp_302_in0;
	reg [0:0] andOp_302_in1;
	wire [0:0] andOp_302_out;
	andOp #(.WIDTH(1)) andOp_302(.in0(andOp_302_in0), .in1(andOp_302_in1), .out(andOp_302_out));

	reg [31:0] eq_303_in0;
	reg [31:0] eq_303_in1;
	wire [0:0] eq_303_out;
	eq #(.WIDTH(32)) eq_303(.in0(eq_303_in0), .in1(eq_303_in1), .out(eq_303_out));

	reg [31:0] eq_304_in0;
	reg [31:0] eq_304_in1;
	wire [0:0] eq_304_out;
	eq #(.WIDTH(32)) eq_304(.in0(eq_304_in0), .in1(eq_304_in1), .out(eq_304_out));

	reg [0:0] andOp_305_in0;
	reg [0:0] andOp_305_in1;
	wire [0:0] andOp_305_out;
	andOp #(.WIDTH(1)) andOp_305(.in0(andOp_305_in0), .in1(andOp_305_in1), .out(andOp_305_out));

	reg [31:0] eq_306_in0;
	reg [31:0] eq_306_in1;
	wire [0:0] eq_306_out;
	eq #(.WIDTH(32)) eq_306(.in0(eq_306_in0), .in1(eq_306_in1), .out(eq_306_out));

	reg [0:0] andOp_307_in0;
	reg [0:0] andOp_307_in1;
	wire [0:0] andOp_307_out;
	andOp #(.WIDTH(1)) andOp_307(.in0(andOp_307_in0), .in1(andOp_307_in1), .out(andOp_307_out));

	reg [0:0] notOp_308_in0;
	wire [0:0] notOp_308_out;
	notOp #(.WIDTH(1)) notOp_308(.in(notOp_308_in0), .out(notOp_308_out));

	reg [0:0] andOp_309_in0;
	reg [0:0] andOp_309_in1;
	wire [0:0] andOp_309_out;
	andOp #(.WIDTH(1)) andOp_309(.in0(andOp_309_in0), .in1(andOp_309_in1), .out(andOp_309_out));

	reg [0:0] notOp_310_in0;
	wire [0:0] notOp_310_out;
	notOp #(.WIDTH(1)) notOp_310(.in(notOp_310_in0), .out(notOp_310_out));

	reg [0:0] andOp_311_in0;
	reg [0:0] andOp_311_in1;
	wire [0:0] andOp_311_out;
	andOp #(.WIDTH(1)) andOp_311(.in0(andOp_311_in0), .in1(andOp_311_in1), .out(andOp_311_out));

	reg [0:0] notOp_312_in0;
	wire [0:0] notOp_312_out;
	notOp #(.WIDTH(1)) notOp_312(.in(notOp_312_in0), .out(notOp_312_out));

	reg [0:0] andOp_313_in0;
	reg [0:0] andOp_313_in1;
	wire [0:0] andOp_313_out;
	andOp #(.WIDTH(1)) andOp_313(.in0(andOp_313_in0), .in1(andOp_313_in1), .out(andOp_313_out));

	reg [0:0] andOp_314_in0;
	reg [0:0] andOp_314_in1;
	wire [0:0] andOp_314_out;
	andOp #(.WIDTH(1)) andOp_314(.in0(andOp_314_in0), .in1(andOp_314_in1), .out(andOp_314_out));

	reg [31:0] eq_315_in0;
	reg [31:0] eq_315_in1;
	wire [0:0] eq_315_out;
	eq #(.WIDTH(32)) eq_315(.in0(eq_315_in0), .in1(eq_315_in1), .out(eq_315_out));

	reg [0:0] andOp_316_in0;
	reg [0:0] andOp_316_in1;
	wire [0:0] andOp_316_out;
	andOp #(.WIDTH(1)) andOp_316(.in0(andOp_316_in0), .in1(andOp_316_in1), .out(andOp_316_out));

	reg [0:0] notOp_317_in0;
	wire [0:0] notOp_317_out;
	notOp #(.WIDTH(1)) notOp_317(.in(notOp_317_in0), .out(notOp_317_out));

	reg [0:0] andOp_318_in0;
	reg [0:0] andOp_318_in1;
	wire [0:0] andOp_318_out;
	andOp #(.WIDTH(1)) andOp_318(.in0(andOp_318_in0), .in1(andOp_318_in1), .out(andOp_318_out));

	reg [0:0] notOp_319_in0;
	wire [0:0] notOp_319_out;
	notOp #(.WIDTH(1)) notOp_319(.in(notOp_319_in0), .out(notOp_319_out));

	reg [0:0] andOp_320_in0;
	reg [0:0] andOp_320_in1;
	wire [0:0] andOp_320_out;
	andOp #(.WIDTH(1)) andOp_320(.in0(andOp_320_in0), .in1(andOp_320_in1), .out(andOp_320_out));

	reg [0:0] notOp_321_in0;
	wire [0:0] notOp_321_out;
	notOp #(.WIDTH(1)) notOp_321(.in(notOp_321_in0), .out(notOp_321_out));

	reg [0:0] andOp_322_in0;
	reg [0:0] andOp_322_in1;
	wire [0:0] andOp_322_out;
	andOp #(.WIDTH(1)) andOp_322(.in0(andOp_322_in0), .in1(andOp_322_in1), .out(andOp_322_out));

	reg [0:0] andOp_323_in0;
	reg [0:0] andOp_323_in1;
	wire [0:0] andOp_323_out;
	andOp #(.WIDTH(1)) andOp_323(.in0(andOp_323_in0), .in1(andOp_323_in1), .out(andOp_323_out));

	reg [31:0] eq_324_in0;
	reg [31:0] eq_324_in1;
	wire [0:0] eq_324_out;
	eq #(.WIDTH(32)) eq_324(.in0(eq_324_in0), .in1(eq_324_in1), .out(eq_324_out));

	reg [0:0] andOp_325_in0;
	reg [0:0] andOp_325_in1;
	wire [0:0] andOp_325_out;
	andOp #(.WIDTH(1)) andOp_325(.in0(andOp_325_in0), .in1(andOp_325_in1), .out(andOp_325_out));

	reg [0:0] notOp_326_in0;
	wire [0:0] notOp_326_out;
	notOp #(.WIDTH(1)) notOp_326(.in(notOp_326_in0), .out(notOp_326_out));

	reg [0:0] andOp_327_in0;
	reg [0:0] andOp_327_in1;
	wire [0:0] andOp_327_out;
	andOp #(.WIDTH(1)) andOp_327(.in0(andOp_327_in0), .in1(andOp_327_in1), .out(andOp_327_out));

	reg [0:0] notOp_328_in0;
	wire [0:0] notOp_328_out;
	notOp #(.WIDTH(1)) notOp_328(.in(notOp_328_in0), .out(notOp_328_out));

	reg [0:0] andOp_329_in0;
	reg [0:0] andOp_329_in1;
	wire [0:0] andOp_329_out;
	andOp #(.WIDTH(1)) andOp_329(.in0(andOp_329_in0), .in1(andOp_329_in1), .out(andOp_329_out));

	reg [0:0] notOp_330_in0;
	wire [0:0] notOp_330_out;
	notOp #(.WIDTH(1)) notOp_330(.in(notOp_330_in0), .out(notOp_330_out));

	reg [0:0] andOp_331_in0;
	reg [0:0] andOp_331_in1;
	wire [0:0] andOp_331_out;
	andOp #(.WIDTH(1)) andOp_331(.in0(andOp_331_in0), .in1(andOp_331_in1), .out(andOp_331_out));

	reg [0:0] andOp_332_in0;
	reg [0:0] andOp_332_in1;
	wire [0:0] andOp_332_out;
	andOp #(.WIDTH(1)) andOp_332(.in0(andOp_332_in0), .in1(andOp_332_in1), .out(andOp_332_out));

	reg [31:0] eq_333_in0;
	reg [31:0] eq_333_in1;
	wire [0:0] eq_333_out;
	eq #(.WIDTH(32)) eq_333(.in0(eq_333_in0), .in1(eq_333_in1), .out(eq_333_out));

	reg [0:0] andOp_334_in0;
	reg [0:0] andOp_334_in1;
	wire [0:0] andOp_334_out;
	andOp #(.WIDTH(1)) andOp_334(.in0(andOp_334_in0), .in1(andOp_334_in1), .out(andOp_334_out));

	reg [0:0] notOp_335_in0;
	wire [0:0] notOp_335_out;
	notOp #(.WIDTH(1)) notOp_335(.in(notOp_335_in0), .out(notOp_335_out));

	reg [0:0] andOp_336_in0;
	reg [0:0] andOp_336_in1;
	wire [0:0] andOp_336_out;
	andOp #(.WIDTH(1)) andOp_336(.in0(andOp_336_in0), .in1(andOp_336_in1), .out(andOp_336_out));

	reg [0:0] notOp_337_in0;
	wire [0:0] notOp_337_out;
	notOp #(.WIDTH(1)) notOp_337(.in(notOp_337_in0), .out(notOp_337_out));

	reg [0:0] andOp_338_in0;
	reg [0:0] andOp_338_in1;
	wire [0:0] andOp_338_out;
	andOp #(.WIDTH(1)) andOp_338(.in0(andOp_338_in0), .in1(andOp_338_in1), .out(andOp_338_out));

	reg [0:0] notOp_339_in0;
	wire [0:0] notOp_339_out;
	notOp #(.WIDTH(1)) notOp_339(.in(notOp_339_in0), .out(notOp_339_out));

	reg [0:0] andOp_340_in0;
	reg [0:0] andOp_340_in1;
	wire [0:0] andOp_340_out;
	andOp #(.WIDTH(1)) andOp_340(.in0(andOp_340_in0), .in1(andOp_340_in1), .out(andOp_340_out));

	reg [31:0] eq_341_in0;
	reg [31:0] eq_341_in1;
	wire [0:0] eq_341_out;
	eq #(.WIDTH(32)) eq_341(.in0(eq_341_in0), .in1(eq_341_in1), .out(eq_341_out));

	reg [31:0] eq_342_in0;
	reg [31:0] eq_342_in1;
	wire [0:0] eq_342_out;
	eq #(.WIDTH(32)) eq_342(.in0(eq_342_in0), .in1(eq_342_in1), .out(eq_342_out));

	reg [0:0] andOp_343_in0;
	reg [0:0] andOp_343_in1;
	wire [0:0] andOp_343_out;
	andOp #(.WIDTH(1)) andOp_343(.in0(andOp_343_in0), .in1(andOp_343_in1), .out(andOp_343_out));

	reg [31:0] eq_344_in0;
	reg [31:0] eq_344_in1;
	wire [0:0] eq_344_out;
	eq #(.WIDTH(32)) eq_344(.in0(eq_344_in0), .in1(eq_344_in1), .out(eq_344_out));

	reg [0:0] andOp_345_in0;
	reg [0:0] andOp_345_in1;
	wire [0:0] andOp_345_out;
	andOp #(.WIDTH(1)) andOp_345(.in0(andOp_345_in0), .in1(andOp_345_in1), .out(andOp_345_out));

	reg [0:0] notOp_346_in0;
	wire [0:0] notOp_346_out;
	notOp #(.WIDTH(1)) notOp_346(.in(notOp_346_in0), .out(notOp_346_out));

	reg [0:0] andOp_347_in0;
	reg [0:0] andOp_347_in1;
	wire [0:0] andOp_347_out;
	andOp #(.WIDTH(1)) andOp_347(.in0(andOp_347_in0), .in1(andOp_347_in1), .out(andOp_347_out));

	reg [0:0] notOp_348_in0;
	wire [0:0] notOp_348_out;
	notOp #(.WIDTH(1)) notOp_348(.in(notOp_348_in0), .out(notOp_348_out));

	reg [0:0] andOp_349_in0;
	reg [0:0] andOp_349_in1;
	wire [0:0] andOp_349_out;
	andOp #(.WIDTH(1)) andOp_349(.in0(andOp_349_in0), .in1(andOp_349_in1), .out(andOp_349_out));

	reg [0:0] notOp_350_in0;
	wire [0:0] notOp_350_out;
	notOp #(.WIDTH(1)) notOp_350(.in(notOp_350_in0), .out(notOp_350_out));

	reg [0:0] andOp_351_in0;
	reg [0:0] andOp_351_in1;
	wire [0:0] andOp_351_out;
	andOp #(.WIDTH(1)) andOp_351(.in0(andOp_351_in0), .in1(andOp_351_in1), .out(andOp_351_out));

	reg [0:0] andOp_352_in0;
	reg [0:0] andOp_352_in1;
	wire [0:0] andOp_352_out;
	andOp #(.WIDTH(1)) andOp_352(.in0(andOp_352_in0), .in1(andOp_352_in1), .out(andOp_352_out));

	reg [31:0] eq_353_in0;
	reg [31:0] eq_353_in1;
	wire [0:0] eq_353_out;
	eq #(.WIDTH(32)) eq_353(.in0(eq_353_in0), .in1(eq_353_in1), .out(eq_353_out));

	reg [0:0] andOp_354_in0;
	reg [0:0] andOp_354_in1;
	wire [0:0] andOp_354_out;
	andOp #(.WIDTH(1)) andOp_354(.in0(andOp_354_in0), .in1(andOp_354_in1), .out(andOp_354_out));

	reg [0:0] notOp_355_in0;
	wire [0:0] notOp_355_out;
	notOp #(.WIDTH(1)) notOp_355(.in(notOp_355_in0), .out(notOp_355_out));

	reg [0:0] andOp_356_in0;
	reg [0:0] andOp_356_in1;
	wire [0:0] andOp_356_out;
	andOp #(.WIDTH(1)) andOp_356(.in0(andOp_356_in0), .in1(andOp_356_in1), .out(andOp_356_out));

	reg [0:0] notOp_357_in0;
	wire [0:0] notOp_357_out;
	notOp #(.WIDTH(1)) notOp_357(.in(notOp_357_in0), .out(notOp_357_out));

	reg [0:0] andOp_358_in0;
	reg [0:0] andOp_358_in1;
	wire [0:0] andOp_358_out;
	andOp #(.WIDTH(1)) andOp_358(.in0(andOp_358_in0), .in1(andOp_358_in1), .out(andOp_358_out));

	reg [0:0] notOp_359_in0;
	wire [0:0] notOp_359_out;
	notOp #(.WIDTH(1)) notOp_359(.in(notOp_359_in0), .out(notOp_359_out));

	reg [0:0] andOp_360_in0;
	reg [0:0] andOp_360_in1;
	wire [0:0] andOp_360_out;
	andOp #(.WIDTH(1)) andOp_360(.in0(andOp_360_in0), .in1(andOp_360_in1), .out(andOp_360_out));

	reg [0:0] andOp_361_in0;
	reg [0:0] andOp_361_in1;
	wire [0:0] andOp_361_out;
	andOp #(.WIDTH(1)) andOp_361(.in0(andOp_361_in0), .in1(andOp_361_in1), .out(andOp_361_out));

	reg [31:0] eq_362_in0;
	reg [31:0] eq_362_in1;
	wire [0:0] eq_362_out;
	eq #(.WIDTH(32)) eq_362(.in0(eq_362_in0), .in1(eq_362_in1), .out(eq_362_out));

	reg [0:0] andOp_363_in0;
	reg [0:0] andOp_363_in1;
	wire [0:0] andOp_363_out;
	andOp #(.WIDTH(1)) andOp_363(.in0(andOp_363_in0), .in1(andOp_363_in1), .out(andOp_363_out));

	reg [0:0] notOp_364_in0;
	wire [0:0] notOp_364_out;
	notOp #(.WIDTH(1)) notOp_364(.in(notOp_364_in0), .out(notOp_364_out));

	reg [0:0] andOp_365_in0;
	reg [0:0] andOp_365_in1;
	wire [0:0] andOp_365_out;
	andOp #(.WIDTH(1)) andOp_365(.in0(andOp_365_in0), .in1(andOp_365_in1), .out(andOp_365_out));

	reg [0:0] notOp_366_in0;
	wire [0:0] notOp_366_out;
	notOp #(.WIDTH(1)) notOp_366(.in(notOp_366_in0), .out(notOp_366_out));

	reg [0:0] andOp_367_in0;
	reg [0:0] andOp_367_in1;
	wire [0:0] andOp_367_out;
	andOp #(.WIDTH(1)) andOp_367(.in0(andOp_367_in0), .in1(andOp_367_in1), .out(andOp_367_out));

	reg [0:0] notOp_368_in0;
	wire [0:0] notOp_368_out;
	notOp #(.WIDTH(1)) notOp_368(.in(notOp_368_in0), .out(notOp_368_out));

	reg [0:0] andOp_369_in0;
	reg [0:0] andOp_369_in1;
	wire [0:0] andOp_369_out;
	andOp #(.WIDTH(1)) andOp_369(.in0(andOp_369_in0), .in1(andOp_369_in1), .out(andOp_369_out));

	reg [0:0] andOp_370_in0;
	reg [0:0] andOp_370_in1;
	wire [0:0] andOp_370_out;
	andOp #(.WIDTH(1)) andOp_370(.in0(andOp_370_in0), .in1(andOp_370_in1), .out(andOp_370_out));

	reg [31:0] eq_371_in0;
	reg [31:0] eq_371_in1;
	wire [0:0] eq_371_out;
	eq #(.WIDTH(32)) eq_371(.in0(eq_371_in0), .in1(eq_371_in1), .out(eq_371_out));

	reg [0:0] andOp_372_in0;
	reg [0:0] andOp_372_in1;
	wire [0:0] andOp_372_out;
	andOp #(.WIDTH(1)) andOp_372(.in0(andOp_372_in0), .in1(andOp_372_in1), .out(andOp_372_out));

	reg [0:0] notOp_373_in0;
	wire [0:0] notOp_373_out;
	notOp #(.WIDTH(1)) notOp_373(.in(notOp_373_in0), .out(notOp_373_out));

	reg [0:0] andOp_374_in0;
	reg [0:0] andOp_374_in1;
	wire [0:0] andOp_374_out;
	andOp #(.WIDTH(1)) andOp_374(.in0(andOp_374_in0), .in1(andOp_374_in1), .out(andOp_374_out));

	reg [0:0] notOp_375_in0;
	wire [0:0] notOp_375_out;
	notOp #(.WIDTH(1)) notOp_375(.in(notOp_375_in0), .out(notOp_375_out));

	reg [0:0] andOp_376_in0;
	reg [0:0] andOp_376_in1;
	wire [0:0] andOp_376_out;
	andOp #(.WIDTH(1)) andOp_376(.in0(andOp_376_in0), .in1(andOp_376_in1), .out(andOp_376_out));

	reg [0:0] notOp_377_in0;
	wire [0:0] notOp_377_out;
	notOp #(.WIDTH(1)) notOp_377(.in(notOp_377_in0), .out(notOp_377_out));

	reg [0:0] andOp_378_in0;
	reg [0:0] andOp_378_in1;
	wire [0:0] andOp_378_out;
	andOp #(.WIDTH(1)) andOp_378(.in0(andOp_378_in0), .in1(andOp_378_in1), .out(andOp_378_out));

	// End Functional Units

	reg [31:0] data_store_0_0;
	reg [31:0] data_store_0_2;
	reg [31:0] data_store_0_4;
	reg [0:0] data_store_0_6;
	reg [31:0] data_store_1_10;
	reg [31:0] data_store_1_12;
	reg [0:0] data_store_1_14;
	reg [31:0] data_store_1_8;
	reg [31:0] data_store_2_16;
	reg [31:0] data_store_2_18;
	reg [31:0] data_store_2_20;
	reg [0:0] data_store_2_22;
	reg [31:0] data_store_3_24;
	reg [31:0] data_store_3_26;
	reg [31:0] data_store_3_28;
	reg [0:0] data_store_3_30;
	reg [31:0] data_store_4_32;
	reg [31:0] data_store_4_34;
	reg [31:0] data_store_4_36;
	reg [0:0] data_store_4_38;
	reg [31:0] global_state;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_3_last_state;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;
	reg [31:0] state_4_last_state;

	// controller for add_add_14.add_in0_add_14
	// controller for add_add_14.add_in1_add_14
	// Insensitive connections
	always @(*) begin
		add_in0_add_14 = valid ? rdata_ram_0 : rdata_ram_0;
		add_in1_add_14 = valid ? tmp_output_160_out_data : tmp_output_160_out_data;
	end
	// controller for add_add_16.add_in0_add_16
	// controller for add_add_16.add_in1_add_16
	// Insensitive connections
	always @(*) begin
		add_in0_add_16 = valid ? data_in_3_27_out_data : data_in_3_27_out_data;
		add_in1_add_16 = valid ? 32'd1 : 32'd1;
	end
	// controller for andOp_117.andOp_117_in0
	// controller for andOp_117.andOp_117_in1
	// Insensitive connections
	always @(*) begin
		andOp_117_in0 = valid ? notOp_116_out : notOp_116_out;
		andOp_117_in1 = valid ? andOp_56_out : andOp_56_out;
	end
	// controller for andOp_120.andOp_120_in0
	// controller for andOp_120.andOp_120_in1
	// Insensitive connections
	always @(*) begin
		andOp_120_in0 = valid ? notOp_119_out : notOp_119_out;
		andOp_120_in1 = valid ? andOp_44_out : andOp_44_out;
	end
	// controller for andOp_124.andOp_124_in0
	// controller for andOp_124.andOp_124_in1
	// Insensitive connections
	always @(*) begin
		andOp_124_in0 = valid ? notOp_123_out : notOp_123_out;
		andOp_124_in1 = valid ? andOp_41_out : andOp_41_out;
	end
	// controller for andOp_128.andOp_128_in0
	// controller for andOp_128.andOp_128_in1
	// Insensitive connections
	always @(*) begin
		andOp_128_in0 = valid ? notOp_127_out : notOp_127_out;
		andOp_128_in1 = valid ? andOp_59_out : andOp_59_out;
	end
	// controller for andOp_132.andOp_132_in0
	// controller for andOp_132.andOp_132_in1
	// Insensitive connections
	always @(*) begin
		andOp_132_in0 = valid ? notOp_131_out : notOp_131_out;
		andOp_132_in1 = valid ? andOp_74_out : andOp_74_out;
	end
	// controller for andOp_135.andOp_135_in0
	// controller for andOp_135.andOp_135_in1
	// Insensitive connections
	always @(*) begin
		andOp_135_in0 = valid ? notOp_134_out : notOp_134_out;
		andOp_135_in1 = valid ? andOp_89_out : andOp_89_out;
	end
	// controller for andOp_138.andOp_138_in0
	// controller for andOp_138.andOp_138_in1
	// Insensitive connections
	always @(*) begin
		andOp_138_in0 = valid ? notOp_137_out : notOp_137_out;
		andOp_138_in1 = valid ? andOp_79_out : andOp_79_out;
	end
	// controller for andOp_141.andOp_141_in0
	// controller for andOp_141.andOp_141_in1
	// Insensitive connections
	always @(*) begin
		andOp_141_in0 = valid ? notOp_140_out : notOp_140_out;
		andOp_141_in1 = valid ? andOp_71_out : andOp_71_out;
	end
	// controller for andOp_145.andOp_145_in0
	// controller for andOp_145.andOp_145_in1
	// Insensitive connections
	always @(*) begin
		andOp_145_in0 = valid ? notOp_144_out : notOp_144_out;
		andOp_145_in1 = valid ? andOp_64_out : andOp_64_out;
	end
	// controller for andOp_146.andOp_146_in0
	// controller for andOp_146.andOp_146_in1
	// Insensitive connections
	always @(*) begin
		andOp_146_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_146_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_147.andOp_147_in0
	// controller for andOp_147.andOp_147_in1
	// Insensitive connections
	always @(*) begin
		andOp_147_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_147_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_148.andOp_148_in0
	// controller for andOp_148.andOp_148_in1
	// Insensitive connections
	always @(*) begin
		andOp_148_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_148_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_149.andOp_149_in0
	// controller for andOp_149.andOp_149_in1
	// Insensitive connections
	always @(*) begin
		andOp_149_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_149_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_150.andOp_150_in0
	// controller for andOp_150.andOp_150_in1
	// Insensitive connections
	always @(*) begin
		andOp_150_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_150_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_151.andOp_151_in0
	// controller for andOp_151.andOp_151_in1
	// Insensitive connections
	always @(*) begin
		andOp_151_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_151_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_152.andOp_152_in0
	// controller for andOp_152.andOp_152_in1
	// Insensitive connections
	always @(*) begin
		andOp_152_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_152_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_153.andOp_153_in0
	// controller for andOp_153.andOp_153_in1
	// Insensitive connections
	always @(*) begin
		andOp_153_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
		andOp_153_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_154.andOp_154_in0
	// controller for andOp_154.andOp_154_in1
	// Insensitive connections
	always @(*) begin
		andOp_154_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_154_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_155.andOp_155_in0
	// controller for andOp_155.andOp_155_in1
	// Insensitive connections
	always @(*) begin
		andOp_155_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_155_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_156.andOp_156_in0
	// controller for andOp_156.andOp_156_in1
	// Insensitive connections
	always @(*) begin
		andOp_156_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_156_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_159.andOp_159_in0
	// controller for andOp_159.andOp_159_in1
	// Insensitive connections
	always @(*) begin
		andOp_159_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_159_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_162.andOp_162_in0
	// controller for andOp_162.andOp_162_in1
	// Insensitive connections
	always @(*) begin
		andOp_162_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_162_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_163.andOp_163_in0
	// controller for andOp_163.andOp_163_in1
	// Insensitive connections
	always @(*) begin
		andOp_163_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_163_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_164.andOp_164_in0
	// controller for andOp_164.andOp_164_in1
	// Insensitive connections
	always @(*) begin
		andOp_164_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
		andOp_164_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_165.andOp_165_in0
	// controller for andOp_165.andOp_165_in1
	// Insensitive connections
	always @(*) begin
		andOp_165_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_165_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_166.andOp_166_in0
	// controller for andOp_166.andOp_166_in1
	// Insensitive connections
	always @(*) begin
		andOp_166_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_166_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_167.andOp_167_in0
	// controller for andOp_167.andOp_167_in1
	// Insensitive connections
	always @(*) begin
		andOp_167_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_167_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_168.andOp_168_in0
	// controller for andOp_168.andOp_168_in1
	// Insensitive connections
	always @(*) begin
		andOp_168_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_168_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_169.andOp_169_in0
	// controller for andOp_169.andOp_169_in1
	// Insensitive connections
	always @(*) begin
		andOp_169_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_169_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_170.andOp_170_in0
	// controller for andOp_170.andOp_170_in1
	// Insensitive connections
	always @(*) begin
		andOp_170_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_170_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_171.andOp_171_in0
	// controller for andOp_171.andOp_171_in1
	// Insensitive connections
	always @(*) begin
		andOp_171_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_171_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_172.andOp_172_in0
	// controller for andOp_172.andOp_172_in1
	// Insensitive connections
	always @(*) begin
		andOp_172_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_172_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_174.andOp_174_in0
	// controller for andOp_174.andOp_174_in1
	// Insensitive connections
	always @(*) begin
		andOp_174_in0 = valid ? notOp_173_out : notOp_173_out;
		andOp_174_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_176.andOp_176_in0
	// controller for andOp_176.andOp_176_in1
	// Insensitive connections
	always @(*) begin
		andOp_176_in0 = valid ? notOp_175_out : notOp_175_out;
		andOp_176_in1 = valid ? andOp_174_out : andOp_174_out;
	end
	// controller for andOp_178.andOp_178_in0
	// controller for andOp_178.andOp_178_in1
	// Insensitive connections
	always @(*) begin
		andOp_178_in0 = valid ? notOp_177_out : notOp_177_out;
		andOp_178_in1 = valid ? andOp_176_out : andOp_176_out;
	end
	// controller for andOp_180.andOp_180_in0
	// controller for andOp_180.andOp_180_in1
	// Insensitive connections
	always @(*) begin
		andOp_180_in0 = valid ? notOp_179_out : notOp_179_out;
		andOp_180_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_182.andOp_182_in0
	// controller for andOp_182.andOp_182_in1
	// Insensitive connections
	always @(*) begin
		andOp_182_in0 = valid ? notOp_181_out : notOp_181_out;
		andOp_182_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_184.andOp_184_in0
	// controller for andOp_184.andOp_184_in1
	// Insensitive connections
	always @(*) begin
		andOp_184_in0 = valid ? notOp_183_out : notOp_183_out;
		andOp_184_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_186.andOp_186_in0
	// controller for andOp_186.andOp_186_in1
	// Insensitive connections
	always @(*) begin
		andOp_186_in0 = valid ? notOp_185_out : notOp_185_out;
		andOp_186_in1 = valid ? andOp_184_out : andOp_184_out;
	end
	// controller for andOp_188.andOp_188_in0
	// controller for andOp_188.andOp_188_in1
	// Insensitive connections
	always @(*) begin
		andOp_188_in0 = valid ? notOp_187_out : notOp_187_out;
		andOp_188_in1 = valid ? andOp_186_out : andOp_186_out;
	end
	// controller for andOp_190.andOp_190_in0
	// controller for andOp_190.andOp_190_in1
	// Insensitive connections
	always @(*) begin
		andOp_190_in0 = valid ? 1'd0 : 1'd0;
		andOp_190_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_192.andOp_192_in0
	// controller for andOp_192.andOp_192_in1
	// Insensitive connections
	always @(*) begin
		andOp_192_in0 = valid ? andOp_190_out : andOp_190_out;
		andOp_192_in1 = valid ? eq_191_out : eq_191_out;
	end
	// controller for andOp_194.andOp_194_in0
	// controller for andOp_194.andOp_194_in1
	// Insensitive connections
	always @(*) begin
		andOp_194_in0 = valid ? andOp_190_out : andOp_190_out;
		andOp_194_in1 = valid ? notOp_193_out : notOp_193_out;
	end
	// controller for andOp_196.andOp_196_in0
	// controller for andOp_196.andOp_196_in1
	// Insensitive connections
	always @(*) begin
		andOp_196_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_196_in1 = valid ? notOp_195_out : notOp_195_out;
	end
	// controller for andOp_198.andOp_198_in0
	// controller for andOp_198.andOp_198_in1
	// Insensitive connections
	always @(*) begin
		andOp_198_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_198_in1 = valid ? notOp_197_out : notOp_197_out;
	end
	// controller for andOp_199.andOp_199_in0
	// controller for andOp_199.andOp_199_in1
	// Insensitive connections
	always @(*) begin
		andOp_199_in0 = valid ? 1'd0 : 1'd0;
		andOp_199_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_201.andOp_201_in0
	// controller for andOp_201.andOp_201_in1
	// Insensitive connections
	always @(*) begin
		andOp_201_in0 = valid ? andOp_199_out : andOp_199_out;
		andOp_201_in1 = valid ? eq_200_out : eq_200_out;
	end
	// controller for andOp_203.andOp_203_in0
	// controller for andOp_203.andOp_203_in1
	// Insensitive connections
	always @(*) begin
		andOp_203_in0 = valid ? andOp_199_out : andOp_199_out;
		andOp_203_in1 = valid ? notOp_202_out : notOp_202_out;
	end
	// controller for andOp_205.andOp_205_in0
	// controller for andOp_205.andOp_205_in1
	// Insensitive connections
	always @(*) begin
		andOp_205_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_205_in1 = valid ? notOp_204_out : notOp_204_out;
	end
	// controller for andOp_207.andOp_207_in0
	// controller for andOp_207.andOp_207_in1
	// Insensitive connections
	always @(*) begin
		andOp_207_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_207_in1 = valid ? notOp_206_out : notOp_206_out;
	end
	// controller for andOp_208.andOp_208_in0
	// controller for andOp_208.andOp_208_in1
	// Insensitive connections
	always @(*) begin
		andOp_208_in0 = valid ? 1'd0 : 1'd0;
		andOp_208_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_210.andOp_210_in0
	// controller for andOp_210.andOp_210_in1
	// Insensitive connections
	always @(*) begin
		andOp_210_in0 = valid ? andOp_208_out : andOp_208_out;
		andOp_210_in1 = valid ? eq_209_out : eq_209_out;
	end
	// controller for andOp_212.andOp_212_in0
	// controller for andOp_212.andOp_212_in1
	// Insensitive connections
	always @(*) begin
		andOp_212_in0 = valid ? andOp_208_out : andOp_208_out;
		andOp_212_in1 = valid ? notOp_211_out : notOp_211_out;
	end
	// controller for andOp_214.andOp_214_in0
	// controller for andOp_214.andOp_214_in1
	// Insensitive connections
	always @(*) begin
		andOp_214_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_214_in1 = valid ? notOp_213_out : notOp_213_out;
	end
	// controller for andOp_216.andOp_216_in0
	// controller for andOp_216.andOp_216_in1
	// Insensitive connections
	always @(*) begin
		andOp_216_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_216_in1 = valid ? notOp_215_out : notOp_215_out;
	end
	// controller for andOp_217.andOp_217_in0
	// controller for andOp_217.andOp_217_in1
	// Insensitive connections
	always @(*) begin
		andOp_217_in0 = valid ? 1'd0 : 1'd0;
		andOp_217_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_219.andOp_219_in0
	// controller for andOp_219.andOp_219_in1
	// Insensitive connections
	always @(*) begin
		andOp_219_in0 = valid ? andOp_217_out : andOp_217_out;
		andOp_219_in1 = valid ? eq_218_out : eq_218_out;
	end
	// controller for andOp_221.andOp_221_in0
	// controller for andOp_221.andOp_221_in1
	// Insensitive connections
	always @(*) begin
		andOp_221_in0 = valid ? andOp_217_out : andOp_217_out;
		andOp_221_in1 = valid ? notOp_220_out : notOp_220_out;
	end
	// controller for andOp_223.andOp_223_in0
	// controller for andOp_223.andOp_223_in1
	// Insensitive connections
	always @(*) begin
		andOp_223_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_223_in1 = valid ? notOp_222_out : notOp_222_out;
	end
	// controller for andOp_225.andOp_225_in0
	// controller for andOp_225.andOp_225_in1
	// Insensitive connections
	always @(*) begin
		andOp_225_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_225_in1 = valid ? notOp_224_out : notOp_224_out;
	end
	// controller for andOp_229.andOp_229_in0
	// controller for andOp_229.andOp_229_in1
	// Insensitive connections
	always @(*) begin
		andOp_229_in0 = valid ? 1'd0 : 1'd0;
		andOp_229_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_231.andOp_231_in0
	// controller for andOp_231.andOp_231_in1
	// Insensitive connections
	always @(*) begin
		andOp_231_in0 = valid ? andOp_229_out : andOp_229_out;
		andOp_231_in1 = valid ? eq_230_out : eq_230_out;
	end
	// controller for andOp_233.andOp_233_in0
	// controller for andOp_233.andOp_233_in1
	// Insensitive connections
	always @(*) begin
		andOp_233_in0 = valid ? andOp_229_out : andOp_229_out;
		andOp_233_in1 = valid ? notOp_232_out : notOp_232_out;
	end
	// controller for andOp_235.andOp_235_in0
	// controller for andOp_235.andOp_235_in1
	// Insensitive connections
	always @(*) begin
		andOp_235_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_235_in1 = valid ? notOp_234_out : notOp_234_out;
	end
	// controller for andOp_237.andOp_237_in0
	// controller for andOp_237.andOp_237_in1
	// Insensitive connections
	always @(*) begin
		andOp_237_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_237_in1 = valid ? notOp_236_out : notOp_236_out;
	end
	// controller for andOp_238.andOp_238_in0
	// controller for andOp_238.andOp_238_in1
	// Insensitive connections
	always @(*) begin
		andOp_238_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_238_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_240.andOp_240_in0
	// controller for andOp_240.andOp_240_in1
	// Insensitive connections
	always @(*) begin
		andOp_240_in0 = valid ? andOp_238_out : andOp_238_out;
		andOp_240_in1 = valid ? eq_239_out : eq_239_out;
	end
	// controller for andOp_242.andOp_242_in0
	// controller for andOp_242.andOp_242_in1
	// Insensitive connections
	always @(*) begin
		andOp_242_in0 = valid ? andOp_238_out : andOp_238_out;
		andOp_242_in1 = valid ? notOp_241_out : notOp_241_out;
	end
	// controller for andOp_244.andOp_244_in0
	// controller for andOp_244.andOp_244_in1
	// Insensitive connections
	always @(*) begin
		andOp_244_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_244_in1 = valid ? notOp_243_out : notOp_243_out;
	end
	// controller for andOp_246.andOp_246_in0
	// controller for andOp_246.andOp_246_in1
	// Insensitive connections
	always @(*) begin
		andOp_246_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_246_in1 = valid ? notOp_245_out : notOp_245_out;
	end
	// controller for andOp_247.andOp_247_in0
	// controller for andOp_247.andOp_247_in1
	// Insensitive connections
	always @(*) begin
		andOp_247_in0 = valid ? 1'd0 : 1'd0;
		andOp_247_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_249.andOp_249_in0
	// controller for andOp_249.andOp_249_in1
	// Insensitive connections
	always @(*) begin
		andOp_249_in0 = valid ? andOp_247_out : andOp_247_out;
		andOp_249_in1 = valid ? eq_248_out : eq_248_out;
	end
	// controller for andOp_251.andOp_251_in0
	// controller for andOp_251.andOp_251_in1
	// Insensitive connections
	always @(*) begin
		andOp_251_in0 = valid ? andOp_247_out : andOp_247_out;
		andOp_251_in1 = valid ? notOp_250_out : notOp_250_out;
	end
	// controller for andOp_253.andOp_253_in0
	// controller for andOp_253.andOp_253_in1
	// Insensitive connections
	always @(*) begin
		andOp_253_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_253_in1 = valid ? notOp_252_out : notOp_252_out;
	end
	// controller for andOp_255.andOp_255_in0
	// controller for andOp_255.andOp_255_in1
	// Insensitive connections
	always @(*) begin
		andOp_255_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_255_in1 = valid ? notOp_254_out : notOp_254_out;
	end
	// controller for andOp_256.andOp_256_in0
	// controller for andOp_256.andOp_256_in1
	// Insensitive connections
	always @(*) begin
		andOp_256_in0 = valid ? 1'd0 : 1'd0;
		andOp_256_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_258.andOp_258_in0
	// controller for andOp_258.andOp_258_in1
	// Insensitive connections
	always @(*) begin
		andOp_258_in0 = valid ? andOp_256_out : andOp_256_out;
		andOp_258_in1 = valid ? eq_257_out : eq_257_out;
	end
	// controller for andOp_260.andOp_260_in0
	// controller for andOp_260.andOp_260_in1
	// Insensitive connections
	always @(*) begin
		andOp_260_in0 = valid ? andOp_256_out : andOp_256_out;
		andOp_260_in1 = valid ? notOp_259_out : notOp_259_out;
	end
	// controller for andOp_262.andOp_262_in0
	// controller for andOp_262.andOp_262_in1
	// Insensitive connections
	always @(*) begin
		andOp_262_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_262_in1 = valid ? notOp_261_out : notOp_261_out;
	end
	// controller for andOp_264.andOp_264_in0
	// controller for andOp_264.andOp_264_in1
	// Insensitive connections
	always @(*) begin
		andOp_264_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_264_in1 = valid ? notOp_263_out : notOp_263_out;
	end
	// controller for andOp_267.andOp_267_in0
	// controller for andOp_267.andOp_267_in1
	// Insensitive connections
	always @(*) begin
		andOp_267_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_267_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_269.andOp_269_in0
	// controller for andOp_269.andOp_269_in1
	// Insensitive connections
	always @(*) begin
		andOp_269_in0 = valid ? andOp_267_out : andOp_267_out;
		andOp_269_in1 = valid ? eq_268_out : eq_268_out;
	end
	// controller for andOp_271.andOp_271_in0
	// controller for andOp_271.andOp_271_in1
	// Insensitive connections
	always @(*) begin
		andOp_271_in0 = valid ? andOp_267_out : andOp_267_out;
		andOp_271_in1 = valid ? notOp_270_out : notOp_270_out;
	end
	// controller for andOp_273.andOp_273_in0
	// controller for andOp_273.andOp_273_in1
	// Insensitive connections
	always @(*) begin
		andOp_273_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_273_in1 = valid ? notOp_272_out : notOp_272_out;
	end
	// controller for andOp_275.andOp_275_in0
	// controller for andOp_275.andOp_275_in1
	// Insensitive connections
	always @(*) begin
		andOp_275_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_275_in1 = valid ? notOp_274_out : notOp_274_out;
	end
	// controller for andOp_276.andOp_276_in0
	// controller for andOp_276.andOp_276_in1
	// Insensitive connections
	always @(*) begin
		andOp_276_in0 = valid ? 1'd0 : 1'd0;
		andOp_276_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_278.andOp_278_in0
	// controller for andOp_278.andOp_278_in1
	// Insensitive connections
	always @(*) begin
		andOp_278_in0 = valid ? andOp_276_out : andOp_276_out;
		andOp_278_in1 = valid ? eq_277_out : eq_277_out;
	end
	// controller for andOp_280.andOp_280_in0
	// controller for andOp_280.andOp_280_in1
	// Insensitive connections
	always @(*) begin
		andOp_280_in0 = valid ? andOp_276_out : andOp_276_out;
		andOp_280_in1 = valid ? notOp_279_out : notOp_279_out;
	end
	// controller for andOp_282.andOp_282_in0
	// controller for andOp_282.andOp_282_in1
	// Insensitive connections
	always @(*) begin
		andOp_282_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_282_in1 = valid ? notOp_281_out : notOp_281_out;
	end
	// controller for andOp_284.andOp_284_in0
	// controller for andOp_284.andOp_284_in1
	// Insensitive connections
	always @(*) begin
		andOp_284_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_284_in1 = valid ? notOp_283_out : notOp_283_out;
	end
	// controller for andOp_285.andOp_285_in0
	// controller for andOp_285.andOp_285_in1
	// Insensitive connections
	always @(*) begin
		andOp_285_in0 = valid ? 1'd0 : 1'd0;
		andOp_285_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_287.andOp_287_in0
	// controller for andOp_287.andOp_287_in1
	// Insensitive connections
	always @(*) begin
		andOp_287_in0 = valid ? andOp_285_out : andOp_285_out;
		andOp_287_in1 = valid ? eq_286_out : eq_286_out;
	end
	// controller for andOp_289.andOp_289_in0
	// controller for andOp_289.andOp_289_in1
	// Insensitive connections
	always @(*) begin
		andOp_289_in0 = valid ? andOp_285_out : andOp_285_out;
		andOp_289_in1 = valid ? notOp_288_out : notOp_288_out;
	end
	// controller for andOp_291.andOp_291_in0
	// controller for andOp_291.andOp_291_in1
	// Insensitive connections
	always @(*) begin
		andOp_291_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_291_in1 = valid ? notOp_290_out : notOp_290_out;
	end
	// controller for andOp_293.andOp_293_in0
	// controller for andOp_293.andOp_293_in1
	// Insensitive connections
	always @(*) begin
		andOp_293_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_293_in1 = valid ? notOp_292_out : notOp_292_out;
	end
	// controller for andOp_294.andOp_294_in0
	// controller for andOp_294.andOp_294_in1
	// Insensitive connections
	always @(*) begin
		andOp_294_in0 = valid ? 1'd0 : 1'd0;
		andOp_294_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_296.andOp_296_in0
	// controller for andOp_296.andOp_296_in1
	// Insensitive connections
	always @(*) begin
		andOp_296_in0 = valid ? andOp_294_out : andOp_294_out;
		andOp_296_in1 = valid ? eq_295_out : eq_295_out;
	end
	// controller for andOp_298.andOp_298_in0
	// controller for andOp_298.andOp_298_in1
	// Insensitive connections
	always @(*) begin
		andOp_298_in0 = valid ? andOp_294_out : andOp_294_out;
		andOp_298_in1 = valid ? notOp_297_out : notOp_297_out;
	end
	// controller for andOp_300.andOp_300_in0
	// controller for andOp_300.andOp_300_in1
	// Insensitive connections
	always @(*) begin
		andOp_300_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_300_in1 = valid ? notOp_299_out : notOp_299_out;
	end
	// controller for andOp_302.andOp_302_in0
	// controller for andOp_302.andOp_302_in1
	// Insensitive connections
	always @(*) begin
		andOp_302_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_302_in1 = valid ? notOp_301_out : notOp_301_out;
	end
	// controller for andOp_305.andOp_305_in0
	// controller for andOp_305.andOp_305_in1
	// Insensitive connections
	always @(*) begin
		andOp_305_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_305_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_307.andOp_307_in0
	// controller for andOp_307.andOp_307_in1
	// Insensitive connections
	always @(*) begin
		andOp_307_in0 = valid ? andOp_305_out : andOp_305_out;
		andOp_307_in1 = valid ? eq_306_out : eq_306_out;
	end
	// controller for andOp_309.andOp_309_in0
	// controller for andOp_309.andOp_309_in1
	// Insensitive connections
	always @(*) begin
		andOp_309_in0 = valid ? andOp_305_out : andOp_305_out;
		andOp_309_in1 = valid ? notOp_308_out : notOp_308_out;
	end
	// controller for andOp_311.andOp_311_in0
	// controller for andOp_311.andOp_311_in1
	// Insensitive connections
	always @(*) begin
		andOp_311_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_311_in1 = valid ? notOp_310_out : notOp_310_out;
	end
	// controller for andOp_313.andOp_313_in0
	// controller for andOp_313.andOp_313_in1
	// Insensitive connections
	always @(*) begin
		andOp_313_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_313_in1 = valid ? notOp_312_out : notOp_312_out;
	end
	// controller for andOp_314.andOp_314_in0
	// controller for andOp_314.andOp_314_in1
	// Insensitive connections
	always @(*) begin
		andOp_314_in0 = valid ? 1'd0 : 1'd0;
		andOp_314_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_316.andOp_316_in0
	// controller for andOp_316.andOp_316_in1
	// Insensitive connections
	always @(*) begin
		andOp_316_in0 = valid ? andOp_314_out : andOp_314_out;
		andOp_316_in1 = valid ? eq_315_out : eq_315_out;
	end
	// controller for andOp_318.andOp_318_in0
	// controller for andOp_318.andOp_318_in1
	// Insensitive connections
	always @(*) begin
		andOp_318_in0 = valid ? andOp_314_out : andOp_314_out;
		andOp_318_in1 = valid ? notOp_317_out : notOp_317_out;
	end
	// controller for andOp_320.andOp_320_in0
	// controller for andOp_320.andOp_320_in1
	// Insensitive connections
	always @(*) begin
		andOp_320_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_320_in1 = valid ? notOp_319_out : notOp_319_out;
	end
	// controller for andOp_322.andOp_322_in0
	// controller for andOp_322.andOp_322_in1
	// Insensitive connections
	always @(*) begin
		andOp_322_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_322_in1 = valid ? notOp_321_out : notOp_321_out;
	end
	// controller for andOp_323.andOp_323_in0
	// controller for andOp_323.andOp_323_in1
	// Insensitive connections
	always @(*) begin
		andOp_323_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_323_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_325.andOp_325_in0
	// controller for andOp_325.andOp_325_in1
	// Insensitive connections
	always @(*) begin
		andOp_325_in0 = valid ? andOp_323_out : andOp_323_out;
		andOp_325_in1 = valid ? eq_324_out : eq_324_out;
	end
	// controller for andOp_327.andOp_327_in0
	// controller for andOp_327.andOp_327_in1
	// Insensitive connections
	always @(*) begin
		andOp_327_in0 = valid ? andOp_323_out : andOp_323_out;
		andOp_327_in1 = valid ? notOp_326_out : notOp_326_out;
	end
	// controller for andOp_329.andOp_329_in0
	// controller for andOp_329.andOp_329_in1
	// Insensitive connections
	always @(*) begin
		andOp_329_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_329_in1 = valid ? notOp_328_out : notOp_328_out;
	end
	// controller for andOp_331.andOp_331_in0
	// controller for andOp_331.andOp_331_in1
	// Insensitive connections
	always @(*) begin
		andOp_331_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_331_in1 = valid ? notOp_330_out : notOp_330_out;
	end
	// controller for andOp_332.andOp_332_in0
	// controller for andOp_332.andOp_332_in1
	// Insensitive connections
	always @(*) begin
		andOp_332_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_332_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_334.andOp_334_in0
	// controller for andOp_334.andOp_334_in1
	// Insensitive connections
	always @(*) begin
		andOp_334_in0 = valid ? andOp_332_out : andOp_332_out;
		andOp_334_in1 = valid ? eq_333_out : eq_333_out;
	end
	// controller for andOp_336.andOp_336_in0
	// controller for andOp_336.andOp_336_in1
	// Insensitive connections
	always @(*) begin
		andOp_336_in0 = valid ? andOp_332_out : andOp_332_out;
		andOp_336_in1 = valid ? notOp_335_out : notOp_335_out;
	end
	// controller for andOp_338.andOp_338_in0
	// controller for andOp_338.andOp_338_in1
	// Insensitive connections
	always @(*) begin
		andOp_338_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_338_in1 = valid ? notOp_337_out : notOp_337_out;
	end
	// controller for andOp_340.andOp_340_in0
	// controller for andOp_340.andOp_340_in1
	// Insensitive connections
	always @(*) begin
		andOp_340_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_340_in1 = valid ? notOp_339_out : notOp_339_out;
	end
	// controller for andOp_343.andOp_343_in0
	// controller for andOp_343.andOp_343_in1
	// Insensitive connections
	always @(*) begin
		andOp_343_in0 = valid ? 1'd0 : 1'd0;
		andOp_343_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_345.andOp_345_in0
	// controller for andOp_345.andOp_345_in1
	// Insensitive connections
	always @(*) begin
		andOp_345_in0 = valid ? andOp_343_out : andOp_343_out;
		andOp_345_in1 = valid ? eq_344_out : eq_344_out;
	end
	// controller for andOp_347.andOp_347_in0
	// controller for andOp_347.andOp_347_in1
	// Insensitive connections
	always @(*) begin
		andOp_347_in0 = valid ? andOp_343_out : andOp_343_out;
		andOp_347_in1 = valid ? notOp_346_out : notOp_346_out;
	end
	// controller for andOp_349.andOp_349_in0
	// controller for andOp_349.andOp_349_in1
	// Insensitive connections
	always @(*) begin
		andOp_349_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_349_in1 = valid ? notOp_348_out : notOp_348_out;
	end
	// controller for andOp_351.andOp_351_in0
	// controller for andOp_351.andOp_351_in1
	// Insensitive connections
	always @(*) begin
		andOp_351_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_351_in1 = valid ? notOp_350_out : notOp_350_out;
	end
	// controller for andOp_352.andOp_352_in0
	// controller for andOp_352.andOp_352_in1
	// Insensitive connections
	always @(*) begin
		andOp_352_in0 = valid ? 1'd0 : 1'd0;
		andOp_352_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_354.andOp_354_in0
	// controller for andOp_354.andOp_354_in1
	// Insensitive connections
	always @(*) begin
		andOp_354_in0 = valid ? andOp_352_out : andOp_352_out;
		andOp_354_in1 = valid ? eq_353_out : eq_353_out;
	end
	// controller for andOp_356.andOp_356_in0
	// controller for andOp_356.andOp_356_in1
	// Insensitive connections
	always @(*) begin
		andOp_356_in0 = valid ? andOp_352_out : andOp_352_out;
		andOp_356_in1 = valid ? notOp_355_out : notOp_355_out;
	end
	// controller for andOp_358.andOp_358_in0
	// controller for andOp_358.andOp_358_in1
	// Insensitive connections
	always @(*) begin
		andOp_358_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_358_in1 = valid ? notOp_357_out : notOp_357_out;
	end
	// controller for andOp_360.andOp_360_in0
	// controller for andOp_360.andOp_360_in1
	// Insensitive connections
	always @(*) begin
		andOp_360_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_360_in1 = valid ? notOp_359_out : notOp_359_out;
	end
	// controller for andOp_361.andOp_361_in0
	// controller for andOp_361.andOp_361_in1
	// Insensitive connections
	always @(*) begin
		andOp_361_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_361_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_363.andOp_363_in0
	// controller for andOp_363.andOp_363_in1
	// Insensitive connections
	always @(*) begin
		andOp_363_in0 = valid ? andOp_361_out : andOp_361_out;
		andOp_363_in1 = valid ? eq_362_out : eq_362_out;
	end
	// controller for andOp_365.andOp_365_in0
	// controller for andOp_365.andOp_365_in1
	// Insensitive connections
	always @(*) begin
		andOp_365_in0 = valid ? andOp_361_out : andOp_361_out;
		andOp_365_in1 = valid ? notOp_364_out : notOp_364_out;
	end
	// controller for andOp_367.andOp_367_in0
	// controller for andOp_367.andOp_367_in1
	// Insensitive connections
	always @(*) begin
		andOp_367_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_367_in1 = valid ? notOp_366_out : notOp_366_out;
	end
	// controller for andOp_369.andOp_369_in0
	// controller for andOp_369.andOp_369_in1
	// Insensitive connections
	always @(*) begin
		andOp_369_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_369_in1 = valid ? notOp_368_out : notOp_368_out;
	end
	// controller for andOp_370.andOp_370_in0
	// controller for andOp_370.andOp_370_in1
	// Insensitive connections
	always @(*) begin
		andOp_370_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_370_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_372.andOp_372_in0
	// controller for andOp_372.andOp_372_in1
	// Insensitive connections
	always @(*) begin
		andOp_372_in0 = valid ? andOp_370_out : andOp_370_out;
		andOp_372_in1 = valid ? eq_371_out : eq_371_out;
	end
	// controller for andOp_374.andOp_374_in0
	// controller for andOp_374.andOp_374_in1
	// Insensitive connections
	always @(*) begin
		andOp_374_in0 = valid ? andOp_370_out : andOp_370_out;
		andOp_374_in1 = valid ? notOp_373_out : notOp_373_out;
	end
	// controller for andOp_376.andOp_376_in0
	// controller for andOp_376.andOp_376_in1
	// Insensitive connections
	always @(*) begin
		andOp_376_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_376_in1 = valid ? notOp_375_out : notOp_375_out;
	end
	// controller for andOp_378.andOp_378_in0
	// controller for andOp_378.andOp_378_in1
	// Insensitive connections
	always @(*) begin
		andOp_378_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_378_in1 = valid ? notOp_377_out : notOp_377_out;
	end
	// controller for andOp_40.andOp_40_in0
	// controller for andOp_40.andOp_40_in1
	// Insensitive connections
	always @(*) begin
		andOp_40_in0 = valid ? bb_0_active_in_state_1_out_data : bb_0_active_in_state_1_out_data;
		andOp_40_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_41.andOp_41_in0
	// controller for andOp_41.andOp_41_in1
	// Insensitive connections
	always @(*) begin
		andOp_41_in0 = valid ? andOp_40_out : andOp_40_out;
		andOp_41_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_43.andOp_43_in0
	// controller for andOp_43.andOp_43_in1
	// Insensitive connections
	always @(*) begin
		andOp_43_in0 = valid ? bb_8_active_in_state_1_out_data : bb_8_active_in_state_1_out_data;
		andOp_43_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_44.andOp_44_in0
	// controller for andOp_44.andOp_44_in1
	// Insensitive connections
	always @(*) begin
		andOp_44_in0 = valid ? andOp_43_out : andOp_43_out;
		andOp_44_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_46.andOp_46_in0
	// controller for andOp_46.andOp_46_in1
	// Insensitive connections
	always @(*) begin
		andOp_46_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
		andOp_46_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_47.andOp_47_in0
	// controller for andOp_47.andOp_47_in1
	// Insensitive connections
	always @(*) begin
		andOp_47_in0 = valid ? andOp_46_out : andOp_46_out;
		andOp_47_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_49.andOp_49_in0
	// controller for andOp_49.andOp_49_in1
	// Insensitive connections
	always @(*) begin
		andOp_49_in0 = valid ? andOp_47_out : andOp_47_out;
		andOp_49_in1 = valid ? in_read_ready : in_read_ready;
	end
	// controller for andOp_51.andOp_51_in0
	// controller for andOp_51.andOp_51_in1
	// Insensitive connections
	always @(*) begin
		andOp_51_in0 = valid ? andOp_47_out : andOp_47_out;
		andOp_51_in1 = valid ? notOp_50_out : notOp_50_out;
	end
	// controller for andOp_52.andOp_52_in0
	// controller for andOp_52.andOp_52_in1
	// Insensitive connections
	always @(*) begin
		andOp_52_in0 = valid ? bb_0_active_in_state_1_out_data : bb_0_active_in_state_1_out_data;
		andOp_52_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_53.andOp_53_in0
	// controller for andOp_53.andOp_53_in1
	// Insensitive connections
	always @(*) begin
		andOp_53_in0 = valid ? andOp_52_out : andOp_52_out;
		andOp_53_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_55.andOp_55_in0
	// controller for andOp_55.andOp_55_in1
	// Insensitive connections
	always @(*) begin
		andOp_55_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_55_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_56.andOp_56_in0
	// controller for andOp_56.andOp_56_in1
	// Insensitive connections
	always @(*) begin
		andOp_56_in0 = valid ? andOp_55_out : andOp_55_out;
		andOp_56_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_58.andOp_58_in0
	// controller for andOp_58.andOp_58_in1
	// Insensitive connections
	always @(*) begin
		andOp_58_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_58_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_59.andOp_59_in0
	// controller for andOp_59.andOp_59_in1
	// Insensitive connections
	always @(*) begin
		andOp_59_in0 = valid ? andOp_58_out : andOp_58_out;
		andOp_59_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_61.andOp_61_in0
	// controller for andOp_61.andOp_61_in1
	// Insensitive connections
	always @(*) begin
		andOp_61_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_61_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_62.andOp_62_in0
	// controller for andOp_62.andOp_62_in1
	// Insensitive connections
	always @(*) begin
		andOp_62_in0 = valid ? andOp_61_out : andOp_61_out;
		andOp_62_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_64.andOp_64_in0
	// controller for andOp_64.andOp_64_in1
	// Insensitive connections
	always @(*) begin
		andOp_64_in0 = valid ? andOp_62_out : andOp_62_out;
		andOp_64_in1 = valid ? data_in_4_39_out_data : data_in_4_39_out_data;
	end
	// controller for andOp_66.andOp_66_in0
	// controller for andOp_66.andOp_66_in1
	// Insensitive connections
	always @(*) begin
		andOp_66_in0 = valid ? andOp_62_out : andOp_62_out;
		andOp_66_in1 = valid ? notOp_65_out : notOp_65_out;
	end
	// controller for andOp_67.andOp_67_in0
	// controller for andOp_67.andOp_67_in1
	// Insensitive connections
	always @(*) begin
		andOp_67_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_67_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_68.andOp_68_in0
	// controller for andOp_68.andOp_68_in1
	// Insensitive connections
	always @(*) begin
		andOp_68_in0 = valid ? andOp_67_out : andOp_67_out;
		andOp_68_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_70.andOp_70_in0
	// controller for andOp_70.andOp_70_in1
	// Insensitive connections
	always @(*) begin
		andOp_70_in0 = valid ? bb_5_active_in_state_4_out_data : bb_5_active_in_state_4_out_data;
		andOp_70_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_71.andOp_71_in0
	// controller for andOp_71.andOp_71_in1
	// Insensitive connections
	always @(*) begin
		andOp_71_in0 = valid ? andOp_70_out : andOp_70_out;
		andOp_71_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_73.andOp_73_in0
	// controller for andOp_73.andOp_73_in1
	// Insensitive connections
	always @(*) begin
		andOp_73_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_73_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_74.andOp_74_in0
	// controller for andOp_74.andOp_74_in1
	// Insensitive connections
	always @(*) begin
		andOp_74_in0 = valid ? andOp_73_out : andOp_73_out;
		andOp_74_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_76.andOp_76_in0
	// controller for andOp_76.andOp_76_in1
	// Insensitive connections
	always @(*) begin
		andOp_76_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
		andOp_76_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_77.andOp_77_in0
	// controller for andOp_77.andOp_77_in1
	// Insensitive connections
	always @(*) begin
		andOp_77_in0 = valid ? andOp_76_out : andOp_76_out;
		andOp_77_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_79.andOp_79_in0
	// controller for andOp_79.andOp_79_in1
	// Insensitive connections
	always @(*) begin
		andOp_79_in0 = valid ? andOp_77_out : andOp_77_out;
		andOp_79_in1 = valid ? out_write_ready : out_write_ready;
	end
	// controller for andOp_81.andOp_81_in0
	// controller for andOp_81.andOp_81_in1
	// Insensitive connections
	always @(*) begin
		andOp_81_in0 = valid ? andOp_77_out : andOp_77_out;
		andOp_81_in1 = valid ? notOp_80_out : notOp_80_out;
	end
	// controller for andOp_82.andOp_82_in0
	// controller for andOp_82.andOp_82_in1
	// Insensitive connections
	always @(*) begin
		andOp_82_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_82_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_83.andOp_83_in0
	// controller for andOp_83.andOp_83_in1
	// Insensitive connections
	always @(*) begin
		andOp_83_in0 = valid ? andOp_82_out : andOp_82_out;
		andOp_83_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_85.andOp_85_in0
	// controller for andOp_85.andOp_85_in1
	// Insensitive connections
	always @(*) begin
		andOp_85_in0 = valid ? andOp_83_out : andOp_83_out;
		andOp_85_in1 = valid ? data_in_4_39_out_data : data_in_4_39_out_data;
	end
	// controller for andOp_87.andOp_87_in0
	// controller for andOp_87.andOp_87_in1
	// Insensitive connections
	always @(*) begin
		andOp_87_in0 = valid ? andOp_83_out : andOp_83_out;
		andOp_87_in1 = valid ? notOp_86_out : notOp_86_out;
	end
	// controller for andOp_88.andOp_88_in0
	// controller for andOp_88.andOp_88_in1
	// Insensitive connections
	always @(*) begin
		andOp_88_in0 = valid ? bb_1_active_in_state_4_out_data : bb_1_active_in_state_4_out_data;
		andOp_88_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_89.andOp_89_in0
	// controller for andOp_89.andOp_89_in1
	// Insensitive connections
	always @(*) begin
		andOp_89_in0 = valid ? andOp_88_out : andOp_88_out;
		andOp_89_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_91_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_active_in_state_1.bb_0_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_1_in_data = eq_96_out;
		end else begin
			bb_0_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_114_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_1.bb_0_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_121_out) begin 
			bb_0_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_2.bb_10_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_2_in_data = eq_99_out;
		end else begin
			bb_10_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_3.bb_10_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_3_in_data = eq_102_out;
		end else begin
			bb_10_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_2.bb_10_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_125_out) begin 
			bb_10_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_3.bb_10_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_129_out) begin 
			bb_10_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_4.bb_1_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_4_in_data = orOp_113_out;
		end else begin
			bb_1_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_4.bb_1_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_145_out) begin 
			bb_1_predecessor_in_state_4_in_data = 32'd4;
		end else if (eq_143_out) begin 
			bb_1_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_4.bb_2_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_4_in_data = orOp_104_out;
		end else begin
			bb_2_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_4.bb_2_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_132_out) begin 
			bb_2_predecessor_in_state_4_in_data = 32'd7;
		end else if (eq_130_out) begin 
			bb_2_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_1.bb_3_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_1_in_data = orOp_98_out;
		end else begin
			bb_3_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_1.bb_3_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_124_out) begin 
			bb_3_predecessor_in_state_1_in_data = 32'd0;
		end else if (eq_122_out) begin 
			bb_3_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_3.bb_4_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_3_in_data = orOp_101_out;
		end else begin
			bb_4_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_4.bb_4_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_4_in_data = eq_111_out;
		end else begin
			bb_4_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_3.bb_4_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_128_out) begin 
			bb_4_predecessor_in_state_3_in_data = 32'd10;
		end else if (eq_126_out) begin 
			bb_4_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_4.bb_4_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_142_out) begin 
			bb_4_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_5_active_in_state_4.bb_5_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_5_active_in_state_4_in_data = orOp_106_out;
		end else begin
			bb_5_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_5_predecessor_in_state_4.bb_5_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_135_out) begin 
			bb_5_predecessor_in_state_4_in_data = 32'd1;
		end else if (eq_133_out) begin 
			bb_5_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_5_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_6_active_in_state_4.bb_6_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_6_active_in_state_4_in_data = orOp_110_out;
		end else begin
			bb_6_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_6_predecessor_in_state_4.bb_6_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_141_out) begin 
			bb_6_predecessor_in_state_4_in_data = 32'd5;
		end else if (eq_139_out) begin 
			bb_6_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_6_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_7_active_in_state_4.bb_7_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_7_active_in_state_4_in_data = orOp_108_out;
		end else begin
			bb_7_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_7_predecessor_in_state_4.bb_7_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_138_out) begin 
			bb_7_predecessor_in_state_4_in_data = 32'd6;
		end else if (eq_136_out) begin 
			bb_7_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_7_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_8_active_in_state_1.bb_8_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_state_1_in_data = orOp_93_out;
		end else begin
			bb_8_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_8_predecessor_in_state_1.bb_8_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_117_out) begin 
			bb_8_predecessor_in_state_1_in_data = 32'd3;
		end else if (eq_115_out) begin 
			bb_8_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_8_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_9_active_in_state_1.bb_9_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_9_active_in_state_1_in_data = orOp_95_out;
		end else begin
			bb_9_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_9_predecessor_in_state_1.bb_9_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_120_out) begin 
			bb_9_predecessor_in_state_1_in_data = 32'd8;
		end else if (eq_118_out) begin 
			bb_9_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_9_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_41_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_42_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_1.br_0_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_53_out) begin 
			br_0_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_54_out) begin 
			br_0_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_2.br_10_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_59_out) begin 
			br_10_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_60_out) begin 
			br_10_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_3.br_10_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_68_out) begin 
			br_10_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_69_out) begin 
			br_10_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_1_happened_in_state_4.br_1_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_89_out) begin 
			br_1_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_90_out) begin 
			br_1_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_1_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_1.br_3_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_56_out) begin 
			br_3_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_57_out) begin 
			br_3_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_3.br_4_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_62_out) begin 
			br_4_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_63_out) begin 
			br_4_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_4.br_4_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_83_out) begin 
			br_4_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_84_out) begin 
			br_4_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_5_happened_in_state_4.br_5_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_71_out) begin 
			br_5_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_72_out) begin 
			br_5_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_5_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_6_happened_in_state_4.br_6_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_77_out) begin 
			br_6_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_78_out) begin 
			br_6_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_6_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_7_happened_in_state_4.br_7_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_74_out) begin 
			br_7_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_75_out) begin 
			br_7_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_7_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_8_happened_in_state_1.br_8_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_44_out) begin 
			br_8_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_45_out) begin 
			br_8_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_8_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_9_happened_in_state_1.br_9_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_47_out) begin 
			br_9_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_48_out) begin 
			br_9_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_9_happened_in_state_1_in_data = 0;
		end
	end
	// controller for concat_157.concat_157_in0
	// controller for concat_157.concat_157_in1
	// Insensitive connections
	always @(*) begin
		concat_157_in0 = valid ? data_in_1_13_out_data : data_in_1_13_out_data;
		concat_157_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for concat_158.concat_158_in0
	// controller for concat_158.concat_158_in1
	// Insensitive connections
	always @(*) begin
		concat_158_in0 = valid ? 32'd4 : 32'd4;
		concat_158_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for data_in_0_1.data_in_0_1_in_data
	always @(*) begin
		if (eq_189_out) begin 
			data_in_0_1_in_data = data_store_0_0;
		end else begin
			data_in_0_1_in_data = 0;
		end
	end
	// controller for data_in_0_3.data_in_0_3_in_data
	always @(*) begin
		if (eq_189_out) begin 
			data_in_0_3_in_data = data_store_0_2;
		end else begin
			data_in_0_3_in_data = 0;
		end
	end
	// controller for data_in_0_5.data_in_0_5_in_data
	always @(*) begin
		if (eq_189_out) begin 
			data_in_0_5_in_data = data_store_0_4;
		end else begin
			data_in_0_5_in_data = 0;
		end
	end
	// controller for data_in_0_7.data_in_0_7_in_data
	always @(*) begin
		if (eq_189_out) begin 
			data_in_0_7_in_data = data_store_0_6;
		end else begin
			data_in_0_7_in_data = 0;
		end
	end
	// controller for data_in_1_11.data_in_1_11_in_data
	always @(*) begin
		if (eq_226_out) begin 
			data_in_1_11_in_data = data_store_0_2;
		end else if (eq_227_out) begin 
			data_in_1_11_in_data = data_store_1_10;
		end else if (eq_228_out) begin 
			data_in_1_11_in_data = data_store_4_34;
		end else begin
			data_in_1_11_in_data = 0;
		end
	end
	// controller for data_in_1_13.data_in_1_13_in_data
	always @(*) begin
		if (eq_226_out) begin 
			data_in_1_13_in_data = data_store_0_4;
		end else if (eq_227_out) begin 
			data_in_1_13_in_data = data_store_1_12;
		end else if (eq_228_out) begin 
			data_in_1_13_in_data = data_store_4_36;
		end else begin
			data_in_1_13_in_data = 0;
		end
	end
	// controller for data_in_1_15.data_in_1_15_in_data
	always @(*) begin
		if (eq_226_out) begin 
			data_in_1_15_in_data = data_store_0_6;
		end else if (eq_227_out) begin 
			data_in_1_15_in_data = data_store_1_14;
		end else if (eq_228_out) begin 
			data_in_1_15_in_data = data_store_4_38;
		end else begin
			data_in_1_15_in_data = 0;
		end
	end
	// controller for data_in_1_9.data_in_1_9_in_data
	always @(*) begin
		if (eq_226_out) begin 
			data_in_1_9_in_data = data_store_0_0;
		end else if (eq_227_out) begin 
			data_in_1_9_in_data = data_store_1_8;
		end else if (eq_228_out) begin 
			data_in_1_9_in_data = data_store_4_32;
		end else begin
			data_in_1_9_in_data = 0;
		end
	end
	// controller for data_in_2_17.data_in_2_17_in_data
	always @(*) begin
		if (eq_265_out) begin 
			data_in_2_17_in_data = data_store_1_8;
		end else if (eq_266_out) begin 
			data_in_2_17_in_data = data_store_2_16;
		end else begin
			data_in_2_17_in_data = 0;
		end
	end
	// controller for data_in_2_19.data_in_2_19_in_data
	always @(*) begin
		if (eq_265_out) begin 
			data_in_2_19_in_data = data_store_1_10;
		end else if (eq_266_out) begin 
			data_in_2_19_in_data = data_store_2_18;
		end else begin
			data_in_2_19_in_data = 0;
		end
	end
	// controller for data_in_2_21.data_in_2_21_in_data
	always @(*) begin
		if (eq_265_out) begin 
			data_in_2_21_in_data = data_store_1_12;
		end else if (eq_266_out) begin 
			data_in_2_21_in_data = data_store_2_20;
		end else begin
			data_in_2_21_in_data = 0;
		end
	end
	// controller for data_in_2_23.data_in_2_23_in_data
	always @(*) begin
		if (eq_265_out) begin 
			data_in_2_23_in_data = data_store_1_14;
		end else if (eq_266_out) begin 
			data_in_2_23_in_data = data_store_2_22;
		end else begin
			data_in_2_23_in_data = 0;
		end
	end
	// controller for data_in_3_25.data_in_3_25_in_data
	always @(*) begin
		if (eq_303_out) begin 
			data_in_3_25_in_data = data_store_2_16;
		end else if (eq_304_out) begin 
			data_in_3_25_in_data = data_store_3_24;
		end else begin
			data_in_3_25_in_data = 0;
		end
	end
	// controller for data_in_3_27.data_in_3_27_in_data
	always @(*) begin
		if (eq_303_out) begin 
			data_in_3_27_in_data = data_store_2_18;
		end else if (eq_304_out) begin 
			data_in_3_27_in_data = data_store_3_26;
		end else begin
			data_in_3_27_in_data = 0;
		end
	end
	// controller for data_in_3_29.data_in_3_29_in_data
	always @(*) begin
		if (eq_303_out) begin 
			data_in_3_29_in_data = data_store_2_20;
		end else if (eq_304_out) begin 
			data_in_3_29_in_data = data_store_3_28;
		end else begin
			data_in_3_29_in_data = 0;
		end
	end
	// controller for data_in_3_31.data_in_3_31_in_data
	always @(*) begin
		if (eq_303_out) begin 
			data_in_3_31_in_data = data_store_2_22;
		end else if (eq_304_out) begin 
			data_in_3_31_in_data = data_store_3_30;
		end else begin
			data_in_3_31_in_data = 0;
		end
	end
	// controller for data_in_4_33.data_in_4_33_in_data
	always @(*) begin
		if (eq_341_out) begin 
			data_in_4_33_in_data = data_store_3_24;
		end else if (eq_342_out) begin 
			data_in_4_33_in_data = data_store_4_32;
		end else begin
			data_in_4_33_in_data = 0;
		end
	end
	// controller for data_in_4_35.data_in_4_35_in_data
	always @(*) begin
		if (eq_341_out) begin 
			data_in_4_35_in_data = data_store_3_26;
		end else if (eq_342_out) begin 
			data_in_4_35_in_data = data_store_4_34;
		end else begin
			data_in_4_35_in_data = 0;
		end
	end
	// controller for data_in_4_37.data_in_4_37_in_data
	always @(*) begin
		if (eq_341_out) begin 
			data_in_4_37_in_data = data_store_3_28;
		end else if (eq_342_out) begin 
			data_in_4_37_in_data = data_store_4_36;
		end else begin
			data_in_4_37_in_data = 0;
		end
	end
	// controller for data_in_4_39.data_in_4_39_in_data
	always @(*) begin
		if (eq_341_out) begin 
			data_in_4_39_in_data = data_store_3_30;
		end else if (eq_342_out) begin 
			data_in_4_39_in_data = data_store_4_38;
		end else begin
			data_in_4_39_in_data = 0;
		end
	end
	// controller for eq_100.eq_100_in0
	// controller for eq_100.eq_100_in1
	// Insensitive connections
	always @(*) begin
		eq_100_in0 = valid ? 32'd4 : 32'd4;
		eq_100_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_102.eq_102_in0
	// controller for eq_102.eq_102_in1
	// Insensitive connections
	always @(*) begin
		eq_102_in0 = valid ? 32'd10 : 32'd10;
		eq_102_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_103.eq_103_in0
	// controller for eq_103.eq_103_in1
	// Insensitive connections
	always @(*) begin
		eq_103_in0 = valid ? 32'd2 : 32'd2;
		eq_103_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_105.eq_105_in0
	// controller for eq_105.eq_105_in1
	// Insensitive connections
	always @(*) begin
		eq_105_in0 = valid ? 32'd5 : 32'd5;
		eq_105_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_107.eq_107_in0
	// controller for eq_107.eq_107_in1
	// Insensitive connections
	always @(*) begin
		eq_107_in0 = valid ? 32'd7 : 32'd7;
		eq_107_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_109.eq_109_in0
	// controller for eq_109.eq_109_in1
	// Insensitive connections
	always @(*) begin
		eq_109_in0 = valid ? 32'd6 : 32'd6;
		eq_109_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_111.eq_111_in0
	// controller for eq_111.eq_111_in1
	// Insensitive connections
	always @(*) begin
		eq_111_in0 = valid ? 32'd4 : 32'd4;
		eq_111_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_112.eq_112_in0
	// controller for eq_112.eq_112_in1
	// Insensitive connections
	always @(*) begin
		eq_112_in0 = valid ? 32'd1 : 32'd1;
		eq_112_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_114.eq_114_in0
	// controller for eq_114.eq_114_in1
	// Insensitive connections
	always @(*) begin
		eq_114_in0 = valid ? 32'd0 : 32'd0;
		eq_114_in1 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
	end
	// controller for eq_115.eq_115_in0
	// controller for eq_115.eq_115_in1
	// Insensitive connections
	always @(*) begin
		eq_115_in0 = valid ? 32'd8 : 32'd8;
		eq_115_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_118.eq_118_in0
	// controller for eq_118.eq_118_in1
	// Insensitive connections
	always @(*) begin
		eq_118_in0 = valid ? 32'd9 : 32'd9;
		eq_118_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_121.eq_121_in0
	// controller for eq_121.eq_121_in1
	// Insensitive connections
	always @(*) begin
		eq_121_in0 = valid ? 32'd0 : 32'd0;
		eq_121_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_122.eq_122_in0
	// controller for eq_122.eq_122_in1
	// Insensitive connections
	always @(*) begin
		eq_122_in0 = valid ? 32'd3 : 32'd3;
		eq_122_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_125.eq_125_in0
	// controller for eq_125.eq_125_in1
	// Insensitive connections
	always @(*) begin
		eq_125_in0 = valid ? 32'd10 : 32'd10;
		eq_125_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_126.eq_126_in0
	// controller for eq_126.eq_126_in1
	// Insensitive connections
	always @(*) begin
		eq_126_in0 = valid ? 32'd4 : 32'd4;
		eq_126_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_129.eq_129_in0
	// controller for eq_129.eq_129_in1
	// Insensitive connections
	always @(*) begin
		eq_129_in0 = valid ? 32'd10 : 32'd10;
		eq_129_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_130.eq_130_in0
	// controller for eq_130.eq_130_in1
	// Insensitive connections
	always @(*) begin
		eq_130_in0 = valid ? 32'd2 : 32'd2;
		eq_130_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_133.eq_133_in0
	// controller for eq_133.eq_133_in1
	// Insensitive connections
	always @(*) begin
		eq_133_in0 = valid ? 32'd5 : 32'd5;
		eq_133_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_136.eq_136_in0
	// controller for eq_136.eq_136_in1
	// Insensitive connections
	always @(*) begin
		eq_136_in0 = valid ? 32'd7 : 32'd7;
		eq_136_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_139.eq_139_in0
	// controller for eq_139.eq_139_in1
	// Insensitive connections
	always @(*) begin
		eq_139_in0 = valid ? 32'd6 : 32'd6;
		eq_139_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_142.eq_142_in0
	// controller for eq_142.eq_142_in1
	// Insensitive connections
	always @(*) begin
		eq_142_in0 = valid ? 32'd4 : 32'd4;
		eq_142_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_143.eq_143_in0
	// controller for eq_143.eq_143_in1
	// Insensitive connections
	always @(*) begin
		eq_143_in0 = valid ? 32'd1 : 32'd1;
		eq_143_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_161.eq_161_in0
	// controller for eq_161.eq_161_in1
	// Insensitive connections
	always @(*) begin
		eq_161_in0 = valid ? 32'd10 : 32'd10;
		eq_161_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_189.eq_189_in0
	// controller for eq_189.eq_189_in1
	// Insensitive connections
	always @(*) begin
		eq_189_in0 = valid ? 32'd0 : 32'd0;
		eq_189_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_191.eq_191_in0
	// controller for eq_191.eq_191_in1
	// Insensitive connections
	always @(*) begin
		eq_191_in0 = valid ? 32'd3 : 32'd3;
		eq_191_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_200.eq_200_in0
	// controller for eq_200.eq_200_in1
	// Insensitive connections
	always @(*) begin
		eq_200_in0 = valid ? 32'd1 : 32'd1;
		eq_200_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_209.eq_209_in0
	// controller for eq_209.eq_209_in1
	// Insensitive connections
	always @(*) begin
		eq_209_in0 = valid ? 32'd3 : 32'd3;
		eq_209_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_218.eq_218_in0
	// controller for eq_218.eq_218_in1
	// Insensitive connections
	always @(*) begin
		eq_218_in0 = valid ? 32'd3 : 32'd3;
		eq_218_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_226.eq_226_in0
	// controller for eq_226.eq_226_in1
	// Insensitive connections
	always @(*) begin
		eq_226_in0 = valid ? 32'd0 : 32'd0;
		eq_226_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_227.eq_227_in0
	// controller for eq_227.eq_227_in1
	// Insensitive connections
	always @(*) begin
		eq_227_in0 = valid ? 32'd1 : 32'd1;
		eq_227_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_228.eq_228_in0
	// controller for eq_228.eq_228_in1
	// Insensitive connections
	always @(*) begin
		eq_228_in0 = valid ? 32'd4 : 32'd4;
		eq_228_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_230.eq_230_in0
	// controller for eq_230.eq_230_in1
	// Insensitive connections
	always @(*) begin
		eq_230_in0 = valid ? 32'd3 : 32'd3;
		eq_230_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_239.eq_239_in0
	// controller for eq_239.eq_239_in1
	// Insensitive connections
	always @(*) begin
		eq_239_in0 = valid ? 32'd1 : 32'd1;
		eq_239_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_248.eq_248_in0
	// controller for eq_248.eq_248_in1
	// Insensitive connections
	always @(*) begin
		eq_248_in0 = valid ? 32'd3 : 32'd3;
		eq_248_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_257.eq_257_in0
	// controller for eq_257.eq_257_in1
	// Insensitive connections
	always @(*) begin
		eq_257_in0 = valid ? 32'd3 : 32'd3;
		eq_257_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_265.eq_265_in0
	// controller for eq_265.eq_265_in1
	// Insensitive connections
	always @(*) begin
		eq_265_in0 = valid ? 32'd1 : 32'd1;
		eq_265_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_266.eq_266_in0
	// controller for eq_266.eq_266_in1
	// Insensitive connections
	always @(*) begin
		eq_266_in0 = valid ? 32'd2 : 32'd2;
		eq_266_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_268.eq_268_in0
	// controller for eq_268.eq_268_in1
	// Insensitive connections
	always @(*) begin
		eq_268_in0 = valid ? 32'd3 : 32'd3;
		eq_268_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_277.eq_277_in0
	// controller for eq_277.eq_277_in1
	// Insensitive connections
	always @(*) begin
		eq_277_in0 = valid ? 32'd1 : 32'd1;
		eq_277_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_286.eq_286_in0
	// controller for eq_286.eq_286_in1
	// Insensitive connections
	always @(*) begin
		eq_286_in0 = valid ? 32'd3 : 32'd3;
		eq_286_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_295.eq_295_in0
	// controller for eq_295.eq_295_in1
	// Insensitive connections
	always @(*) begin
		eq_295_in0 = valid ? 32'd3 : 32'd3;
		eq_295_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_303.eq_303_in0
	// controller for eq_303.eq_303_in1
	// Insensitive connections
	always @(*) begin
		eq_303_in0 = valid ? 32'd2 : 32'd2;
		eq_303_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_304.eq_304_in0
	// controller for eq_304.eq_304_in1
	// Insensitive connections
	always @(*) begin
		eq_304_in0 = valid ? 32'd3 : 32'd3;
		eq_304_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_306.eq_306_in0
	// controller for eq_306.eq_306_in1
	// Insensitive connections
	always @(*) begin
		eq_306_in0 = valid ? 32'd3 : 32'd3;
		eq_306_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_315.eq_315_in0
	// controller for eq_315.eq_315_in1
	// Insensitive connections
	always @(*) begin
		eq_315_in0 = valid ? 32'd1 : 32'd1;
		eq_315_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_324.eq_324_in0
	// controller for eq_324.eq_324_in1
	// Insensitive connections
	always @(*) begin
		eq_324_in0 = valid ? 32'd3 : 32'd3;
		eq_324_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_333.eq_333_in0
	// controller for eq_333.eq_333_in1
	// Insensitive connections
	always @(*) begin
		eq_333_in0 = valid ? 32'd3 : 32'd3;
		eq_333_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_341.eq_341_in0
	// controller for eq_341.eq_341_in1
	// Insensitive connections
	always @(*) begin
		eq_341_in0 = valid ? 32'd3 : 32'd3;
		eq_341_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_342.eq_342_in0
	// controller for eq_342.eq_342_in1
	// Insensitive connections
	always @(*) begin
		eq_342_in0 = valid ? 32'd4 : 32'd4;
		eq_342_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_344.eq_344_in0
	// controller for eq_344.eq_344_in1
	// Insensitive connections
	always @(*) begin
		eq_344_in0 = valid ? 32'd3 : 32'd3;
		eq_344_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_353.eq_353_in0
	// controller for eq_353.eq_353_in1
	// Insensitive connections
	always @(*) begin
		eq_353_in0 = valid ? 32'd1 : 32'd1;
		eq_353_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_362.eq_362_in0
	// controller for eq_362.eq_362_in1
	// Insensitive connections
	always @(*) begin
		eq_362_in0 = valid ? 32'd3 : 32'd3;
		eq_362_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_371.eq_371_in0
	// controller for eq_371.eq_371_in1
	// Insensitive connections
	always @(*) begin
		eq_371_in0 = valid ? 32'd3 : 32'd3;
		eq_371_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_91.eq_91_in0
	// controller for eq_91.eq_91_in1
	// Insensitive connections
	always @(*) begin
		eq_91_in0 = valid ? 32'd0 : 32'd0;
		eq_91_in1 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
	end
	// controller for eq_92.eq_92_in0
	// controller for eq_92.eq_92_in1
	// Insensitive connections
	always @(*) begin
		eq_92_in0 = valid ? 32'd8 : 32'd8;
		eq_92_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_94.eq_94_in0
	// controller for eq_94.eq_94_in1
	// Insensitive connections
	always @(*) begin
		eq_94_in0 = valid ? 32'd9 : 32'd9;
		eq_94_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_96.eq_96_in0
	// controller for eq_96.eq_96_in1
	// Insensitive connections
	always @(*) begin
		eq_96_in0 = valid ? 32'd0 : 32'd0;
		eq_96_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_97.eq_97_in0
	// controller for eq_97.eq_97_in1
	// Insensitive connections
	always @(*) begin
		eq_97_in0 = valid ? 32'd3 : 32'd3;
		eq_97_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_99.eq_99_in0
	// controller for eq_99.eq_99_in1
	// Insensitive connections
	always @(*) begin
		eq_99_in0 = valid ? 32'd10 : 32'd10;
		eq_99_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for icmp_17.cmp_in0_icmp_17
	// controller for icmp_17.cmp_in1_icmp_17
	// Insensitive connections
	always @(*) begin
		cmp_in0_icmp_17 = valid ? add_out_add_16 : add_out_add_16;
		cmp_in1_icmp_17 = valid ? 32'd4 : 32'd4;
	end
	// controller for in.in_read_valid_reg
	always @(*) begin
		if (andOp_154_out) begin 
			in_read_valid_reg = -(1'd1);
		end else begin
			in_read_valid_reg = 0;
		end
	end
	// controller for notOp_116.notOp_116_in0
	// Insensitive connections
	always @(*) begin
		notOp_116_in0 = valid ? eq_115_out : eq_115_out;
	end
	// controller for notOp_119.notOp_119_in0
	// Insensitive connections
	always @(*) begin
		notOp_119_in0 = valid ? eq_118_out : eq_118_out;
	end
	// controller for notOp_123.notOp_123_in0
	// Insensitive connections
	always @(*) begin
		notOp_123_in0 = valid ? eq_122_out : eq_122_out;
	end
	// controller for notOp_127.notOp_127_in0
	// Insensitive connections
	always @(*) begin
		notOp_127_in0 = valid ? eq_126_out : eq_126_out;
	end
	// controller for notOp_131.notOp_131_in0
	// Insensitive connections
	always @(*) begin
		notOp_131_in0 = valid ? eq_130_out : eq_130_out;
	end
	// controller for notOp_134.notOp_134_in0
	// Insensitive connections
	always @(*) begin
		notOp_134_in0 = valid ? eq_133_out : eq_133_out;
	end
	// controller for notOp_137.notOp_137_in0
	// Insensitive connections
	always @(*) begin
		notOp_137_in0 = valid ? eq_136_out : eq_136_out;
	end
	// controller for notOp_140.notOp_140_in0
	// Insensitive connections
	always @(*) begin
		notOp_140_in0 = valid ? eq_139_out : eq_139_out;
	end
	// controller for notOp_144.notOp_144_in0
	// Insensitive connections
	always @(*) begin
		notOp_144_in0 = valid ? eq_143_out : eq_143_out;
	end
	// controller for notOp_173.notOp_173_in0
	// Insensitive connections
	always @(*) begin
		notOp_173_in0 = valid ? andOp_169_out : andOp_169_out;
	end
	// controller for notOp_175.notOp_175_in0
	// Insensitive connections
	always @(*) begin
		notOp_175_in0 = valid ? andOp_51_out : andOp_51_out;
	end
	// controller for notOp_177.notOp_177_in0
	// Insensitive connections
	always @(*) begin
		notOp_177_in0 = valid ? andOp_66_out : andOp_66_out;
	end
	// controller for notOp_179.notOp_179_in0
	// Insensitive connections
	always @(*) begin
		notOp_179_in0 = valid ? andOp_49_out : andOp_49_out;
	end
	// controller for notOp_181.notOp_181_in0
	// Insensitive connections
	always @(*) begin
		notOp_181_in0 = valid ? andOp_170_out : andOp_170_out;
	end
	// controller for notOp_183.notOp_183_in0
	// Insensitive connections
	always @(*) begin
		notOp_183_in0 = valid ? andOp_171_out : andOp_171_out;
	end
	// controller for notOp_185.notOp_185_in0
	// Insensitive connections
	always @(*) begin
		notOp_185_in0 = valid ? andOp_172_out : andOp_172_out;
	end
	// controller for notOp_187.notOp_187_in0
	// Insensitive connections
	always @(*) begin
		notOp_187_in0 = valid ? andOp_81_out : andOp_81_out;
	end
	// controller for notOp_193.notOp_193_in0
	// Insensitive connections
	always @(*) begin
		notOp_193_in0 = valid ? eq_191_out : eq_191_out;
	end
	// controller for notOp_195.notOp_195_in0
	// Insensitive connections
	always @(*) begin
		notOp_195_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_197.notOp_197_in0
	// Insensitive connections
	always @(*) begin
		notOp_197_in0 = valid ? andOp_192_out : andOp_192_out;
	end
	// controller for notOp_202.notOp_202_in0
	// Insensitive connections
	always @(*) begin
		notOp_202_in0 = valid ? eq_200_out : eq_200_out;
	end
	// controller for notOp_204.notOp_204_in0
	// Insensitive connections
	always @(*) begin
		notOp_204_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_206.notOp_206_in0
	// Insensitive connections
	always @(*) begin
		notOp_206_in0 = valid ? andOp_201_out : andOp_201_out;
	end
	// controller for notOp_211.notOp_211_in0
	// Insensitive connections
	always @(*) begin
		notOp_211_in0 = valid ? eq_209_out : eq_209_out;
	end
	// controller for notOp_213.notOp_213_in0
	// Insensitive connections
	always @(*) begin
		notOp_213_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_215.notOp_215_in0
	// Insensitive connections
	always @(*) begin
		notOp_215_in0 = valid ? andOp_210_out : andOp_210_out;
	end
	// controller for notOp_220.notOp_220_in0
	// Insensitive connections
	always @(*) begin
		notOp_220_in0 = valid ? eq_218_out : eq_218_out;
	end
	// controller for notOp_222.notOp_222_in0
	// Insensitive connections
	always @(*) begin
		notOp_222_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_224.notOp_224_in0
	// Insensitive connections
	always @(*) begin
		notOp_224_in0 = valid ? andOp_219_out : andOp_219_out;
	end
	// controller for notOp_232.notOp_232_in0
	// Insensitive connections
	always @(*) begin
		notOp_232_in0 = valid ? eq_230_out : eq_230_out;
	end
	// controller for notOp_234.notOp_234_in0
	// Insensitive connections
	always @(*) begin
		notOp_234_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_236.notOp_236_in0
	// Insensitive connections
	always @(*) begin
		notOp_236_in0 = valid ? andOp_231_out : andOp_231_out;
	end
	// controller for notOp_241.notOp_241_in0
	// Insensitive connections
	always @(*) begin
		notOp_241_in0 = valid ? eq_239_out : eq_239_out;
	end
	// controller for notOp_243.notOp_243_in0
	// Insensitive connections
	always @(*) begin
		notOp_243_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
	end
	// controller for notOp_245.notOp_245_in0
	// Insensitive connections
	always @(*) begin
		notOp_245_in0 = valid ? andOp_240_out : andOp_240_out;
	end
	// controller for notOp_250.notOp_250_in0
	// Insensitive connections
	always @(*) begin
		notOp_250_in0 = valid ? eq_248_out : eq_248_out;
	end
	// controller for notOp_252.notOp_252_in0
	// Insensitive connections
	always @(*) begin
		notOp_252_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_254.notOp_254_in0
	// Insensitive connections
	always @(*) begin
		notOp_254_in0 = valid ? andOp_249_out : andOp_249_out;
	end
	// controller for notOp_259.notOp_259_in0
	// Insensitive connections
	always @(*) begin
		notOp_259_in0 = valid ? eq_257_out : eq_257_out;
	end
	// controller for notOp_261.notOp_261_in0
	// Insensitive connections
	always @(*) begin
		notOp_261_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_263.notOp_263_in0
	// Insensitive connections
	always @(*) begin
		notOp_263_in0 = valid ? andOp_258_out : andOp_258_out;
	end
	// controller for notOp_270.notOp_270_in0
	// Insensitive connections
	always @(*) begin
		notOp_270_in0 = valid ? eq_268_out : eq_268_out;
	end
	// controller for notOp_272.notOp_272_in0
	// Insensitive connections
	always @(*) begin
		notOp_272_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
	end
	// controller for notOp_274.notOp_274_in0
	// Insensitive connections
	always @(*) begin
		notOp_274_in0 = valid ? andOp_269_out : andOp_269_out;
	end
	// controller for notOp_279.notOp_279_in0
	// Insensitive connections
	always @(*) begin
		notOp_279_in0 = valid ? eq_277_out : eq_277_out;
	end
	// controller for notOp_281.notOp_281_in0
	// Insensitive connections
	always @(*) begin
		notOp_281_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_283.notOp_283_in0
	// Insensitive connections
	always @(*) begin
		notOp_283_in0 = valid ? andOp_278_out : andOp_278_out;
	end
	// controller for notOp_288.notOp_288_in0
	// Insensitive connections
	always @(*) begin
		notOp_288_in0 = valid ? eq_286_out : eq_286_out;
	end
	// controller for notOp_290.notOp_290_in0
	// Insensitive connections
	always @(*) begin
		notOp_290_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_292.notOp_292_in0
	// Insensitive connections
	always @(*) begin
		notOp_292_in0 = valid ? andOp_287_out : andOp_287_out;
	end
	// controller for notOp_297.notOp_297_in0
	// Insensitive connections
	always @(*) begin
		notOp_297_in0 = valid ? eq_295_out : eq_295_out;
	end
	// controller for notOp_299.notOp_299_in0
	// Insensitive connections
	always @(*) begin
		notOp_299_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_301.notOp_301_in0
	// Insensitive connections
	always @(*) begin
		notOp_301_in0 = valid ? andOp_296_out : andOp_296_out;
	end
	// controller for notOp_308.notOp_308_in0
	// Insensitive connections
	always @(*) begin
		notOp_308_in0 = valid ? eq_306_out : eq_306_out;
	end
	// controller for notOp_310.notOp_310_in0
	// Insensitive connections
	always @(*) begin
		notOp_310_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
	end
	// controller for notOp_312.notOp_312_in0
	// Insensitive connections
	always @(*) begin
		notOp_312_in0 = valid ? andOp_307_out : andOp_307_out;
	end
	// controller for notOp_317.notOp_317_in0
	// Insensitive connections
	always @(*) begin
		notOp_317_in0 = valid ? eq_315_out : eq_315_out;
	end
	// controller for notOp_319.notOp_319_in0
	// Insensitive connections
	always @(*) begin
		notOp_319_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_321.notOp_321_in0
	// Insensitive connections
	always @(*) begin
		notOp_321_in0 = valid ? andOp_316_out : andOp_316_out;
	end
	// controller for notOp_326.notOp_326_in0
	// Insensitive connections
	always @(*) begin
		notOp_326_in0 = valid ? eq_324_out : eq_324_out;
	end
	// controller for notOp_328.notOp_328_in0
	// Insensitive connections
	always @(*) begin
		notOp_328_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
	end
	// controller for notOp_330.notOp_330_in0
	// Insensitive connections
	always @(*) begin
		notOp_330_in0 = valid ? andOp_325_out : andOp_325_out;
	end
	// controller for notOp_335.notOp_335_in0
	// Insensitive connections
	always @(*) begin
		notOp_335_in0 = valid ? eq_333_out : eq_333_out;
	end
	// controller for notOp_337.notOp_337_in0
	// Insensitive connections
	always @(*) begin
		notOp_337_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
	end
	// controller for notOp_339.notOp_339_in0
	// Insensitive connections
	always @(*) begin
		notOp_339_in0 = valid ? andOp_334_out : andOp_334_out;
	end
	// controller for notOp_346.notOp_346_in0
	// Insensitive connections
	always @(*) begin
		notOp_346_in0 = valid ? eq_344_out : eq_344_out;
	end
	// controller for notOp_348.notOp_348_in0
	// Insensitive connections
	always @(*) begin
		notOp_348_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_350.notOp_350_in0
	// Insensitive connections
	always @(*) begin
		notOp_350_in0 = valid ? andOp_345_out : andOp_345_out;
	end
	// controller for notOp_355.notOp_355_in0
	// Insensitive connections
	always @(*) begin
		notOp_355_in0 = valid ? eq_353_out : eq_353_out;
	end
	// controller for notOp_357.notOp_357_in0
	// Insensitive connections
	always @(*) begin
		notOp_357_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_359.notOp_359_in0
	// Insensitive connections
	always @(*) begin
		notOp_359_in0 = valid ? andOp_354_out : andOp_354_out;
	end
	// controller for notOp_364.notOp_364_in0
	// Insensitive connections
	always @(*) begin
		notOp_364_in0 = valid ? eq_362_out : eq_362_out;
	end
	// controller for notOp_366.notOp_366_in0
	// Insensitive connections
	always @(*) begin
		notOp_366_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
	end
	// controller for notOp_368.notOp_368_in0
	// Insensitive connections
	always @(*) begin
		notOp_368_in0 = valid ? andOp_363_out : andOp_363_out;
	end
	// controller for notOp_373.notOp_373_in0
	// Insensitive connections
	always @(*) begin
		notOp_373_in0 = valid ? eq_371_out : eq_371_out;
	end
	// controller for notOp_375.notOp_375_in0
	// Insensitive connections
	always @(*) begin
		notOp_375_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
	end
	// controller for notOp_377.notOp_377_in0
	// Insensitive connections
	always @(*) begin
		notOp_377_in0 = valid ? andOp_372_out : andOp_372_out;
	end
	// controller for notOp_42.notOp_42_in0
	// Insensitive connections
	always @(*) begin
		notOp_42_in0 = valid ? andOp_41_out : andOp_41_out;
	end
	// controller for notOp_45.notOp_45_in0
	// Insensitive connections
	always @(*) begin
		notOp_45_in0 = valid ? andOp_44_out : andOp_44_out;
	end
	// controller for notOp_48.notOp_48_in0
	// Insensitive connections
	always @(*) begin
		notOp_48_in0 = valid ? andOp_47_out : andOp_47_out;
	end
	// controller for notOp_50.notOp_50_in0
	// Insensitive connections
	always @(*) begin
		notOp_50_in0 = valid ? in_read_ready : in_read_ready;
	end
	// controller for notOp_54.notOp_54_in0
	// Insensitive connections
	always @(*) begin
		notOp_54_in0 = valid ? andOp_53_out : andOp_53_out;
	end
	// controller for notOp_57.notOp_57_in0
	// Insensitive connections
	always @(*) begin
		notOp_57_in0 = valid ? andOp_56_out : andOp_56_out;
	end
	// controller for notOp_60.notOp_60_in0
	// Insensitive connections
	always @(*) begin
		notOp_60_in0 = valid ? andOp_59_out : andOp_59_out;
	end
	// controller for notOp_63.notOp_63_in0
	// Insensitive connections
	always @(*) begin
		notOp_63_in0 = valid ? andOp_62_out : andOp_62_out;
	end
	// controller for notOp_65.notOp_65_in0
	// Insensitive connections
	always @(*) begin
		notOp_65_in0 = valid ? data_in_4_39_out_data : data_in_4_39_out_data;
	end
	// controller for notOp_69.notOp_69_in0
	// Insensitive connections
	always @(*) begin
		notOp_69_in0 = valid ? andOp_68_out : andOp_68_out;
	end
	// controller for notOp_72.notOp_72_in0
	// Insensitive connections
	always @(*) begin
		notOp_72_in0 = valid ? andOp_71_out : andOp_71_out;
	end
	// controller for notOp_75.notOp_75_in0
	// Insensitive connections
	always @(*) begin
		notOp_75_in0 = valid ? andOp_74_out : andOp_74_out;
	end
	// controller for notOp_78.notOp_78_in0
	// Insensitive connections
	always @(*) begin
		notOp_78_in0 = valid ? andOp_77_out : andOp_77_out;
	end
	// controller for notOp_80.notOp_80_in0
	// Insensitive connections
	always @(*) begin
		notOp_80_in0 = valid ? out_write_ready : out_write_ready;
	end
	// controller for notOp_84.notOp_84_in0
	// Insensitive connections
	always @(*) begin
		notOp_84_in0 = valid ? andOp_83_out : andOp_83_out;
	end
	// controller for notOp_86.notOp_86_in0
	// Insensitive connections
	always @(*) begin
		notOp_86_in0 = valid ? data_in_4_39_out_data : data_in_4_39_out_data;
	end
	// controller for notOp_90.notOp_90_in0
	// Insensitive connections
	always @(*) begin
		notOp_90_in0 = valid ? andOp_89_out : andOp_89_out;
	end
	// controller for orOp_101.orOp_101_in0
	// controller for orOp_101.orOp_101_in1
	// Insensitive connections
	always @(*) begin
		orOp_101_in0 = valid ? eq_100_out : eq_100_out;
		orOp_101_in1 = valid ? andOp_59_out : andOp_59_out;
	end
	// controller for orOp_104.orOp_104_in0
	// controller for orOp_104.orOp_104_in1
	// Insensitive connections
	always @(*) begin
		orOp_104_in0 = valid ? eq_103_out : eq_103_out;
		orOp_104_in1 = valid ? andOp_74_out : andOp_74_out;
	end
	// controller for orOp_106.orOp_106_in0
	// controller for orOp_106.orOp_106_in1
	// Insensitive connections
	always @(*) begin
		orOp_106_in0 = valid ? eq_105_out : eq_105_out;
		orOp_106_in1 = valid ? andOp_89_out : andOp_89_out;
	end
	// controller for orOp_108.orOp_108_in0
	// controller for orOp_108.orOp_108_in1
	// Insensitive connections
	always @(*) begin
		orOp_108_in0 = valid ? eq_107_out : eq_107_out;
		orOp_108_in1 = valid ? andOp_79_out : andOp_79_out;
	end
	// controller for orOp_110.orOp_110_in0
	// controller for orOp_110.orOp_110_in1
	// Insensitive connections
	always @(*) begin
		orOp_110_in0 = valid ? eq_109_out : eq_109_out;
		orOp_110_in1 = valid ? andOp_71_out : andOp_71_out;
	end
	// controller for orOp_113.orOp_113_in0
	// controller for orOp_113.orOp_113_in1
	// Insensitive connections
	always @(*) begin
		orOp_113_in0 = valid ? eq_112_out : eq_112_out;
		orOp_113_in1 = valid ? andOp_64_out : andOp_64_out;
	end
	// controller for orOp_93.orOp_93_in0
	// controller for orOp_93.orOp_93_in1
	// Insensitive connections
	always @(*) begin
		orOp_93_in0 = valid ? eq_92_out : eq_92_out;
		orOp_93_in1 = valid ? andOp_56_out : andOp_56_out;
	end
	// controller for orOp_95.orOp_95_in0
	// controller for orOp_95.orOp_95_in1
	// Insensitive connections
	always @(*) begin
		orOp_95_in0 = valid ? eq_94_out : eq_94_out;
		orOp_95_in1 = valid ? andOp_44_out : andOp_44_out;
	end
	// controller for orOp_98.orOp_98_in0
	// controller for orOp_98.orOp_98_in1
	// Insensitive connections
	always @(*) begin
		orOp_98_in0 = valid ? eq_97_out : eq_97_out;
		orOp_98_in1 = valid ? andOp_41_out : andOp_41_out;
	end
	// controller for out.out_in_data_reg
	always @(*) begin
		if (andOp_166_out) begin 
			out_in_data_reg = rdata_ram_0;
		end else begin
			out_in_data_reg = 0;
		end
	end
	// controller for out.out_write_valid_reg
	always @(*) begin
		if (andOp_165_out) begin 
			out_write_valid_reg = -(1'd1);
		end else begin
			out_write_valid_reg = 0;
		end
	end
	// controller for phi_9.phi_in_phi_9
	// controller for phi_9.phi_last_block_phi_9
	// controller for phi_9.phi_s_phi_9
	// Insensitive connections
	always @(*) begin
		phi_in_phi_9 = valid ? concat_157_out : concat_157_out;
		phi_last_block_phi_9 = valid ? bb_3_predecessor_in_state_1_out_data : bb_3_predecessor_in_state_1_out_data;
		phi_s_phi_9 = valid ? concat_158_out : concat_158_out;
	end
	// controller for ram_0.raddr_ram_0_reg
	always @(*) begin
		if (andOp_150_out) begin 
			raddr_ram_0_reg = 32'd0;
		end else if (andOp_152_out) begin 
			raddr_ram_0_reg = 32'd0;
		end else begin
			raddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.waddr_ram_0_reg
	always @(*) begin
		if (andOp_149_out) begin 
			waddr_ram_0_reg = 32'd0;
		end else if (andOp_151_out) begin 
			waddr_ram_0_reg = 32'd0;
		end else begin
			waddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wdata_ram_0_reg
	always @(*) begin
		if (andOp_149_out) begin 
			wdata_ram_0_reg = 32'd0;
		end else if (andOp_151_out) begin 
			wdata_ram_0_reg = add_out_add_14;
		end else begin
			wdata_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wen_ram_0_reg
	always @(*) begin
		if (andOp_149_out) begin 
			wen_ram_0_reg = 1'd1;
		end else if (andOp_151_out) begin 
			wen_ram_0_reg = 1'd1;
		end else begin
			wen_ram_0_reg = 0;
		end
	end
	// controller for ret_27.valid_reg
	always @(*) begin
		if (andOp_168_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// controller for tmp_output_160.tmp_output_160_in_data
	always @(*) begin
		if (eq_161_out) begin 
			tmp_output_160_in_data = in_out_data;
		end else begin
			tmp_output_160_in_data = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			data_store_0_0 <= 0;
		end else begin
			if (andOp_192_out) begin
				data_store_0_0 <= in_out_data;
			end
			if (andOp_198_out) begin
				data_store_0_0 <= data_in_0_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_2 <= 0;
		end else begin
			if (andOp_201_out) begin
				data_store_0_2 <= phi_out_phi_9;
			end
			if (andOp_207_out) begin
				data_store_0_2 <= data_in_0_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_4 <= 0;
		end else begin
			if (andOp_210_out) begin
				data_store_0_4 <= add_out_add_16;
			end
			if (andOp_216_out) begin
				data_store_0_4 <= data_in_0_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_6 <= 0;
		end else begin
			if (andOp_219_out) begin
				data_store_0_6 <= cmp_out_icmp_17;
			end
			if (andOp_225_out) begin
				data_store_0_6 <= data_in_0_7_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_10 <= 0;
		end else begin
			if (andOp_240_out) begin
				data_store_1_10 <= phi_out_phi_9;
			end
			if (andOp_246_out) begin
				data_store_1_10 <= data_in_1_11_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_12 <= 0;
		end else begin
			if (andOp_249_out) begin
				data_store_1_12 <= add_out_add_16;
			end
			if (andOp_255_out) begin
				data_store_1_12 <= data_in_1_13_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_14 <= 0;
		end else begin
			if (andOp_258_out) begin
				data_store_1_14 <= cmp_out_icmp_17;
			end
			if (andOp_264_out) begin
				data_store_1_14 <= data_in_1_15_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_8 <= 0;
		end else begin
			if (andOp_231_out) begin
				data_store_1_8 <= in_out_data;
			end
			if (andOp_237_out) begin
				data_store_1_8 <= data_in_1_9_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_16 <= 0;
		end else begin
			if (andOp_269_out) begin
				data_store_2_16 <= in_out_data;
			end
			if (andOp_275_out) begin
				data_store_2_16 <= data_in_2_17_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_18 <= 0;
		end else begin
			if (andOp_278_out) begin
				data_store_2_18 <= phi_out_phi_9;
			end
			if (andOp_284_out) begin
				data_store_2_18 <= data_in_2_19_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_20 <= 0;
		end else begin
			if (andOp_287_out) begin
				data_store_2_20 <= add_out_add_16;
			end
			if (andOp_293_out) begin
				data_store_2_20 <= data_in_2_21_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_22 <= 0;
		end else begin
			if (andOp_296_out) begin
				data_store_2_22 <= cmp_out_icmp_17;
			end
			if (andOp_302_out) begin
				data_store_2_22 <= data_in_2_23_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_24 <= 0;
		end else begin
			if (andOp_307_out) begin
				data_store_3_24 <= in_out_data;
			end
			if (andOp_313_out) begin
				data_store_3_24 <= data_in_3_25_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_26 <= 0;
		end else begin
			if (andOp_316_out) begin
				data_store_3_26 <= phi_out_phi_9;
			end
			if (andOp_322_out) begin
				data_store_3_26 <= data_in_3_27_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_28 <= 0;
		end else begin
			if (andOp_325_out) begin
				data_store_3_28 <= add_out_add_16;
			end
			if (andOp_331_out) begin
				data_store_3_28 <= data_in_3_29_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_30 <= 0;
		end else begin
			if (andOp_334_out) begin
				data_store_3_30 <= cmp_out_icmp_17;
			end
			if (andOp_340_out) begin
				data_store_3_30 <= data_in_3_31_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_32 <= 0;
		end else begin
			if (andOp_345_out) begin
				data_store_4_32 <= in_out_data;
			end
			if (andOp_351_out) begin
				data_store_4_32 <= data_in_4_33_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_34 <= 0;
		end else begin
			if (andOp_354_out) begin
				data_store_4_34 <= phi_out_phi_9;
			end
			if (andOp_360_out) begin
				data_store_4_34 <= data_in_4_35_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_36 <= 0;
		end else begin
			if (andOp_363_out) begin
				data_store_4_36 <= add_out_add_16;
			end
			if (andOp_369_out) begin
				data_store_4_36 <= data_in_4_37_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_38 <= 0;
		end else begin
			if (andOp_372_out) begin
				data_store_4_38 <= cmp_out_icmp_17;
			end
			if (andOp_378_out) begin
				data_store_4_38 <= data_in_4_39_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_169_out) begin
				global_state <= 32'd1;
			end
			if (andOp_170_out) begin
				global_state <= 32'd3;
			end
			if (andOp_171_out) begin
				global_state <= 32'd4;
			end
			if (andOp_172_out) begin
				global_state <= 32'd4;
			end
			if (andOp_49_out) begin
				global_state <= 32'd2;
			end
			if (andOp_51_out) begin
				global_state <= 32'd1;
			end
			if (andOp_66_out) begin
				global_state <= 32'd1;
			end
			if (andOp_81_out) begin
				global_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (1'd1) begin
				state_0_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_169_out) begin
				state_1_entry_BB_reg <= 32'd0;
			end
			if (andOp_51_out) begin
				state_1_entry_BB_reg <= 32'd9;
			end
			if (andOp_66_out) begin
				state_1_entry_BB_reg <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_169_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_178_out) begin
				state_1_is_active <= 1'd0;
			end
			if (andOp_51_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_66_out) begin
				state_1_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_169_out) begin
				state_1_last_BB_reg <= bb_0_predecessor_in_state_0_out_data;
			end
			if (andOp_51_out) begin
				state_1_last_BB_reg <= 32'd9;
			end
			if (andOp_66_out) begin
				state_1_last_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_169_out) begin
				state_1_last_state <= 32'd0;
			end
			if (andOp_51_out) begin
				state_1_last_state <= 32'd1;
			end
			if (andOp_66_out) begin
				state_1_last_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_49_out) begin
				state_2_entry_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_180_out) begin
				state_2_is_active <= 1'd0;
			end
			if (andOp_49_out) begin
				state_2_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_49_out) begin
				state_2_last_BB_reg <= 32'd9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_49_out) begin
				state_2_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_170_out) begin
				state_3_entry_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_170_out) begin
				state_3_is_active <= 1'd1;
			end
			if (andOp_182_out) begin
				state_3_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_170_out) begin
				state_3_last_BB_reg <= bb_10_predecessor_in_state_2_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_state <= 0;
		end else begin
			if (andOp_170_out) begin
				state_3_last_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_171_out) begin
				state_4_entry_BB_reg <= 32'd4;
			end
			if (andOp_172_out) begin
				state_4_entry_BB_reg <= 32'd2;
			end
			if (andOp_81_out) begin
				state_4_entry_BB_reg <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_171_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_172_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_188_out) begin
				state_4_is_active <= 1'd0;
			end
			if (andOp_81_out) begin
				state_4_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_171_out) begin
				state_4_last_BB_reg <= bb_4_predecessor_in_state_3_out_data;
			end
			if (andOp_172_out) begin
				state_4_last_BB_reg <= bb_2_predecessor_in_state_4_out_data;
			end
			if (andOp_81_out) begin
				state_4_last_BB_reg <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_state <= 0;
		end else begin
			if (andOp_171_out) begin
				state_4_last_state <= 32'd3;
			end
			if (andOp_172_out) begin
				state_4_last_state <= 32'd4;
			end
			if (andOp_81_out) begin
				state_4_last_state <= 32'd4;
			end
		end
	end

endmodule

