module smul_fifo(input [0:0] clk, input [0:0] rst, output [0:0] valid, output [31:0] arg_0_in_data, input [31:0] arg_0_out_data, input [0:0] arg_0_read_ready, output [0:0] arg_0_read_valid, input [0:0] arg_0_write_ready, output [0:0] arg_0_write_valid, output [31:0] arg_1_in_data, input [31:0] arg_1_out_data, input [0:0] arg_1_read_ready, output [0:0] arg_1_read_valid, input [0:0] arg_1_write_ready, output [0:0] arg_1_write_valid);

	reg [0:0] valid_reg;
	reg [31:0] arg_0_in_data_reg;
	reg [0:0] arg_0_read_valid_reg;
	reg [0:0] arg_0_write_valid_reg;
	reg [31:0] arg_1_in_data_reg;
	reg [0:0] arg_1_read_valid_reg;
	reg [0:0] arg_1_write_valid_reg;

	assign valid = valid_reg;
	assign arg_0_in_data = arg_0_in_data_reg;
	assign arg_0_read_valid = arg_0_read_valid_reg;
	assign arg_0_write_valid = arg_0_write_valid_reg;
	assign arg_1_in_data = arg_1_in_data_reg;
	assign arg_1_read_valid = arg_1_read_valid_reg;
	assign arg_1_write_valid = arg_1_write_valid_reg;

	// Start debug wires and ports

	initial begin
	end



	always @(posedge clk) begin
		if (!((!(andOp_33_out === 1) || andOp_49_out !== 1))) begin $display("assertion((!(andOp_33_out === 1) || andOp_49_out !== 1)) failed: Problem: Overlapping last basic block transition"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_49_out === 1) || andOp_33_out !== 1))) begin $display("assertion((!(andOp_49_out === 1) || andOp_33_out !== 1)) failed: Problem: Overlapping last basic block transition"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_34_out === 1) || andOp_46_out !== 1))) begin $display("assertion((!(andOp_34_out === 1) || andOp_46_out !== 1)) failed: Problem: Overlapping last basic block transition"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_46_out === 1) || andOp_34_out !== 1))) begin $display("assertion((!(andOp_46_out === 1) || andOp_34_out !== 1)) failed: Problem: Overlapping last basic block transition"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_113_out === 1) || andOp_44_out !== 1))) begin $display("assertion((!(andOp_113_out === 1) || andOp_44_out !== 1)) failed: Problem: Overlapping last basic block transition"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_44_out === 1) || andOp_113_out !== 1))) begin $display("assertion((!(andOp_44_out === 1) || andOp_113_out !== 1)) failed: Problem: Overlapping last basic block transition"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_33_out === 1) || andOp_49_out !== 1))) begin $display("assertion((!(andOp_33_out === 1) || andOp_49_out !== 1)) failed: Problem: Overlapping block transition"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_49_out === 1) || andOp_33_out !== 1))) begin $display("assertion((!(andOp_49_out === 1) || andOp_33_out !== 1)) failed: Problem: Overlapping block transition"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_34_out === 1) || andOp_46_out !== 1))) begin $display("assertion((!(andOp_34_out === 1) || andOp_46_out !== 1)) failed: Problem: Overlapping block transition"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_46_out === 1) || andOp_34_out !== 1))) begin $display("assertion((!(andOp_46_out === 1) || andOp_34_out !== 1)) failed: Problem: Overlapping block transition"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_113_out === 1) || andOp_44_out !== 1))) begin $display("assertion((!(andOp_113_out === 1) || andOp_44_out !== 1)) failed: Problem: Overlapping block transition"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_44_out === 1) || andOp_113_out !== 1))) begin $display("assertion((!(andOp_44_out === 1) || andOp_113_out !== 1)) failed: Problem: Overlapping block transition"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_117_out === 1) || andOp_33_out !== 1))) begin $display("assertion((!(andOp_117_out === 1) || andOp_33_out !== 1)) failed: Overlapping state active transition for state 0"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_117_out === 1) || andOp_49_out !== 1))) begin $display("assertion((!(andOp_117_out === 1) || andOp_49_out !== 1)) failed: Overlapping state active transition for state 0"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_33_out === 1) || andOp_117_out !== 1))) begin $display("assertion((!(andOp_33_out === 1) || andOp_117_out !== 1)) failed: Overlapping state active transition for state 0"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_33_out === 1) || andOp_49_out !== 1))) begin $display("assertion((!(andOp_33_out === 1) || andOp_49_out !== 1)) failed: Overlapping state active transition for state 0"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_49_out === 1) || andOp_117_out !== 1))) begin $display("assertion((!(andOp_49_out === 1) || andOp_117_out !== 1)) failed: Overlapping state active transition for state 0"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_49_out === 1) || andOp_33_out !== 1))) begin $display("assertion((!(andOp_49_out === 1) || andOp_33_out !== 1)) failed: Overlapping state active transition for state 0"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_119_out === 1) || andOp_31_out !== 1))) begin $display("assertion((!(andOp_119_out === 1) || andOp_31_out !== 1)) failed: Overlapping state active transition for state 1"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_31_out === 1) || andOp_119_out !== 1))) begin $display("assertion((!(andOp_31_out === 1) || andOp_119_out !== 1)) failed: Overlapping state active transition for state 1"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_112_out === 1) || andOp_121_out !== 1))) begin $display("assertion((!(andOp_112_out === 1) || andOp_121_out !== 1)) failed: Overlapping state active transition for state 2"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_121_out === 1) || andOp_112_out !== 1))) begin $display("assertion((!(andOp_121_out === 1) || andOp_112_out !== 1)) failed: Overlapping state active transition for state 2"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_125_out === 1) || andOp_34_out !== 1))) begin $display("assertion((!(andOp_125_out === 1) || andOp_34_out !== 1)) failed: Overlapping state active transition for state 3"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_125_out === 1) || andOp_46_out !== 1))) begin $display("assertion((!(andOp_125_out === 1) || andOp_46_out !== 1)) failed: Overlapping state active transition for state 3"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_34_out === 1) || andOp_125_out !== 1))) begin $display("assertion((!(andOp_34_out === 1) || andOp_125_out !== 1)) failed: Overlapping state active transition for state 3"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_34_out === 1) || andOp_46_out !== 1))) begin $display("assertion((!(andOp_34_out === 1) || andOp_46_out !== 1)) failed: Overlapping state active transition for state 3"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_46_out === 1) || andOp_125_out !== 1))) begin $display("assertion((!(andOp_46_out === 1) || andOp_125_out !== 1)) failed: Overlapping state active transition for state 3"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_46_out === 1) || andOp_34_out !== 1))) begin $display("assertion((!(andOp_46_out === 1) || andOp_34_out !== 1)) failed: Overlapping state active transition for state 3"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_113_out === 1) || andOp_129_out !== 1))) begin $display("assertion((!(andOp_113_out === 1) || andOp_129_out !== 1)) failed: Overlapping state active transition for state 4"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_113_out === 1) || andOp_44_out !== 1))) begin $display("assertion((!(andOp_113_out === 1) || andOp_44_out !== 1)) failed: Overlapping state active transition for state 4"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_129_out === 1) || andOp_113_out !== 1))) begin $display("assertion((!(andOp_129_out === 1) || andOp_113_out !== 1)) failed: Overlapping state active transition for state 4"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_129_out === 1) || andOp_44_out !== 1))) begin $display("assertion((!(andOp_129_out === 1) || andOp_44_out !== 1)) failed: Overlapping state active transition for state 4"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_44_out === 1) || andOp_113_out !== 1))) begin $display("assertion((!(andOp_44_out === 1) || andOp_113_out !== 1)) failed: Overlapping state active transition for state 4"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_44_out === 1) || andOp_129_out !== 1))) begin $display("assertion((!(andOp_44_out === 1) || andOp_129_out !== 1)) failed: Overlapping state active transition for state 4"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_1_is_active) || !(1'd0)))) begin $display("assertion((!(state_1_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_2_is_active) || !(1'd0)))) begin $display("assertion((!(state_2_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_3_is_active) || !(1'd0)))) begin $display("assertion((!(state_3_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_4_is_active) || !(1'd0)))) begin $display("assertion((!(state_4_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_1_is_active) || !(1'd0)))) begin $display("assertion((!(state_1_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_2_is_active) || !(1'd0)))) begin $display("assertion((!(state_2_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_3_is_active) || !(1'd0)))) begin $display("assertion((!(state_3_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_4_is_active) || !(1'd0)))) begin $display("assertion((!(state_4_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_0_is_active) || !(1'd0)))) begin $display("assertion((!(state_0_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_1_is_active) || !(1'd0)))) begin $display("assertion((!(state_1_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_2_is_active) || !(1'd0)))) begin $display("assertion((!(state_2_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_4_is_active) || !(1'd0)))) begin $display("assertion((!(state_4_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_0_is_active) || !(1'd0)))) begin $display("assertion((!(state_0_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_1_is_active) || !(1'd0)))) begin $display("assertion((!(state_1_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_2_is_active) || !(1'd0)))) begin $display("assertion((!(state_2_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_3_is_active) || !(1'd0)))) begin $display("assertion((!(state_3_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_0_is_active) || !(1'd0)))) begin $display("assertion((!(state_0_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_1_is_active) || !(1'd0)))) begin $display("assertion((!(state_1_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_2_is_active) || !(1'd0)))) begin $display("assertion((!(state_2_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_3_is_active) || !(1'd0)))) begin $display("assertion((!(state_3_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_1_is_active) || !(1'd0)))) begin $display("assertion((!(state_1_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_2_is_active) || !(1'd0)))) begin $display("assertion((!(state_2_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_3_is_active) || !(1'd0)))) begin $display("assertion((!(state_3_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_4_is_active) || !(1'd0)))) begin $display("assertion((!(state_4_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_1_is_active) || !(1'd0)))) begin $display("assertion((!(state_1_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_2_is_active) || !(1'd0)))) begin $display("assertion((!(state_2_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_3_is_active) || !(1'd0)))) begin $display("assertion((!(state_3_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_4_is_active) || !(1'd0)))) begin $display("assertion((!(state_4_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_0_is_active) || !(1'd0)))) begin $display("assertion((!(state_0_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_3_is_active) || !(1'd0)))) begin $display("assertion((!(state_3_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_4_is_active) || !(1'd0)))) begin $display("assertion((!(state_4_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_0_is_active) || !(1'd0)))) begin $display("assertion((!(state_0_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_1_is_active) || !(1'd0)))) begin $display("assertion((!(state_1_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_2_is_active) || !(1'd0)))) begin $display("assertion((!(state_2_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_4_is_active) || !(1'd0)))) begin $display("assertion((!(state_4_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_0_is_active) || !(1'd0)))) begin $display("assertion((!(state_0_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_1_is_active) || !(1'd0)))) begin $display("assertion((!(state_1_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_2_is_active) || !(1'd0)))) begin $display("assertion((!(state_2_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_4_is_active) || !(1'd0)))) begin $display("assertion((!(state_4_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_0_is_active) || !(1'd0)))) begin $display("assertion((!(state_0_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_1_is_active) || !(1'd0)))) begin $display("assertion((!(state_1_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_2_is_active) || !(1'd0)))) begin $display("assertion((!(state_2_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(state_3_is_active) || !(1'd0)))) begin $display("assertion((!(state_3_is_active) || !(1'd0)))"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(notOp_143_out || icmp_icmp18_in0 !== 32'dx)) begin $display("assertion(notOp_143_out || icmp_icmp18_in0 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(notOp_144_out || icmp_icmp18_in1 !== 32'dx)) begin $display("assertion(notOp_144_out || icmp_icmp18_in1 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_145_out) || add_add6_in0 !== 32'dx)) begin $display("assertion(!(andOp_145_out) || add_add6_in0 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_145_out) || add_add6_in1 !== 32'dx)) begin $display("assertion(!(andOp_145_out) || add_add6_in1 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_146_out) || mul_mul14_in0 !== 32'dx)) begin $display("assertion(!(andOp_146_out) || mul_mul14_in0 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!(!(andOp_146_out) || mul_mul14_in1 !== 32'dx)) begin $display("assertion(!(andOp_146_out) || mul_mul14_in1 !== 32'dx)"); $finish(); end
	end

	always @(posedge clk) begin
		if (!((!(andOp_147_out) || phi_phi5_out !== 'dx))) begin $display("assertion((!(andOp_147_out) || phi_phi5_out !== 'dx))"); $finish(); end
	end




	// End debug wires and ports

	// Start Functional Units
	br_dummy br_unit();

	wire [63:0] phi_phi5_in;
	wire [31:0] phi_phi5_last_block;
	wire [63:0] phi_phi5_s;
	wire [31:0] phi_phi5_out;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_phi5(.in(phi_phi5_in), .last_block(phi_phi5_last_block), .out(phi_phi5_out), .s(phi_phi5_s));

	wire [31:0] add_add6_in0;
	wire [31:0] add_add6_in1;
	wire [31:0] add_add6_out;
	add #(.WIDTH(32)) add_add6(.in0(add_add6_in0), .in1(add_add6_in1), .out(add_add6_out));

	wire [31:0] mul_mul14_in0;
	wire [31:0] mul_mul14_in1;
	wire [31:0] mul_mul14_out;
	mul #(.WIDTH(32)) mul_mul14(.in0(mul_mul14_in0), .in1(mul_mul14_in1), .out(mul_mul14_out));

	wire [31:0] icmp_icmp18_in0;
	wire [31:0] icmp_icmp18_in1;
	wire [0:0] icmp_icmp18_out;
	ne #(.WIDTH(32)) icmp_icmp18(.in0(icmp_icmp18_in0), .in1(icmp_icmp18_in1), .out(icmp_icmp18_out));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] bb_1_active_in_state_0_in_data;
	wire [0:0] bb_1_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_0(.in_data(bb_1_active_in_state_0_in_data), .out_data(bb_1_active_in_state_0_out_data));

	reg [31:0] bb_1_predecessor_in_state_0_in_data;
	wire [31:0] bb_1_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_0(.in_data(bb_1_predecessor_in_state_0_in_data), .out_data(bb_1_predecessor_in_state_0_out_data));

	reg [0:0] br_1_happened_in_state_0_in_data;
	wire [0:0] br_1_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened_in_state_0(.in_data(br_1_happened_in_state_0_in_data), .out_data(br_1_happened_in_state_0_out_data));

	reg [0:0] bb_5_active_in_state_0_in_data;
	wire [0:0] bb_5_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_5_active_in_state_0(.in_data(bb_5_active_in_state_0_in_data), .out_data(bb_5_active_in_state_0_out_data));

	reg [31:0] bb_5_predecessor_in_state_0_in_data;
	wire [31:0] bb_5_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_5_predecessor_in_state_0(.in_data(bb_5_predecessor_in_state_0_in_data), .out_data(bb_5_predecessor_in_state_0_out_data));

	reg [0:0] br_5_happened_in_state_0_in_data;
	wire [0:0] br_5_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_5_happened_in_state_0(.in_data(br_5_happened_in_state_0_in_data), .out_data(br_5_happened_in_state_0_out_data));

	reg [0:0] bb_6_active_in_state_0_in_data;
	wire [0:0] bb_6_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_6_active_in_state_0(.in_data(bb_6_active_in_state_0_in_data), .out_data(bb_6_active_in_state_0_out_data));

	reg [31:0] bb_6_predecessor_in_state_0_in_data;
	wire [31:0] bb_6_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_6_predecessor_in_state_0(.in_data(bb_6_predecessor_in_state_0_in_data), .out_data(bb_6_predecessor_in_state_0_out_data));

	reg [0:0] br_6_happened_in_state_0_in_data;
	wire [0:0] br_6_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_6_happened_in_state_0(.in_data(br_6_happened_in_state_0_in_data), .out_data(br_6_happened_in_state_0_out_data));

	reg [0:0] bb_7_active_in_state_1_in_data;
	wire [0:0] bb_7_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_7_active_in_state_1(.in_data(bb_7_active_in_state_1_in_data), .out_data(bb_7_active_in_state_1_out_data));

	reg [31:0] bb_7_predecessor_in_state_1_in_data;
	wire [31:0] bb_7_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_7_predecessor_in_state_1(.in_data(bb_7_predecessor_in_state_1_in_data), .out_data(bb_7_predecessor_in_state_1_out_data));

	reg [0:0] br_7_happened_in_state_1_in_data;
	wire [0:0] br_7_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_7_happened_in_state_1(.in_data(br_7_happened_in_state_1_in_data), .out_data(br_7_happened_in_state_1_out_data));

	reg [0:0] bb_7_active_in_state_2_in_data;
	wire [0:0] bb_7_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_7_active_in_state_2(.in_data(bb_7_active_in_state_2_in_data), .out_data(bb_7_active_in_state_2_out_data));

	reg [31:0] bb_7_predecessor_in_state_2_in_data;
	wire [31:0] bb_7_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_7_predecessor_in_state_2(.in_data(bb_7_predecessor_in_state_2_in_data), .out_data(bb_7_predecessor_in_state_2_out_data));

	reg [0:0] br_7_happened_in_state_2_in_data;
	wire [0:0] br_7_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_7_happened_in_state_2(.in_data(br_7_happened_in_state_2_in_data), .out_data(br_7_happened_in_state_2_out_data));

	reg [0:0] bb_2_active_in_state_3_in_data;
	wire [0:0] bb_2_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_3(.in_data(bb_2_active_in_state_3_in_data), .out_data(bb_2_active_in_state_3_out_data));

	reg [31:0] bb_2_predecessor_in_state_3_in_data;
	wire [31:0] bb_2_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_3(.in_data(bb_2_predecessor_in_state_3_in_data), .out_data(bb_2_predecessor_in_state_3_out_data));

	reg [0:0] br_2_happened_in_state_3_in_data;
	wire [0:0] br_2_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_2_happened_in_state_3(.in_data(br_2_happened_in_state_3_in_data), .out_data(br_2_happened_in_state_3_out_data));

	reg [0:0] bb_8_active_in_state_3_in_data;
	wire [0:0] bb_8_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active_in_state_3(.in_data(bb_8_active_in_state_3_in_data), .out_data(bb_8_active_in_state_3_out_data));

	reg [31:0] bb_8_predecessor_in_state_3_in_data;
	wire [31:0] bb_8_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor_in_state_3(.in_data(bb_8_predecessor_in_state_3_in_data), .out_data(bb_8_predecessor_in_state_3_out_data));

	reg [0:0] br_8_happened_in_state_3_in_data;
	wire [0:0] br_8_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_8_happened_in_state_3(.in_data(br_8_happened_in_state_3_in_data), .out_data(br_8_happened_in_state_3_out_data));

	reg [0:0] bb_9_active_in_state_3_in_data;
	wire [0:0] bb_9_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_9_active_in_state_3(.in_data(bb_9_active_in_state_3_in_data), .out_data(bb_9_active_in_state_3_out_data));

	reg [31:0] bb_9_predecessor_in_state_3_in_data;
	wire [31:0] bb_9_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_9_predecessor_in_state_3(.in_data(bb_9_predecessor_in_state_3_in_data), .out_data(bb_9_predecessor_in_state_3_out_data));

	reg [0:0] br_9_happened_in_state_3_in_data;
	wire [0:0] br_9_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_9_happened_in_state_3(.in_data(br_9_happened_in_state_3_in_data), .out_data(br_9_happened_in_state_3_out_data));

	reg [0:0] bb_4_active_in_state_4_in_data;
	wire [0:0] bb_4_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_4(.in_data(bb_4_active_in_state_4_in_data), .out_data(bb_4_active_in_state_4_out_data));

	reg [31:0] bb_4_predecessor_in_state_4_in_data;
	wire [31:0] bb_4_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_4(.in_data(bb_4_predecessor_in_state_4_in_data), .out_data(bb_4_predecessor_in_state_4_out_data));

	reg [0:0] bb_3_active_in_state_4_in_data;
	wire [0:0] bb_3_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_4(.in_data(bb_3_active_in_state_4_in_data), .out_data(bb_3_active_in_state_4_out_data));

	reg [31:0] bb_3_predecessor_in_state_4_in_data;
	wire [31:0] bb_3_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_4(.in_data(bb_3_predecessor_in_state_4_in_data), .out_data(bb_3_predecessor_in_state_4_out_data));

	reg [0:0] br_3_happened_in_state_4_in_data;
	wire [0:0] br_3_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_4(.in_data(br_3_happened_in_state_4_in_data), .out_data(br_3_happened_in_state_4_out_data));

	reg [0:0] bb_10_active_in_state_4_in_data;
	wire [0:0] bb_10_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_4(.in_data(bb_10_active_in_state_4_in_data), .out_data(bb_10_active_in_state_4_out_data));

	reg [31:0] bb_10_predecessor_in_state_4_in_data;
	wire [31:0] bb_10_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_4(.in_data(bb_10_predecessor_in_state_4_in_data), .out_data(bb_10_predecessor_in_state_4_out_data));

	reg [0:0] br_10_happened_in_state_4_in_data;
	wire [0:0] br_10_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_4(.in_data(br_10_happened_in_state_4_in_data), .out_data(br_10_happened_in_state_4_out_data));

	reg [31:0] data_in_0_1_in_data;
	wire [31:0] data_in_0_1_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_1(.in_data(data_in_0_1_in_data), .out_data(data_in_0_1_out_data));

	reg [31:0] data_in_0_3_in_data;
	wire [31:0] data_in_0_3_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_3(.in_data(data_in_0_3_in_data), .out_data(data_in_0_3_out_data));

	reg [31:0] data_in_1_5_in_data;
	wire [31:0] data_in_1_5_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_5(.in_data(data_in_1_5_in_data), .out_data(data_in_1_5_out_data));

	reg [31:0] data_in_1_7_in_data;
	wire [31:0] data_in_1_7_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_7(.in_data(data_in_1_7_in_data), .out_data(data_in_1_7_out_data));

	reg [31:0] data_in_2_10_in_data;
	wire [31:0] data_in_2_10_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_10(.in_data(data_in_2_10_in_data), .out_data(data_in_2_10_out_data));

	reg [31:0] data_in_2_12_in_data;
	wire [31:0] data_in_2_12_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_12(.in_data(data_in_2_12_in_data), .out_data(data_in_2_12_out_data));

	reg [31:0] data_in_3_14_in_data;
	wire [31:0] data_in_3_14_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_14(.in_data(data_in_3_14_in_data), .out_data(data_in_3_14_out_data));

	reg [31:0] data_in_3_16_in_data;
	wire [31:0] data_in_3_16_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_16(.in_data(data_in_3_16_in_data), .out_data(data_in_3_16_out_data));

	reg [31:0] data_in_3_18_in_data;
	wire [31:0] data_in_3_18_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_18(.in_data(data_in_3_18_in_data), .out_data(data_in_3_18_out_data));

	reg [31:0] data_in_4_20_in_data;
	wire [31:0] data_in_4_20_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_20(.in_data(data_in_4_20_in_data), .out_data(data_in_4_20_out_data));

	reg [31:0] data_in_4_22_in_data;
	wire [31:0] data_in_4_22_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_22(.in_data(data_in_4_22_in_data), .out_data(data_in_4_22_out_data));

	wire [0:0] andOp_23_in0;
	wire [0:0] andOp_23_in1;
	wire [0:0] andOp_23_out;
	andOp #(.WIDTH(1)) andOp_23(.in0(andOp_23_in0), .in1(andOp_23_in1), .out(andOp_23_out));

	wire [0:0] notOp_24_in0;
	wire [0:0] notOp_24_out;
	notOp #(.WIDTH(1)) notOp_24(.in(notOp_24_in0), .out(notOp_24_out));

	wire [0:0] andOp_25_in0;
	wire [0:0] andOp_25_in1;
	wire [0:0] andOp_25_out;
	andOp #(.WIDTH(1)) andOp_25(.in0(andOp_25_in0), .in1(andOp_25_in1), .out(andOp_25_out));

	wire [0:0] notOp_26_in0;
	wire [0:0] notOp_26_out;
	notOp #(.WIDTH(1)) notOp_26(.in(notOp_26_in0), .out(notOp_26_out));

	wire [0:0] andOp_27_in0;
	wire [0:0] andOp_27_in1;
	wire [0:0] andOp_27_out;
	andOp #(.WIDTH(1)) andOp_27(.in0(andOp_27_in0), .in1(andOp_27_in1), .out(andOp_27_out));

	wire [0:0] notOp_28_in0;
	wire [0:0] notOp_28_out;
	notOp #(.WIDTH(1)) notOp_28(.in(notOp_28_in0), .out(notOp_28_out));

	wire [0:0] andOp_29_in0;
	wire [0:0] andOp_29_in1;
	wire [0:0] andOp_29_out;
	andOp #(.WIDTH(1)) andOp_29(.in0(andOp_29_in0), .in1(andOp_29_in1), .out(andOp_29_out));

	wire [0:0] notOp_30_in0;
	wire [0:0] notOp_30_out;
	notOp #(.WIDTH(1)) notOp_30(.in(notOp_30_in0), .out(notOp_30_out));

	wire [0:0] andOp_31_in0;
	wire [0:0] andOp_31_in1;
	wire [0:0] andOp_31_out;
	andOp #(.WIDTH(1)) andOp_31(.in0(andOp_31_in0), .in1(andOp_31_in1), .out(andOp_31_out));

	wire [0:0] notOp_32_in0;
	wire [0:0] notOp_32_out;
	notOp #(.WIDTH(1)) notOp_32(.in(notOp_32_in0), .out(notOp_32_out));

	wire [0:0] andOp_33_in0;
	wire [0:0] andOp_33_in1;
	wire [0:0] andOp_33_out;
	andOp #(.WIDTH(1)) andOp_33(.in0(andOp_33_in0), .in1(andOp_33_in1), .out(andOp_33_out));

	wire [0:0] andOp_34_in0;
	wire [0:0] andOp_34_in1;
	wire [0:0] andOp_34_out;
	andOp #(.WIDTH(1)) andOp_34(.in0(andOp_34_in0), .in1(andOp_34_in1), .out(andOp_34_out));

	wire [0:0] notOp_35_in0;
	wire [0:0] notOp_35_out;
	notOp #(.WIDTH(1)) notOp_35(.in(notOp_35_in0), .out(notOp_35_out));

	wire [0:0] andOp_36_in0;
	wire [0:0] andOp_36_in1;
	wire [0:0] andOp_36_out;
	andOp #(.WIDTH(1)) andOp_36(.in0(andOp_36_in0), .in1(andOp_36_in1), .out(andOp_36_out));

	wire [0:0] notOp_37_in0;
	wire [0:0] notOp_37_out;
	notOp #(.WIDTH(1)) notOp_37(.in(notOp_37_in0), .out(notOp_37_out));

	wire [0:0] andOp_38_in0;
	wire [0:0] andOp_38_in1;
	wire [0:0] andOp_38_out;
	andOp #(.WIDTH(1)) andOp_38(.in0(andOp_38_in0), .in1(andOp_38_in1), .out(andOp_38_out));

	wire [0:0] notOp_39_in0;
	wire [0:0] notOp_39_out;
	notOp #(.WIDTH(1)) notOp_39(.in(notOp_39_in0), .out(notOp_39_out));

	wire [0:0] andOp_40_in0;
	wire [0:0] andOp_40_in1;
	wire [0:0] andOp_40_out;
	andOp #(.WIDTH(1)) andOp_40(.in0(andOp_40_in0), .in1(andOp_40_in1), .out(andOp_40_out));

	wire [0:0] notOp_41_in0;
	wire [0:0] notOp_41_out;
	notOp #(.WIDTH(1)) notOp_41(.in(notOp_41_in0), .out(notOp_41_out));

	wire [0:0] andOp_42_in0;
	wire [0:0] andOp_42_in1;
	wire [0:0] andOp_42_out;
	andOp #(.WIDTH(1)) andOp_42(.in0(andOp_42_in0), .in1(andOp_42_in1), .out(andOp_42_out));

	wire [0:0] notOp_43_in0;
	wire [0:0] notOp_43_out;
	notOp #(.WIDTH(1)) notOp_43(.in(notOp_43_in0), .out(notOp_43_out));

	wire [0:0] andOp_44_in0;
	wire [0:0] andOp_44_in1;
	wire [0:0] andOp_44_out;
	andOp #(.WIDTH(1)) andOp_44(.in0(andOp_44_in0), .in1(andOp_44_in1), .out(andOp_44_out));

	wire [0:0] notOp_45_in0;
	wire [0:0] notOp_45_out;
	notOp #(.WIDTH(1)) notOp_45(.in(notOp_45_in0), .out(notOp_45_out));

	wire [0:0] andOp_46_in0;
	wire [0:0] andOp_46_in1;
	wire [0:0] andOp_46_out;
	andOp #(.WIDTH(1)) andOp_46(.in0(andOp_46_in0), .in1(andOp_46_in1), .out(andOp_46_out));

	wire [0:0] andOp_47_in0;
	wire [0:0] andOp_47_in1;
	wire [0:0] andOp_47_out;
	andOp #(.WIDTH(1)) andOp_47(.in0(andOp_47_in0), .in1(andOp_47_in1), .out(andOp_47_out));

	wire [0:0] notOp_48_in0;
	wire [0:0] notOp_48_out;
	notOp #(.WIDTH(1)) notOp_48(.in(notOp_48_in0), .out(notOp_48_out));

	wire [0:0] andOp_49_in0;
	wire [0:0] andOp_49_in1;
	wire [0:0] andOp_49_out;
	andOp #(.WIDTH(1)) andOp_49(.in0(andOp_49_in0), .in1(andOp_49_in1), .out(andOp_49_out));

	wire [0:0] notOp_50_in0;
	wire [0:0] notOp_50_out;
	notOp #(.WIDTH(1)) notOp_50(.in(notOp_50_in0), .out(notOp_50_out));

	wire [0:0] andOp_51_in0;
	wire [0:0] andOp_51_in1;
	wire [0:0] andOp_51_out;
	andOp #(.WIDTH(1)) andOp_51(.in0(andOp_51_in0), .in1(andOp_51_in1), .out(andOp_51_out));

	wire [0:0] andOp_52_in0;
	wire [0:0] andOp_52_in1;
	wire [0:0] andOp_52_out;
	andOp #(.WIDTH(1)) andOp_52(.in0(andOp_52_in0), .in1(andOp_52_in1), .out(andOp_52_out));

	wire [0:0] notOp_53_in0;
	wire [0:0] notOp_53_out;
	notOp #(.WIDTH(1)) notOp_53(.in(notOp_53_in0), .out(notOp_53_out));

	wire [31:0] eq_54_in0;
	wire [31:0] eq_54_in1;
	wire [0:0] eq_54_out;
	eq #(.WIDTH(32)) eq_54(.in0(eq_54_in0), .in1(eq_54_in1), .out(eq_54_out));

	wire [31:0] eq_55_in0;
	wire [31:0] eq_55_in1;
	wire [0:0] eq_55_out;
	eq #(.WIDTH(32)) eq_55(.in0(eq_55_in0), .in1(eq_55_in1), .out(eq_55_out));

	wire [0:0] orOp_56_in0;
	wire [0:0] orOp_56_in1;
	wire [0:0] orOp_56_out;
	orOp #(.WIDTH(1)) orOp_56(.in0(orOp_56_in0), .in1(orOp_56_in1), .out(orOp_56_out));

	wire [31:0] eq_57_in0;
	wire [31:0] eq_57_in1;
	wire [0:0] eq_57_out;
	eq #(.WIDTH(32)) eq_57(.in0(eq_57_in0), .in1(eq_57_in1), .out(eq_57_out));

	wire [0:0] orOp_58_in0;
	wire [0:0] orOp_58_in1;
	wire [0:0] orOp_58_out;
	orOp #(.WIDTH(1)) orOp_58(.in0(orOp_58_in0), .in1(orOp_58_in1), .out(orOp_58_out));

	wire [31:0] eq_59_in0;
	wire [31:0] eq_59_in1;
	wire [0:0] eq_59_out;
	eq #(.WIDTH(32)) eq_59(.in0(eq_59_in0), .in1(eq_59_in1), .out(eq_59_out));

	wire [0:0] orOp_60_in0;
	wire [0:0] orOp_60_in1;
	wire [0:0] orOp_60_out;
	orOp #(.WIDTH(1)) orOp_60(.in0(orOp_60_in0), .in1(orOp_60_in1), .out(orOp_60_out));

	wire [31:0] eq_61_in0;
	wire [31:0] eq_61_in1;
	wire [0:0] eq_61_out;
	eq #(.WIDTH(32)) eq_61(.in0(eq_61_in0), .in1(eq_61_in1), .out(eq_61_out));

	wire [31:0] eq_62_in0;
	wire [31:0] eq_62_in1;
	wire [0:0] eq_62_out;
	eq #(.WIDTH(32)) eq_62(.in0(eq_62_in0), .in1(eq_62_in1), .out(eq_62_out));

	wire [31:0] eq_63_in0;
	wire [31:0] eq_63_in1;
	wire [0:0] eq_63_out;
	eq #(.WIDTH(32)) eq_63(.in0(eq_63_in0), .in1(eq_63_in1), .out(eq_63_out));

	wire [31:0] eq_64_in0;
	wire [31:0] eq_64_in1;
	wire [0:0] eq_64_out;
	eq #(.WIDTH(32)) eq_64(.in0(eq_64_in0), .in1(eq_64_in1), .out(eq_64_out));

	wire [0:0] orOp_65_in0;
	wire [0:0] orOp_65_in1;
	wire [0:0] orOp_65_out;
	orOp #(.WIDTH(1)) orOp_65(.in0(orOp_65_in0), .in1(orOp_65_in1), .out(orOp_65_out));

	wire [31:0] eq_66_in0;
	wire [31:0] eq_66_in1;
	wire [0:0] eq_66_out;
	eq #(.WIDTH(32)) eq_66(.in0(eq_66_in0), .in1(eq_66_in1), .out(eq_66_out));

	wire [0:0] orOp_67_in0;
	wire [0:0] orOp_67_in1;
	wire [0:0] orOp_67_out;
	orOp #(.WIDTH(1)) orOp_67(.in0(orOp_67_in0), .in1(orOp_67_in1), .out(orOp_67_out));

	wire [31:0] eq_68_in0;
	wire [31:0] eq_68_in1;
	wire [0:0] eq_68_out;
	eq #(.WIDTH(32)) eq_68(.in0(eq_68_in0), .in1(eq_68_in1), .out(eq_68_out));

	wire [0:0] orOp_69_in0;
	wire [0:0] orOp_69_in1;
	wire [0:0] orOp_69_out;
	orOp #(.WIDTH(1)) orOp_69(.in0(orOp_69_in0), .in1(orOp_69_in1), .out(orOp_69_out));

	wire [31:0] eq_70_in0;
	wire [31:0] eq_70_in1;
	wire [0:0] eq_70_out;
	eq #(.WIDTH(32)) eq_70(.in0(eq_70_in0), .in1(eq_70_in1), .out(eq_70_out));

	wire [0:0] orOp_71_in0;
	wire [0:0] orOp_71_in1;
	wire [0:0] orOp_71_out;
	orOp #(.WIDTH(1)) orOp_71(.in0(orOp_71_in0), .in1(orOp_71_in1), .out(orOp_71_out));

	wire [31:0] eq_72_in0;
	wire [31:0] eq_72_in1;
	wire [0:0] eq_72_out;
	eq #(.WIDTH(32)) eq_72(.in0(eq_72_in0), .in1(eq_72_in1), .out(eq_72_out));

	wire [31:0] eq_73_in0;
	wire [31:0] eq_73_in1;
	wire [0:0] eq_73_out;
	eq #(.WIDTH(32)) eq_73(.in0(eq_73_in0), .in1(eq_73_in1), .out(eq_73_out));

	wire [31:0] eq_74_in0;
	wire [31:0] eq_74_in1;
	wire [0:0] eq_74_out;
	eq #(.WIDTH(32)) eq_74(.in0(eq_74_in0), .in1(eq_74_in1), .out(eq_74_out));

	wire [0:0] notOp_75_in0;
	wire [0:0] notOp_75_out;
	notOp #(.WIDTH(1)) notOp_75(.in(notOp_75_in0), .out(notOp_75_out));

	wire [0:0] andOp_76_in0;
	wire [0:0] andOp_76_in1;
	wire [0:0] andOp_76_out;
	andOp #(.WIDTH(1)) andOp_76(.in0(andOp_76_in0), .in1(andOp_76_in1), .out(andOp_76_out));

	wire [31:0] eq_77_in0;
	wire [31:0] eq_77_in1;
	wire [0:0] eq_77_out;
	eq #(.WIDTH(32)) eq_77(.in0(eq_77_in0), .in1(eq_77_in1), .out(eq_77_out));

	wire [0:0] notOp_78_in0;
	wire [0:0] notOp_78_out;
	notOp #(.WIDTH(1)) notOp_78(.in(notOp_78_in0), .out(notOp_78_out));

	wire [0:0] andOp_79_in0;
	wire [0:0] andOp_79_in1;
	wire [0:0] andOp_79_out;
	andOp #(.WIDTH(1)) andOp_79(.in0(andOp_79_in0), .in1(andOp_79_in1), .out(andOp_79_out));

	wire [31:0] eq_80_in0;
	wire [31:0] eq_80_in1;
	wire [0:0] eq_80_out;
	eq #(.WIDTH(32)) eq_80(.in0(eq_80_in0), .in1(eq_80_in1), .out(eq_80_out));

	wire [0:0] notOp_81_in0;
	wire [0:0] notOp_81_out;
	notOp #(.WIDTH(1)) notOp_81(.in(notOp_81_in0), .out(notOp_81_out));

	wire [0:0] andOp_82_in0;
	wire [0:0] andOp_82_in1;
	wire [0:0] andOp_82_out;
	andOp #(.WIDTH(1)) andOp_82(.in0(andOp_82_in0), .in1(andOp_82_in1), .out(andOp_82_out));

	wire [31:0] eq_83_in0;
	wire [31:0] eq_83_in1;
	wire [0:0] eq_83_out;
	eq #(.WIDTH(32)) eq_83(.in0(eq_83_in0), .in1(eq_83_in1), .out(eq_83_out));

	wire [31:0] eq_84_in0;
	wire [31:0] eq_84_in1;
	wire [0:0] eq_84_out;
	eq #(.WIDTH(32)) eq_84(.in0(eq_84_in0), .in1(eq_84_in1), .out(eq_84_out));

	wire [31:0] eq_85_in0;
	wire [31:0] eq_85_in1;
	wire [0:0] eq_85_out;
	eq #(.WIDTH(32)) eq_85(.in0(eq_85_in0), .in1(eq_85_in1), .out(eq_85_out));

	wire [31:0] eq_86_in0;
	wire [31:0] eq_86_in1;
	wire [0:0] eq_86_out;
	eq #(.WIDTH(32)) eq_86(.in0(eq_86_in0), .in1(eq_86_in1), .out(eq_86_out));

	wire [0:0] notOp_87_in0;
	wire [0:0] notOp_87_out;
	notOp #(.WIDTH(1)) notOp_87(.in(notOp_87_in0), .out(notOp_87_out));

	wire [0:0] andOp_88_in0;
	wire [0:0] andOp_88_in1;
	wire [0:0] andOp_88_out;
	andOp #(.WIDTH(1)) andOp_88(.in0(andOp_88_in0), .in1(andOp_88_in1), .out(andOp_88_out));

	wire [31:0] eq_89_in0;
	wire [31:0] eq_89_in1;
	wire [0:0] eq_89_out;
	eq #(.WIDTH(32)) eq_89(.in0(eq_89_in0), .in1(eq_89_in1), .out(eq_89_out));

	wire [0:0] notOp_90_in0;
	wire [0:0] notOp_90_out;
	notOp #(.WIDTH(1)) notOp_90(.in(notOp_90_in0), .out(notOp_90_out));

	wire [0:0] andOp_91_in0;
	wire [0:0] andOp_91_in1;
	wire [0:0] andOp_91_out;
	andOp #(.WIDTH(1)) andOp_91(.in0(andOp_91_in0), .in1(andOp_91_in1), .out(andOp_91_out));

	wire [31:0] eq_92_in0;
	wire [31:0] eq_92_in1;
	wire [0:0] eq_92_out;
	eq #(.WIDTH(32)) eq_92(.in0(eq_92_in0), .in1(eq_92_in1), .out(eq_92_out));

	wire [0:0] notOp_93_in0;
	wire [0:0] notOp_93_out;
	notOp #(.WIDTH(1)) notOp_93(.in(notOp_93_in0), .out(notOp_93_out));

	wire [0:0] andOp_94_in0;
	wire [0:0] andOp_94_in1;
	wire [0:0] andOp_94_out;
	andOp #(.WIDTH(1)) andOp_94(.in0(andOp_94_in0), .in1(andOp_94_in1), .out(andOp_94_out));

	wire [31:0] eq_95_in0;
	wire [31:0] eq_95_in1;
	wire [0:0] eq_95_out;
	eq #(.WIDTH(32)) eq_95(.in0(eq_95_in0), .in1(eq_95_in1), .out(eq_95_out));

	wire [0:0] notOp_96_in0;
	wire [0:0] notOp_96_out;
	notOp #(.WIDTH(1)) notOp_96(.in(notOp_96_in0), .out(notOp_96_out));

	wire [0:0] andOp_97_in0;
	wire [0:0] andOp_97_in1;
	wire [0:0] andOp_97_out;
	andOp #(.WIDTH(1)) andOp_97(.in0(andOp_97_in0), .in1(andOp_97_in1), .out(andOp_97_out));

	wire [31:0] eq_98_in0;
	wire [31:0] eq_98_in1;
	wire [0:0] eq_98_out;
	eq #(.WIDTH(32)) eq_98(.in0(eq_98_in0), .in1(eq_98_in1), .out(eq_98_out));

	wire [0:0] andOp_99_in0;
	wire [0:0] andOp_99_in1;
	wire [0:0] andOp_99_out;
	andOp #(.WIDTH(1)) andOp_99(.in0(andOp_99_in0), .in1(andOp_99_in1), .out(andOp_99_out));

	wire [0:0] andOp_100_in0;
	wire [0:0] andOp_100_in1;
	wire [0:0] andOp_100_out;
	andOp #(.WIDTH(1)) andOp_100(.in0(andOp_100_in0), .in1(andOp_100_in1), .out(andOp_100_out));

	wire [0:0] andOp_101_in0;
	wire [0:0] andOp_101_in1;
	wire [0:0] andOp_101_out;
	andOp #(.WIDTH(1)) andOp_101(.in0(andOp_101_in0), .in1(andOp_101_in1), .out(andOp_101_out));

	wire [0:0] andOp_102_in0;
	wire [0:0] andOp_102_in1;
	wire [0:0] andOp_102_out;
	andOp #(.WIDTH(1)) andOp_102(.in0(andOp_102_in0), .in1(andOp_102_in1), .out(andOp_102_out));

	wire [31:0] concat_103_in0;
	wire [31:0] concat_103_in1;
	wire [63:0] concat_103_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_103(.in0(concat_103_in0), .in1(concat_103_in1), .out(concat_103_out));

	wire [31:0] concat_104_in0;
	wire [31:0] concat_104_in1;
	wire [63:0] concat_104_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_104(.in0(concat_104_in0), .in1(concat_104_in1), .out(concat_104_out));

	wire [0:0] andOp_105_in0;
	wire [0:0] andOp_105_in1;
	wire [0:0] andOp_105_out;
	andOp #(.WIDTH(1)) andOp_105(.in0(andOp_105_in0), .in1(andOp_105_in1), .out(andOp_105_out));

	wire [0:0] andOp_106_in0;
	wire [0:0] andOp_106_in1;
	wire [0:0] andOp_106_out;
	andOp #(.WIDTH(1)) andOp_106(.in0(andOp_106_in0), .in1(andOp_106_in1), .out(andOp_106_out));

	wire [0:0] andOp_107_in0;
	wire [0:0] andOp_107_in1;
	wire [0:0] andOp_107_out;
	andOp #(.WIDTH(1)) andOp_107(.in0(andOp_107_in0), .in1(andOp_107_in1), .out(andOp_107_out));

	wire [0:0] andOp_108_in0;
	wire [0:0] andOp_108_in1;
	wire [0:0] andOp_108_out;
	andOp #(.WIDTH(1)) andOp_108(.in0(andOp_108_in0), .in1(andOp_108_in1), .out(andOp_108_out));

	wire [0:0] andOp_109_in0;
	wire [0:0] andOp_109_in1;
	wire [0:0] andOp_109_out;
	andOp #(.WIDTH(1)) andOp_109(.in0(andOp_109_in0), .in1(andOp_109_in1), .out(andOp_109_out));

	wire [0:0] andOp_110_in0;
	wire [0:0] andOp_110_in1;
	wire [0:0] andOp_110_out;
	andOp #(.WIDTH(1)) andOp_110(.in0(andOp_110_in0), .in1(andOp_110_in1), .out(andOp_110_out));

	wire [0:0] andOp_111_in0;
	wire [0:0] andOp_111_in1;
	wire [0:0] andOp_111_out;
	andOp #(.WIDTH(1)) andOp_111(.in0(andOp_111_in0), .in1(andOp_111_in1), .out(andOp_111_out));

	wire [0:0] andOp_112_in0;
	wire [0:0] andOp_112_in1;
	wire [0:0] andOp_112_out;
	andOp #(.WIDTH(1)) andOp_112(.in0(andOp_112_in0), .in1(andOp_112_in1), .out(andOp_112_out));

	wire [0:0] andOp_113_in0;
	wire [0:0] andOp_113_in1;
	wire [0:0] andOp_113_out;
	andOp #(.WIDTH(1)) andOp_113(.in0(andOp_113_in0), .in1(andOp_113_in1), .out(andOp_113_out));

	wire [0:0] notOp_114_in0;
	wire [0:0] notOp_114_out;
	notOp #(.WIDTH(1)) notOp_114(.in(notOp_114_in0), .out(notOp_114_out));

	wire [0:0] andOp_115_in0;
	wire [0:0] andOp_115_in1;
	wire [0:0] andOp_115_out;
	andOp #(.WIDTH(1)) andOp_115(.in0(andOp_115_in0), .in1(andOp_115_in1), .out(andOp_115_out));

	wire [0:0] notOp_116_in0;
	wire [0:0] notOp_116_out;
	notOp #(.WIDTH(1)) notOp_116(.in(notOp_116_in0), .out(notOp_116_out));

	wire [0:0] andOp_117_in0;
	wire [0:0] andOp_117_in1;
	wire [0:0] andOp_117_out;
	andOp #(.WIDTH(1)) andOp_117(.in0(andOp_117_in0), .in1(andOp_117_in1), .out(andOp_117_out));

	wire [0:0] notOp_118_in0;
	wire [0:0] notOp_118_out;
	notOp #(.WIDTH(1)) notOp_118(.in(notOp_118_in0), .out(notOp_118_out));

	wire [0:0] andOp_119_in0;
	wire [0:0] andOp_119_in1;
	wire [0:0] andOp_119_out;
	andOp #(.WIDTH(1)) andOp_119(.in0(andOp_119_in0), .in1(andOp_119_in1), .out(andOp_119_out));

	wire [0:0] notOp_120_in0;
	wire [0:0] notOp_120_out;
	notOp #(.WIDTH(1)) notOp_120(.in(notOp_120_in0), .out(notOp_120_out));

	wire [0:0] andOp_121_in0;
	wire [0:0] andOp_121_in1;
	wire [0:0] andOp_121_out;
	andOp #(.WIDTH(1)) andOp_121(.in0(andOp_121_in0), .in1(andOp_121_in1), .out(andOp_121_out));

	wire [0:0] notOp_122_in0;
	wire [0:0] notOp_122_out;
	notOp #(.WIDTH(1)) notOp_122(.in(notOp_122_in0), .out(notOp_122_out));

	wire [0:0] andOp_123_in0;
	wire [0:0] andOp_123_in1;
	wire [0:0] andOp_123_out;
	andOp #(.WIDTH(1)) andOp_123(.in0(andOp_123_in0), .in1(andOp_123_in1), .out(andOp_123_out));

	wire [0:0] notOp_124_in0;
	wire [0:0] notOp_124_out;
	notOp #(.WIDTH(1)) notOp_124(.in(notOp_124_in0), .out(notOp_124_out));

	wire [0:0] andOp_125_in0;
	wire [0:0] andOp_125_in1;
	wire [0:0] andOp_125_out;
	andOp #(.WIDTH(1)) andOp_125(.in0(andOp_125_in0), .in1(andOp_125_in1), .out(andOp_125_out));

	wire [0:0] notOp_126_in0;
	wire [0:0] notOp_126_out;
	notOp #(.WIDTH(1)) notOp_126(.in(notOp_126_in0), .out(notOp_126_out));

	wire [0:0] andOp_127_in0;
	wire [0:0] andOp_127_in1;
	wire [0:0] andOp_127_out;
	andOp #(.WIDTH(1)) andOp_127(.in0(andOp_127_in0), .in1(andOp_127_in1), .out(andOp_127_out));

	wire [0:0] notOp_128_in0;
	wire [0:0] notOp_128_out;
	notOp #(.WIDTH(1)) notOp_128(.in(notOp_128_in0), .out(notOp_128_out));

	wire [0:0] andOp_129_in0;
	wire [0:0] andOp_129_in1;
	wire [0:0] andOp_129_out;
	andOp #(.WIDTH(1)) andOp_129(.in0(andOp_129_in0), .in1(andOp_129_in1), .out(andOp_129_out));

	wire [31:0] eq_130_in0;
	wire [31:0] eq_130_in1;
	wire [0:0] eq_130_out;
	eq #(.WIDTH(32)) eq_130(.in0(eq_130_in0), .in1(eq_130_in1), .out(eq_130_out));

	wire [31:0] eq_131_in0;
	wire [31:0] eq_131_in1;
	wire [0:0] eq_131_out;
	eq #(.WIDTH(32)) eq_131(.in0(eq_131_in0), .in1(eq_131_in1), .out(eq_131_out));

	wire [0:0] andOp_132_in0;
	wire [0:0] andOp_132_in1;
	wire [0:0] andOp_132_out;
	andOp #(.WIDTH(1)) andOp_132(.in0(andOp_132_in0), .in1(andOp_132_in1), .out(andOp_132_out));

	wire [31:0] eq_133_in0;
	wire [31:0] eq_133_in1;
	wire [0:0] eq_133_out;
	eq #(.WIDTH(32)) eq_133(.in0(eq_133_in0), .in1(eq_133_in1), .out(eq_133_out));

	wire [31:0] eq_134_in0;
	wire [31:0] eq_134_in1;
	wire [0:0] eq_134_out;
	eq #(.WIDTH(32)) eq_134(.in0(eq_134_in0), .in1(eq_134_in1), .out(eq_134_out));

	wire [31:0] eq_135_in0;
	wire [31:0] eq_135_in1;
	wire [0:0] eq_135_out;
	eq #(.WIDTH(32)) eq_135(.in0(eq_135_in0), .in1(eq_135_in1), .out(eq_135_out));

	wire [31:0] eq_136_in0;
	wire [31:0] eq_136_in1;
	wire [0:0] eq_136_out;
	eq #(.WIDTH(32)) eq_136(.in0(eq_136_in0), .in1(eq_136_in1), .out(eq_136_out));

	wire [0:0] andOp_137_in0;
	wire [0:0] andOp_137_in1;
	wire [0:0] andOp_137_out;
	andOp #(.WIDTH(1)) andOp_137(.in0(andOp_137_in0), .in1(andOp_137_in1), .out(andOp_137_out));

	wire [31:0] eq_138_in0;
	wire [31:0] eq_138_in1;
	wire [0:0] eq_138_out;
	eq #(.WIDTH(32)) eq_138(.in0(eq_138_in0), .in1(eq_138_in1), .out(eq_138_out));

	wire [31:0] eq_139_in0;
	wire [31:0] eq_139_in1;
	wire [0:0] eq_139_out;
	eq #(.WIDTH(32)) eq_139(.in0(eq_139_in0), .in1(eq_139_in1), .out(eq_139_out));

	wire [0:0] andOp_140_in0;
	wire [0:0] andOp_140_in1;
	wire [0:0] andOp_140_out;
	andOp #(.WIDTH(1)) andOp_140(.in0(andOp_140_in0), .in1(andOp_140_in1), .out(andOp_140_out));

	wire [31:0] eq_141_in0;
	wire [31:0] eq_141_in1;
	wire [0:0] eq_141_out;
	eq #(.WIDTH(32)) eq_141(.in0(eq_141_in0), .in1(eq_141_in1), .out(eq_141_out));

	wire [31:0] eq_142_in0;
	wire [31:0] eq_142_in1;
	wire [0:0] eq_142_out;
	eq #(.WIDTH(32)) eq_142(.in0(eq_142_in0), .in1(eq_142_in1), .out(eq_142_out));

	wire [0:0] notOp_143_in0;
	wire [0:0] notOp_143_out;
	notOp #(.WIDTH(1)) notOp_143(.in(notOp_143_in0), .out(notOp_143_out));

	wire [0:0] notOp_144_in0;
	wire [0:0] notOp_144_out;
	notOp #(.WIDTH(1)) notOp_144(.in(notOp_144_in0), .out(notOp_144_out));

	wire [0:0] andOp_145_in0;
	wire [0:0] andOp_145_in1;
	wire [0:0] andOp_145_out;
	andOp #(.WIDTH(1)) andOp_145(.in0(andOp_145_in0), .in1(andOp_145_in1), .out(andOp_145_out));

	wire [0:0] andOp_146_in0;
	wire [0:0] andOp_146_in1;
	wire [0:0] andOp_146_out;
	andOp #(.WIDTH(1)) andOp_146(.in0(andOp_146_in0), .in1(andOp_146_in1), .out(andOp_146_out));

	wire [0:0] andOp_147_in0;
	wire [0:0] andOp_147_in1;
	wire [0:0] andOp_147_out;
	andOp #(.WIDTH(1)) andOp_147(.in0(andOp_147_in0), .in1(andOp_147_in1), .out(andOp_147_out));

	// End Functional Units

	reg [31:0] data_store_0_0;
	reg [31:0] data_store_0_2;
	reg [31:0] data_store_1_4;
	reg [31:0] data_store_1_6;
	reg [31:0] data_store_2_11;
	reg [31:0] data_store_2_8;
	reg [31:0] data_store_2_9;
	reg [31:0] data_store_3_13;
	reg [31:0] data_store_3_15;
	reg [31:0] data_store_3_17;
	reg [31:0] data_store_4_19;
	reg [31:0] data_store_4_21;
	reg [31:0] global_state;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_3_last_state;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;
	reg [31:0] state_4_last_state;

	// controller for add_add6.add_add6_in0
	// controller for add_add6.add_add6_in1
	// Insensitive connections
	assign add_add6_in0 = phi_phi5_out;
	assign add_add6_in1 = 32'd1;
	// controller for andOp_100.andOp_100_in0
	// controller for andOp_100.andOp_100_in1
	// Insensitive connections
	assign andOp_100_in0 = bb_7_active_in_state_1_out_data;
	assign andOp_100_in1 = state_1_is_active;
	// controller for andOp_101.andOp_101_in0
	// controller for andOp_101.andOp_101_in1
	// Insensitive connections
	assign andOp_101_in0 = bb_7_active_in_state_2_out_data;
	assign andOp_101_in1 = state_2_is_active;
	// controller for andOp_102.andOp_102_in0
	// controller for andOp_102.andOp_102_in1
	// Insensitive connections
	assign andOp_102_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_102_in1 = state_0_is_active;
	// controller for andOp_105.andOp_105_in0
	// controller for andOp_105.andOp_105_in1
	// Insensitive connections
	assign andOp_105_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_105_in1 = state_0_is_active;
	// controller for andOp_106.andOp_106_in0
	// controller for andOp_106.andOp_106_in1
	// Insensitive connections
	assign andOp_106_in0 = bb_9_active_in_state_3_out_data;
	assign andOp_106_in1 = state_3_is_active;
	// controller for andOp_107.andOp_107_in0
	// controller for andOp_107.andOp_107_in1
	// Insensitive connections
	assign andOp_107_in0 = bb_10_active_in_state_4_out_data;
	assign andOp_107_in1 = state_4_is_active;
	// controller for andOp_108.andOp_108_in0
	// controller for andOp_108.andOp_108_in1
	// Insensitive connections
	assign andOp_108_in0 = bb_10_active_in_state_4_out_data;
	assign andOp_108_in1 = state_4_is_active;
	// controller for andOp_109.andOp_109_in0
	// controller for andOp_109.andOp_109_in1
	// Insensitive connections
	assign andOp_109_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_109_in1 = state_3_is_active;
	// controller for andOp_110.andOp_110_in0
	// controller for andOp_110.andOp_110_in1
	// Insensitive connections
	assign andOp_110_in0 = bb_3_active_in_state_4_out_data;
	assign andOp_110_in1 = state_4_is_active;
	// controller for andOp_111.andOp_111_in0
	// controller for andOp_111.andOp_111_in1
	// Insensitive connections
	assign andOp_111_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_111_in1 = state_4_is_active;
	// controller for andOp_112.andOp_112_in0
	// controller for andOp_112.andOp_112_in1
	// Insensitive connections
	assign andOp_112_in0 = bb_7_active_in_state_1_out_data;
	assign andOp_112_in1 = state_1_is_active;
	// controller for andOp_113.andOp_113_in0
	// controller for andOp_113.andOp_113_in1
	// Insensitive connections
	assign andOp_113_in0 = bb_4_active_in_state_4_out_data;
	assign andOp_113_in1 = state_4_is_active;
	// controller for andOp_115.andOp_115_in0
	// controller for andOp_115.andOp_115_in1
	// Insensitive connections
	assign andOp_115_in0 = notOp_114_out;
	assign andOp_115_in1 = 1'd1;
	// controller for andOp_117.andOp_117_in0
	// controller for andOp_117.andOp_117_in1
	// Insensitive connections
	assign andOp_117_in0 = notOp_116_out;
	assign andOp_117_in1 = andOp_115_out;
	// controller for andOp_119.andOp_119_in0
	// controller for andOp_119.andOp_119_in1
	// Insensitive connections
	assign andOp_119_in0 = notOp_118_out;
	assign andOp_119_in1 = 1'd1;
	// controller for andOp_121.andOp_121_in0
	// controller for andOp_121.andOp_121_in1
	// Insensitive connections
	assign andOp_121_in0 = notOp_120_out;
	assign andOp_121_in1 = 1'd1;
	// controller for andOp_123.andOp_123_in0
	// controller for andOp_123.andOp_123_in1
	// Insensitive connections
	assign andOp_123_in0 = notOp_122_out;
	assign andOp_123_in1 = 1'd1;
	// controller for andOp_125.andOp_125_in0
	// controller for andOp_125.andOp_125_in1
	// Insensitive connections
	assign andOp_125_in0 = notOp_124_out;
	assign andOp_125_in1 = andOp_123_out;
	// controller for andOp_127.andOp_127_in0
	// controller for andOp_127.andOp_127_in1
	// Insensitive connections
	assign andOp_127_in0 = notOp_126_out;
	assign andOp_127_in1 = 1'd1;
	// controller for andOp_129.andOp_129_in0
	// controller for andOp_129.andOp_129_in1
	// Insensitive connections
	assign andOp_129_in0 = notOp_128_out;
	assign andOp_129_in1 = andOp_127_out;
	// controller for andOp_132.andOp_132_in0
	// controller for andOp_132.andOp_132_in1
	// Insensitive connections
	assign andOp_132_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_132_in1 = state_0_is_active;
	// controller for andOp_137.andOp_137_in0
	// controller for andOp_137.andOp_137_in1
	// Insensitive connections
	assign andOp_137_in0 = bb_7_active_in_state_2_out_data;
	assign andOp_137_in1 = state_2_is_active;
	// controller for andOp_140.andOp_140_in0
	// controller for andOp_140.andOp_140_in1
	// Insensitive connections
	assign andOp_140_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_140_in1 = state_3_is_active;
	// controller for andOp_145.andOp_145_in0
	// controller for andOp_145.andOp_145_in1
	// Insensitive connections
	assign andOp_145_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_145_in1 = state_0_is_active;
	// controller for andOp_146.andOp_146_in0
	// controller for andOp_146.andOp_146_in1
	// Insensitive connections
	assign andOp_146_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_146_in1 = state_3_is_active;
	// controller for andOp_147.andOp_147_in0
	// controller for andOp_147.andOp_147_in1
	// Insensitive connections
	assign andOp_147_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_147_in1 = state_0_is_active;
	// controller for andOp_23.andOp_23_in0
	// controller for andOp_23.andOp_23_in1
	// Insensitive connections
	assign andOp_23_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_23_in1 = state_0_is_active;
	// controller for andOp_25.andOp_25_in0
	// controller for andOp_25.andOp_25_in1
	// Insensitive connections
	assign andOp_25_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_25_in1 = state_0_is_active;
	// controller for andOp_27.andOp_27_in0
	// controller for andOp_27.andOp_27_in1
	// Insensitive connections
	assign andOp_27_in0 = bb_5_active_in_state_0_out_data;
	assign andOp_27_in1 = state_0_is_active;
	// controller for andOp_29.andOp_29_in0
	// controller for andOp_29.andOp_29_in1
	// Insensitive connections
	assign andOp_29_in0 = bb_6_active_in_state_0_out_data;
	assign andOp_29_in1 = state_0_is_active;
	// controller for andOp_31.andOp_31_in0
	// controller for andOp_31.andOp_31_in1
	// Insensitive connections
	assign andOp_31_in0 = andOp_29_out;
	assign andOp_31_in1 = arg_0_read_ready;
	// controller for andOp_33.andOp_33_in0
	// controller for andOp_33.andOp_33_in1
	// Insensitive connections
	assign andOp_33_in0 = andOp_29_out;
	assign andOp_33_in1 = notOp_32_out;
	// controller for andOp_34.andOp_34_in0
	// controller for andOp_34.andOp_34_in1
	// Insensitive connections
	assign andOp_34_in0 = bb_7_active_in_state_2_out_data;
	assign andOp_34_in1 = state_2_is_active;
	// controller for andOp_36.andOp_36_in0
	// controller for andOp_36.andOp_36_in1
	// Insensitive connections
	assign andOp_36_in0 = bb_7_active_in_state_2_out_data;
	assign andOp_36_in1 = state_2_is_active;
	// controller for andOp_38.andOp_38_in0
	// controller for andOp_38.andOp_38_in1
	// Insensitive connections
	assign andOp_38_in0 = bb_2_active_in_state_3_out_data;
	assign andOp_38_in1 = state_3_is_active;
	// controller for andOp_40.andOp_40_in0
	// controller for andOp_40.andOp_40_in1
	// Insensitive connections
	assign andOp_40_in0 = bb_8_active_in_state_3_out_data;
	assign andOp_40_in1 = state_3_is_active;
	// controller for andOp_42.andOp_42_in0
	// controller for andOp_42.andOp_42_in1
	// Insensitive connections
	assign andOp_42_in0 = bb_9_active_in_state_3_out_data;
	assign andOp_42_in1 = state_3_is_active;
	// controller for andOp_44.andOp_44_in0
	// controller for andOp_44.andOp_44_in1
	// Insensitive connections
	assign andOp_44_in0 = andOp_42_out;
	assign andOp_44_in1 = arg_1_write_ready;
	// controller for andOp_46.andOp_46_in0
	// controller for andOp_46.andOp_46_in1
	// Insensitive connections
	assign andOp_46_in0 = andOp_42_out;
	assign andOp_46_in1 = notOp_45_out;
	// controller for andOp_47.andOp_47_in0
	// controller for andOp_47.andOp_47_in1
	// Insensitive connections
	assign andOp_47_in0 = bb_3_active_in_state_4_out_data;
	assign andOp_47_in1 = state_4_is_active;
	// controller for andOp_49.andOp_49_in0
	// controller for andOp_49.andOp_49_in1
	// Insensitive connections
	assign andOp_49_in0 = andOp_47_out;
	assign andOp_49_in1 = icmp_icmp18_out;
	// controller for andOp_51.andOp_51_in0
	// controller for andOp_51.andOp_51_in1
	// Insensitive connections
	assign andOp_51_in0 = andOp_47_out;
	assign andOp_51_in1 = notOp_50_out;
	// controller for andOp_52.andOp_52_in0
	// controller for andOp_52.andOp_52_in1
	// Insensitive connections
	assign andOp_52_in0 = bb_10_active_in_state_4_out_data;
	assign andOp_52_in1 = state_4_is_active;
	// controller for andOp_76.andOp_76_in0
	// controller for andOp_76.andOp_76_in1
	// Insensitive connections
	assign andOp_76_in0 = notOp_75_out;
	assign andOp_76_in1 = andOp_23_out;
	// controller for andOp_79.andOp_79_in0
	// controller for andOp_79.andOp_79_in1
	// Insensitive connections
	assign andOp_79_in0 = notOp_78_out;
	assign andOp_79_in1 = andOp_25_out;
	// controller for andOp_82.andOp_82_in0
	// controller for andOp_82.andOp_82_in1
	// Insensitive connections
	assign andOp_82_in0 = notOp_81_out;
	assign andOp_82_in1 = andOp_27_out;
	// controller for andOp_88.andOp_88_in0
	// controller for andOp_88.andOp_88_in1
	// Insensitive connections
	assign andOp_88_in0 = notOp_87_out;
	assign andOp_88_in1 = andOp_38_out;
	// controller for andOp_91.andOp_91_in0
	// controller for andOp_91.andOp_91_in1
	// Insensitive connections
	assign andOp_91_in0 = notOp_90_out;
	assign andOp_91_in1 = andOp_40_out;
	// controller for andOp_94.andOp_94_in0
	// controller for andOp_94.andOp_94_in1
	// Insensitive connections
	assign andOp_94_in0 = notOp_93_out;
	assign andOp_94_in1 = andOp_51_out;
	// controller for andOp_97.andOp_97_in0
	// controller for andOp_97.andOp_97_in1
	// Insensitive connections
	assign andOp_97_in0 = notOp_96_out;
	assign andOp_97_in1 = andOp_52_out;
	// controller for andOp_99.andOp_99_in0
	// controller for andOp_99.andOp_99_in1
	// Insensitive connections
	assign andOp_99_in0 = bb_6_active_in_state_0_out_data;
	assign andOp_99_in1 = state_0_is_active;
	// controller for arg_0.arg_0_read_valid_reg
	always @(*) begin
		if (andOp_100_out) begin 
			arg_0_read_valid_reg = -(1'd1);
		end else begin
			arg_0_read_valid_reg = 0;
		end
	end
	// controller for arg_1.arg_1_in_data_reg
	always @(*) begin
		if (andOp_108_out) begin 
			arg_1_in_data_reg = data_in_4_22_out_data;
		end else begin
			arg_1_in_data_reg = 0;
		end
	end
	// controller for arg_1.arg_1_write_valid_reg
	always @(*) begin
		if (andOp_107_out) begin 
			arg_1_write_valid_reg = -(1'd1);
		end else begin
			arg_1_write_valid_reg = 0;
		end
	end
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_54_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_73_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_4.bb_10_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_4_in_data = eq_72_out;
		end else begin
			bb_10_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_4.bb_10_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_98_out) begin 
			bb_10_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_0.bb_1_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_0_in_data = orOp_56_out;
		end else begin
			bb_1_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_0.bb_1_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_76_out) begin 
			bb_1_predecessor_in_state_0_in_data = 32'd0;
		end else if (eq_74_out) begin 
			bb_1_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_3.bb_2_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_3_in_data = eq_63_out;
		end else begin
			bb_2_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_3.bb_2_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_85_out) begin 
			bb_2_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_4.bb_3_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_4_in_data = orOp_71_out;
		end else begin
			bb_3_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_4.bb_3_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_97_out) begin 
			bb_3_predecessor_in_state_4_in_data = 32'd10;
		end else if (eq_95_out) begin 
			bb_3_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_4.bb_4_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_4_in_data = orOp_69_out;
		end else begin
			bb_4_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_4.bb_4_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_94_out) begin 
			bb_4_predecessor_in_state_4_in_data = 32'd3;
		end else if (eq_92_out) begin 
			bb_4_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_5_active_in_state_0.bb_5_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_5_active_in_state_0_in_data = orOp_58_out;
		end else begin
			bb_5_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_5_predecessor_in_state_0.bb_5_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_79_out) begin 
			bb_5_predecessor_in_state_0_in_data = 32'd1;
		end else if (eq_77_out) begin 
			bb_5_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_5_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_6_active_in_state_0.bb_6_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_6_active_in_state_0_in_data = orOp_60_out;
		end else begin
			bb_6_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_6_predecessor_in_state_0.bb_6_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_82_out) begin 
			bb_6_predecessor_in_state_0_in_data = 32'd5;
		end else if (eq_80_out) begin 
			bb_6_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_6_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_7_active_in_state_1.bb_7_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_7_active_in_state_1_in_data = eq_61_out;
		end else begin
			bb_7_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_7_active_in_state_2.bb_7_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_7_active_in_state_2_in_data = eq_62_out;
		end else begin
			bb_7_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_7_predecessor_in_state_1.bb_7_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_83_out) begin 
			bb_7_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_7_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_7_predecessor_in_state_2.bb_7_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_84_out) begin 
			bb_7_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_7_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_8_active_in_state_3.bb_8_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_state_3_in_data = orOp_65_out;
		end else begin
			bb_8_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_8_predecessor_in_state_3.bb_8_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_88_out) begin 
			bb_8_predecessor_in_state_3_in_data = 32'd2;
		end else if (eq_86_out) begin 
			bb_8_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_8_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_9_active_in_state_3.bb_9_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_9_active_in_state_3_in_data = orOp_67_out;
		end else begin
			bb_9_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_9_predecessor_in_state_3.bb_9_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_91_out) begin 
			bb_9_predecessor_in_state_3_in_data = 32'd8;
		end else if (eq_89_out) begin 
			bb_9_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_9_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_23_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_24_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_4.br_10_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_52_out) begin 
			br_10_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_53_out) begin 
			br_10_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_1_happened_in_state_0.br_1_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_25_out) begin 
			br_1_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_26_out) begin 
			br_1_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_1_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_2_happened_in_state_3.br_2_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_38_out) begin 
			br_2_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_39_out) begin 
			br_2_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_2_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_4.br_3_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_47_out) begin 
			br_3_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_48_out) begin 
			br_3_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_5_happened_in_state_0.br_5_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_27_out) begin 
			br_5_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_28_out) begin 
			br_5_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_5_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_6_happened_in_state_0.br_6_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_29_out) begin 
			br_6_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_30_out) begin 
			br_6_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_6_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_7_happened_in_state_1.br_7_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_34_out) begin 
			br_7_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_35_out) begin 
			br_7_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_7_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_7_happened_in_state_2.br_7_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_36_out) begin 
			br_7_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_37_out) begin 
			br_7_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_7_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_8_happened_in_state_3.br_8_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_40_out) begin 
			br_8_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_41_out) begin 
			br_8_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_8_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_9_happened_in_state_3.br_9_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_42_out) begin 
			br_9_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_43_out) begin 
			br_9_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_9_happened_in_state_3_in_data = 0;
		end
	end
	// controller for concat_103.concat_103_in0
	// controller for concat_103.concat_103_in1
	// Insensitive connections
	assign concat_103_in0 = data_in_0_1_out_data;
	assign concat_103_in1 = 32'd0;
	// controller for concat_104.concat_104_in0
	// controller for concat_104.concat_104_in1
	// Insensitive connections
	assign concat_104_in0 = 32'd3;
	assign concat_104_in1 = 32'd0;
	// controller for data_in_0_1.data_in_0_1_in_data
	always @(*) begin
		if (eq_130_out) begin 
			data_in_0_1_in_data = data_store_0_0;
		end else if (eq_131_out) begin 
			data_in_0_1_in_data = data_store_4_19;
		end else begin
			data_in_0_1_in_data = 0;
		end
	end
	// controller for data_in_0_3.data_in_0_3_in_data
	always @(*) begin
		if (eq_130_out) begin 
			data_in_0_3_in_data = data_store_0_2;
		end else if (eq_131_out) begin 
			data_in_0_3_in_data = data_store_4_21;
		end else begin
			data_in_0_3_in_data = 0;
		end
	end
	// controller for data_in_1_5.data_in_1_5_in_data
	always @(*) begin
		if (eq_133_out) begin 
			data_in_1_5_in_data = data_store_0_0;
		end else if (eq_134_out) begin 
			data_in_1_5_in_data = data_store_1_4;
		end else begin
			data_in_1_5_in_data = 0;
		end
	end
	// controller for data_in_1_7.data_in_1_7_in_data
	always @(*) begin
		if (eq_133_out) begin 
			data_in_1_7_in_data = data_store_0_2;
		end else if (eq_134_out) begin 
			data_in_1_7_in_data = data_store_1_6;
		end else begin
			data_in_1_7_in_data = 0;
		end
	end
	// controller for data_in_2_10.data_in_2_10_in_data
	always @(*) begin
		if (eq_135_out) begin 
			data_in_2_10_in_data = data_store_1_4;
		end else if (eq_136_out) begin 
			data_in_2_10_in_data = data_store_2_9;
		end else begin
			data_in_2_10_in_data = 0;
		end
	end
	// controller for data_in_2_12.data_in_2_12_in_data
	always @(*) begin
		if (eq_135_out) begin 
			data_in_2_12_in_data = data_store_1_6;
		end else if (eq_136_out) begin 
			data_in_2_12_in_data = data_store_2_11;
		end else begin
			data_in_2_12_in_data = 0;
		end
	end
	// controller for data_in_3_14.data_in_3_14_in_data
	always @(*) begin
		if (eq_138_out) begin 
			data_in_3_14_in_data = data_store_2_8;
		end else if (eq_139_out) begin 
			data_in_3_14_in_data = data_store_3_13;
		end else begin
			data_in_3_14_in_data = 0;
		end
	end
	// controller for data_in_3_16.data_in_3_16_in_data
	always @(*) begin
		if (eq_138_out) begin 
			data_in_3_16_in_data = data_store_2_9;
		end else if (eq_139_out) begin 
			data_in_3_16_in_data = data_store_3_15;
		end else begin
			data_in_3_16_in_data = 0;
		end
	end
	// controller for data_in_3_18.data_in_3_18_in_data
	always @(*) begin
		if (eq_138_out) begin 
			data_in_3_18_in_data = data_store_2_11;
		end else if (eq_139_out) begin 
			data_in_3_18_in_data = data_store_3_17;
		end else begin
			data_in_3_18_in_data = 0;
		end
	end
	// controller for data_in_4_20.data_in_4_20_in_data
	always @(*) begin
		if (eq_141_out) begin 
			data_in_4_20_in_data = data_store_3_15;
		end else if (eq_142_out) begin 
			data_in_4_20_in_data = data_store_4_19;
		end else begin
			data_in_4_20_in_data = 0;
		end
	end
	// controller for data_in_4_22.data_in_4_22_in_data
	always @(*) begin
		if (eq_141_out) begin 
			data_in_4_22_in_data = data_store_3_17;
		end else if (eq_142_out) begin 
			data_in_4_22_in_data = data_store_4_21;
		end else begin
			data_in_4_22_in_data = 0;
		end
	end
	// controller for eq_130.eq_130_in0
	// controller for eq_130.eq_130_in1
	// Insensitive connections
	assign eq_130_in0 = 32'd0;
	assign eq_130_in1 = state_0_last_state;
	// controller for eq_131.eq_131_in0
	// controller for eq_131.eq_131_in1
	// Insensitive connections
	assign eq_131_in0 = 32'd4;
	assign eq_131_in1 = state_0_last_state;
	// controller for eq_133.eq_133_in0
	// controller for eq_133.eq_133_in1
	// Insensitive connections
	assign eq_133_in0 = 32'd0;
	assign eq_133_in1 = state_1_last_state;
	// controller for eq_134.eq_134_in0
	// controller for eq_134.eq_134_in1
	// Insensitive connections
	assign eq_134_in0 = 32'd1;
	assign eq_134_in1 = state_1_last_state;
	// controller for eq_135.eq_135_in0
	// controller for eq_135.eq_135_in1
	// Insensitive connections
	assign eq_135_in0 = 32'd1;
	assign eq_135_in1 = state_2_last_state;
	// controller for eq_136.eq_136_in0
	// controller for eq_136.eq_136_in1
	// Insensitive connections
	assign eq_136_in0 = 32'd2;
	assign eq_136_in1 = state_2_last_state;
	// controller for eq_138.eq_138_in0
	// controller for eq_138.eq_138_in1
	// Insensitive connections
	assign eq_138_in0 = 32'd2;
	assign eq_138_in1 = state_3_last_state;
	// controller for eq_139.eq_139_in0
	// controller for eq_139.eq_139_in1
	// Insensitive connections
	assign eq_139_in0 = 32'd3;
	assign eq_139_in1 = state_3_last_state;
	// controller for eq_141.eq_141_in0
	// controller for eq_141.eq_141_in1
	// Insensitive connections
	assign eq_141_in0 = 32'd3;
	assign eq_141_in1 = state_4_last_state;
	// controller for eq_142.eq_142_in0
	// controller for eq_142.eq_142_in1
	// Insensitive connections
	assign eq_142_in0 = 32'd4;
	assign eq_142_in1 = state_4_last_state;
	// controller for eq_54.eq_54_in0
	// controller for eq_54.eq_54_in1
	// Insensitive connections
	assign eq_54_in0 = 32'd0;
	assign eq_54_in1 = state_0_entry_BB_reg;
	// controller for eq_55.eq_55_in0
	// controller for eq_55.eq_55_in1
	// Insensitive connections
	assign eq_55_in0 = 32'd1;
	assign eq_55_in1 = state_0_entry_BB_reg;
	// controller for eq_57.eq_57_in0
	// controller for eq_57.eq_57_in1
	// Insensitive connections
	assign eq_57_in0 = 32'd5;
	assign eq_57_in1 = state_0_entry_BB_reg;
	// controller for eq_59.eq_59_in0
	// controller for eq_59.eq_59_in1
	// Insensitive connections
	assign eq_59_in0 = 32'd6;
	assign eq_59_in1 = state_0_entry_BB_reg;
	// controller for eq_61.eq_61_in0
	// controller for eq_61.eq_61_in1
	// Insensitive connections
	assign eq_61_in0 = 32'd7;
	assign eq_61_in1 = state_1_entry_BB_reg;
	// controller for eq_62.eq_62_in0
	// controller for eq_62.eq_62_in1
	// Insensitive connections
	assign eq_62_in0 = 32'd7;
	assign eq_62_in1 = state_2_entry_BB_reg;
	// controller for eq_63.eq_63_in0
	// controller for eq_63.eq_63_in1
	// Insensitive connections
	assign eq_63_in0 = 32'd2;
	assign eq_63_in1 = state_3_entry_BB_reg;
	// controller for eq_64.eq_64_in0
	// controller for eq_64.eq_64_in1
	// Insensitive connections
	assign eq_64_in0 = 32'd8;
	assign eq_64_in1 = state_3_entry_BB_reg;
	// controller for eq_66.eq_66_in0
	// controller for eq_66.eq_66_in1
	// Insensitive connections
	assign eq_66_in0 = 32'd9;
	assign eq_66_in1 = state_3_entry_BB_reg;
	// controller for eq_68.eq_68_in0
	// controller for eq_68.eq_68_in1
	// Insensitive connections
	assign eq_68_in0 = 32'd4;
	assign eq_68_in1 = state_4_entry_BB_reg;
	// controller for eq_70.eq_70_in0
	// controller for eq_70.eq_70_in1
	// Insensitive connections
	assign eq_70_in0 = 32'd3;
	assign eq_70_in1 = state_4_entry_BB_reg;
	// controller for eq_72.eq_72_in0
	// controller for eq_72.eq_72_in1
	// Insensitive connections
	assign eq_72_in0 = 32'd10;
	assign eq_72_in1 = state_4_entry_BB_reg;
	// controller for eq_73.eq_73_in0
	// controller for eq_73.eq_73_in1
	// Insensitive connections
	assign eq_73_in0 = 32'd0;
	assign eq_73_in1 = state_0_entry_BB_reg;
	// controller for eq_74.eq_74_in0
	// controller for eq_74.eq_74_in1
	// Insensitive connections
	assign eq_74_in0 = 32'd1;
	assign eq_74_in1 = state_0_entry_BB_reg;
	// controller for eq_77.eq_77_in0
	// controller for eq_77.eq_77_in1
	// Insensitive connections
	assign eq_77_in0 = 32'd5;
	assign eq_77_in1 = state_0_entry_BB_reg;
	// controller for eq_80.eq_80_in0
	// controller for eq_80.eq_80_in1
	// Insensitive connections
	assign eq_80_in0 = 32'd6;
	assign eq_80_in1 = state_0_entry_BB_reg;
	// controller for eq_83.eq_83_in0
	// controller for eq_83.eq_83_in1
	// Insensitive connections
	assign eq_83_in0 = 32'd7;
	assign eq_83_in1 = state_1_entry_BB_reg;
	// controller for eq_84.eq_84_in0
	// controller for eq_84.eq_84_in1
	// Insensitive connections
	assign eq_84_in0 = 32'd7;
	assign eq_84_in1 = state_2_entry_BB_reg;
	// controller for eq_85.eq_85_in0
	// controller for eq_85.eq_85_in1
	// Insensitive connections
	assign eq_85_in0 = 32'd2;
	assign eq_85_in1 = state_3_entry_BB_reg;
	// controller for eq_86.eq_86_in0
	// controller for eq_86.eq_86_in1
	// Insensitive connections
	assign eq_86_in0 = 32'd8;
	assign eq_86_in1 = state_3_entry_BB_reg;
	// controller for eq_89.eq_89_in0
	// controller for eq_89.eq_89_in1
	// Insensitive connections
	assign eq_89_in0 = 32'd9;
	assign eq_89_in1 = state_3_entry_BB_reg;
	// controller for eq_92.eq_92_in0
	// controller for eq_92.eq_92_in1
	// Insensitive connections
	assign eq_92_in0 = 32'd4;
	assign eq_92_in1 = state_4_entry_BB_reg;
	// controller for eq_95.eq_95_in0
	// controller for eq_95.eq_95_in1
	// Insensitive connections
	assign eq_95_in0 = 32'd3;
	assign eq_95_in1 = state_4_entry_BB_reg;
	// controller for eq_98.eq_98_in0
	// controller for eq_98.eq_98_in1
	// Insensitive connections
	assign eq_98_in0 = 32'd10;
	assign eq_98_in1 = state_4_entry_BB_reg;
	// controller for icmp_icmp18.icmp_icmp18_in0
	// controller for icmp_icmp18.icmp_icmp18_in1
	// Insensitive connections
	assign icmp_icmp18_in0 = data_in_4_20_out_data;
	assign icmp_icmp18_in1 = 32'd15;
	// controller for mul_mul14.mul_mul14_in0
	// controller for mul_mul14.mul_mul14_in1
	// Insensitive connections
	assign mul_mul14_in0 = 32'd2;
	assign mul_mul14_in1 = data_in_3_14_out_data;
	// controller for notOp_114.notOp_114_in0
	// Insensitive connections
	assign notOp_114_in0 = andOp_33_out;
	// controller for notOp_116.notOp_116_in0
	// Insensitive connections
	assign notOp_116_in0 = andOp_49_out;
	// controller for notOp_118.notOp_118_in0
	// Insensitive connections
	assign notOp_118_in0 = andOp_31_out;
	// controller for notOp_120.notOp_120_in0
	// Insensitive connections
	assign notOp_120_in0 = andOp_112_out;
	// controller for notOp_122.notOp_122_in0
	// Insensitive connections
	assign notOp_122_in0 = andOp_34_out;
	// controller for notOp_124.notOp_124_in0
	// Insensitive connections
	assign notOp_124_in0 = andOp_46_out;
	// controller for notOp_126.notOp_126_in0
	// Insensitive connections
	assign notOp_126_in0 = andOp_113_out;
	// controller for notOp_128.notOp_128_in0
	// Insensitive connections
	assign notOp_128_in0 = andOp_44_out;
	// controller for notOp_143.notOp_143_in0
	// Insensitive connections
	assign notOp_143_in0 = state_4_is_active;
	// controller for notOp_144.notOp_144_in0
	// Insensitive connections
	assign notOp_144_in0 = state_4_is_active;
	// controller for notOp_24.notOp_24_in0
	// Insensitive connections
	assign notOp_24_in0 = andOp_23_out;
	// controller for notOp_26.notOp_26_in0
	// Insensitive connections
	assign notOp_26_in0 = andOp_25_out;
	// controller for notOp_28.notOp_28_in0
	// Insensitive connections
	assign notOp_28_in0 = andOp_27_out;
	// controller for notOp_30.notOp_30_in0
	// Insensitive connections
	assign notOp_30_in0 = andOp_29_out;
	// controller for notOp_32.notOp_32_in0
	// Insensitive connections
	assign notOp_32_in0 = arg_0_read_ready;
	// controller for notOp_35.notOp_35_in0
	// Insensitive connections
	assign notOp_35_in0 = andOp_34_out;
	// controller for notOp_37.notOp_37_in0
	// Insensitive connections
	assign notOp_37_in0 = andOp_36_out;
	// controller for notOp_39.notOp_39_in0
	// Insensitive connections
	assign notOp_39_in0 = andOp_38_out;
	// controller for notOp_41.notOp_41_in0
	// Insensitive connections
	assign notOp_41_in0 = andOp_40_out;
	// controller for notOp_43.notOp_43_in0
	// Insensitive connections
	assign notOp_43_in0 = andOp_42_out;
	// controller for notOp_45.notOp_45_in0
	// Insensitive connections
	assign notOp_45_in0 = arg_1_write_ready;
	// controller for notOp_48.notOp_48_in0
	// Insensitive connections
	assign notOp_48_in0 = andOp_47_out;
	// controller for notOp_50.notOp_50_in0
	// Insensitive connections
	assign notOp_50_in0 = icmp_icmp18_out;
	// controller for notOp_53.notOp_53_in0
	// Insensitive connections
	assign notOp_53_in0 = andOp_52_out;
	// controller for notOp_75.notOp_75_in0
	// Insensitive connections
	assign notOp_75_in0 = eq_74_out;
	// controller for notOp_78.notOp_78_in0
	// Insensitive connections
	assign notOp_78_in0 = eq_77_out;
	// controller for notOp_81.notOp_81_in0
	// Insensitive connections
	assign notOp_81_in0 = eq_80_out;
	// controller for notOp_87.notOp_87_in0
	// Insensitive connections
	assign notOp_87_in0 = eq_86_out;
	// controller for notOp_90.notOp_90_in0
	// Insensitive connections
	assign notOp_90_in0 = eq_89_out;
	// controller for notOp_93.notOp_93_in0
	// Insensitive connections
	assign notOp_93_in0 = eq_92_out;
	// controller for notOp_96.notOp_96_in0
	// Insensitive connections
	assign notOp_96_in0 = eq_95_out;
	// controller for orOp_56.orOp_56_in0
	// controller for orOp_56.orOp_56_in1
	// Insensitive connections
	assign orOp_56_in0 = eq_55_out;
	assign orOp_56_in1 = andOp_23_out;
	// controller for orOp_58.orOp_58_in0
	// controller for orOp_58.orOp_58_in1
	// Insensitive connections
	assign orOp_58_in0 = eq_57_out;
	assign orOp_58_in1 = andOp_25_out;
	// controller for orOp_60.orOp_60_in0
	// controller for orOp_60.orOp_60_in1
	// Insensitive connections
	assign orOp_60_in0 = eq_59_out;
	assign orOp_60_in1 = andOp_27_out;
	// controller for orOp_65.orOp_65_in0
	// controller for orOp_65.orOp_65_in1
	// Insensitive connections
	assign orOp_65_in0 = eq_64_out;
	assign orOp_65_in1 = andOp_38_out;
	// controller for orOp_67.orOp_67_in0
	// controller for orOp_67.orOp_67_in1
	// Insensitive connections
	assign orOp_67_in0 = eq_66_out;
	assign orOp_67_in1 = andOp_40_out;
	// controller for orOp_69.orOp_69_in0
	// controller for orOp_69.orOp_69_in1
	// Insensitive connections
	assign orOp_69_in0 = eq_68_out;
	assign orOp_69_in1 = andOp_51_out;
	// controller for orOp_71.orOp_71_in0
	// controller for orOp_71.orOp_71_in1
	// Insensitive connections
	assign orOp_71_in0 = eq_70_out;
	assign orOp_71_in1 = andOp_52_out;
	// controller for phi_phi5.phi_phi5_in
	// controller for phi_phi5.phi_phi5_last_block
	// controller for phi_phi5.phi_phi5_s
	// Insensitive connections
	assign phi_phi5_in = concat_103_out;
	assign phi_phi5_last_block = bb_1_predecessor_in_state_0_out_data;
	assign phi_phi5_s = concat_104_out;
	// controller for ret20.valid_reg
	always @(*) begin
		if (andOp_111_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			data_store_0_0 <= 0;
		end else begin
			if (andOp_132_out) begin
				data_store_0_0 <= add_add6_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_2 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_2 <= data_in_0_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_4 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_4 <= data_in_1_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_6 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_6 <= data_in_1_7_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_11 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_11 <= data_in_2_12_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_8 <= 0;
		end else begin
			if (andOp_137_out) begin
				data_store_2_8 <= arg_0_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_9 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_9 <= data_in_2_10_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_13 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_13 <= data_in_3_14_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_15 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_15 <= data_in_3_16_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_17 <= 0;
		end else begin
			if (andOp_140_out) begin
				data_store_3_17 <= mul_mul14_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_19 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_19 <= data_in_4_20_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_21 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_21 <= data_in_4_22_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_112_out) begin
				global_state <= 32'd2;
			end
			if (andOp_113_out) begin
				global_state <= 32'd4;
			end
			if (andOp_31_out) begin
				global_state <= 32'd1;
			end
			if (andOp_33_out) begin
				global_state <= 32'd0;
			end
			if (andOp_34_out) begin
				global_state <= 32'd3;
			end
			if (andOp_44_out) begin
				global_state <= 32'd4;
			end
			if (andOp_46_out) begin
				global_state <= 32'd3;
			end
			if (andOp_49_out) begin
				global_state <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
			if (andOp_33_out) begin
				state_0_entry_BB_reg <= 32'd6;
			end
			if (andOp_49_out) begin
				state_0_entry_BB_reg <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (andOp_117_out) begin
				state_0_is_active <= 1'd0;
			end
			if (andOp_33_out) begin
				state_0_is_active <= 1'd1;
			end
			if (andOp_49_out) begin
				state_0_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
			if (andOp_33_out) begin
				state_0_last_BB_reg <= 32'd6;
			end
			if (andOp_49_out) begin
				state_0_last_BB_reg <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
			if (andOp_33_out) begin
				state_0_last_state <= 32'd0;
			end
			if (andOp_49_out) begin
				state_0_last_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_31_out) begin
				state_1_entry_BB_reg <= 32'd7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_119_out) begin
				state_1_is_active <= 1'd0;
			end
			if (andOp_31_out) begin
				state_1_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_31_out) begin
				state_1_last_BB_reg <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_31_out) begin
				state_1_last_state <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_112_out) begin
				state_2_entry_BB_reg <= 32'd7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_112_out) begin
				state_2_is_active <= 1'd1;
			end
			if (andOp_121_out) begin
				state_2_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_112_out) begin
				state_2_last_BB_reg <= bb_7_predecessor_in_state_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_112_out) begin
				state_2_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_34_out) begin
				state_3_entry_BB_reg <= 32'd2;
			end
			if (andOp_46_out) begin
				state_3_entry_BB_reg <= 32'd9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_125_out) begin
				state_3_is_active <= 1'd0;
			end
			if (andOp_34_out) begin
				state_3_is_active <= 1'd1;
			end
			if (andOp_46_out) begin
				state_3_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_34_out) begin
				state_3_last_BB_reg <= 32'd7;
			end
			if (andOp_46_out) begin
				state_3_last_BB_reg <= 32'd9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_state <= 0;
		end else begin
			if (andOp_34_out) begin
				state_3_last_state <= 32'd2;
			end
			if (andOp_46_out) begin
				state_3_last_state <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_113_out) begin
				state_4_entry_BB_reg <= 32'd4;
			end
			if (andOp_44_out) begin
				state_4_entry_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_113_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_129_out) begin
				state_4_is_active <= 1'd0;
			end
			if (andOp_44_out) begin
				state_4_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_113_out) begin
				state_4_last_BB_reg <= bb_4_predecessor_in_state_4_out_data;
			end
			if (andOp_44_out) begin
				state_4_last_BB_reg <= 32'd9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_state <= 0;
		end else begin
			if (andOp_113_out) begin
				state_4_last_state <= 32'd4;
			end
			if (andOp_44_out) begin
				state_4_last_state <= 32'd3;
			end
		end
	end

endmodule

