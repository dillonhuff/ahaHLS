module mvmul(input [0:0] clk, input [0:0] rst, output [0:0] valid, output [4:0] ram_debug_addr, input [31:0] ram_debug_data, output [4:0] ram_debug_write_addr, output [31:0] ram_debug_write_data, output [0:0] ram_debug_write_en, output [4:0] ram_raddr_0, output [4:0] ram_raddr_1, output [4:0] ram_raddr_2, input [31:0] ram_rdata_0, input [31:0] ram_rdata_1, input [31:0] ram_rdata_2, output [0:0] ram_rst, output [4:0] ram_waddr_0, output [31:0] ram_wdata_0, output [0:0] ram_wen_0);

	reg [0:0] valid_reg;
	reg [4:0] ram_debug_addr_reg;
	reg [4:0] ram_debug_write_addr_reg;
	reg [31:0] ram_debug_write_data_reg;
	reg [0:0] ram_debug_write_en_reg;
	reg [4:0] ram_raddr_0_reg;
	reg [4:0] ram_raddr_1_reg;
	reg [4:0] ram_raddr_2_reg;
	reg [0:0] ram_rst_reg;
	reg [4:0] ram_waddr_0_reg;
	reg [31:0] ram_wdata_0_reg;
	reg [0:0] ram_wen_0_reg;

	assign valid = valid_reg;
	assign ram_debug_addr = ram_debug_addr_reg;
	assign ram_debug_write_addr = ram_debug_write_addr_reg;
	assign ram_debug_write_data = ram_debug_write_data_reg;
	assign ram_debug_write_en = ram_debug_write_en_reg;
	assign ram_raddr_0 = ram_raddr_0_reg;
	assign ram_raddr_1 = ram_raddr_1_reg;
	assign ram_raddr_2 = ram_raddr_2_reg;
	assign ram_rst = ram_rst_reg;
	assign ram_waddr_0 = ram_waddr_0_reg;
	assign ram_wdata_0 = ram_wdata_0_reg;
	assign ram_wen_0 = ram_wen_0_reg;

	// Start debug wires and ports

	initial begin
	end






	// End debug wires and ports

	// Start Functional Units
	wire [31:0] add_add12_in0;
	wire [31:0] add_add12_in1;
	wire [31:0] add_add12_out;
	add #(.WIDTH(32)) add_add12(.in0(add_add12_in0), .in1(add_add12_in1), .out(add_add12_out));

	wire [31:0] icmp_icmp0_in0;
	wire [31:0] icmp_icmp0_in1;
	wire [0:0] icmp_icmp0_out;
	eq #(.WIDTH(32)) icmp_icmp0(.in0(icmp_icmp0_in0), .in1(icmp_icmp0_in1), .out(icmp_icmp0_out));

	wire [31:0] mul_mul1_in0;
	wire [31:0] mul_mul1_in1;
	wire [31:0] mul_mul1_out;
	mul #(.WIDTH(32)) mul_mul1(.in0(mul_mul1_in0), .in1(mul_mul1_in1), .out(mul_mul1_out));

	wire [31:0] add_add3_in0;
	wire [31:0] add_add3_in1;
	wire [31:0] add_add3_out;
	add #(.WIDTH(32)) add_add3(.in0(add_add3_in0), .in1(add_add3_in1), .out(add_add3_out));

	wire [31:0] mul_mul14_in0;
	wire [31:0] mul_mul14_in1;
	wire [31:0] mul_mul14_out;
	mul #(.WIDTH(32)) mul_mul14(.in0(mul_mul14_in0), .in1(mul_mul14_in1), .out(mul_mul14_out));

	br_dummy br_unit();

	wire [63:0] phi_phi5_in;
	wire [31:0] phi_phi5_last_block;
	wire [63:0] phi_phi5_s;
	wire [31:0] phi_phi5_out;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_phi5(.in(phi_phi5_in), .last_block(phi_phi5_last_block), .out(phi_phi5_out), .s(phi_phi5_s));

	wire [31:0] icmp_icmp16_in0;
	wire [31:0] icmp_icmp16_in1;
	wire [0:0] icmp_icmp16_out;
	eq #(.WIDTH(32)) icmp_icmp16(.in0(icmp_icmp16_in0), .in1(icmp_icmp16_in1), .out(icmp_icmp16_out));

	wire [63:0] phi_phi6_in;
	wire [31:0] phi_phi6_last_block;
	wire [63:0] phi_phi6_s;
	wire [31:0] phi_phi6_out;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_phi6(.in(phi_phi6_in), .last_block(phi_phi6_last_block), .out(phi_phi6_out), .s(phi_phi6_s));

	wire [63:0] phi_phi7_in;
	wire [31:0] phi_phi7_last_block;
	wire [63:0] phi_phi7_s;
	wire [31:0] phi_phi7_out;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_phi7(.in(phi_phi7_in), .last_block(phi_phi7_last_block), .out(phi_phi7_out), .s(phi_phi7_s));

	wire [31:0] add_add8_in0;
	wire [31:0] add_add8_in1;
	wire [31:0] add_add8_out;
	add #(.WIDTH(32)) add_add8(.in0(add_add8_in0), .in1(add_add8_in1), .out(add_add8_out));

	wire [31:0] add_add17_in0;
	wire [31:0] add_add17_in1;
	wire [31:0] add_add17_out;
	add #(.WIDTH(32)) add_add17(.in0(add_add17_in0), .in1(add_add17_in1), .out(add_add17_out));

	wire [31:0] add_add21_in0;
	wire [31:0] add_add21_in1;
	wire [31:0] add_add21_out;
	add #(.WIDTH(32)) add_add21(.in0(add_add21_in0), .in1(add_add21_in1), .out(add_add21_out));

	wire [31:0] add_add10_in0;
	wire [31:0] add_add10_in1;
	wire [31:0] add_add10_out;
	add #(.WIDTH(32)) add_add10(.in0(add_add10_in0), .in1(add_add10_in1), .out(add_add10_out));

	reg [0:0] bb_4_active_in_state_0_in_data;
	wire [0:0] bb_4_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_0(.in_data(bb_4_active_in_state_0_in_data), .out_data(bb_4_active_in_state_0_out_data));

	reg [31:0] bb_4_predecessor_in_state_0_in_data;
	wire [31:0] bb_4_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_0(.in_data(bb_4_predecessor_in_state_0_in_data), .out_data(bb_4_predecessor_in_state_0_out_data));

	reg [0:0] br_4_happened_in_state_0_in_data;
	wire [0:0] br_4_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_0(.in_data(br_4_happened_in_state_0_in_data), .out_data(br_4_happened_in_state_0_out_data));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] bb_1_active_in_state_0_in_data;
	wire [0:0] bb_1_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_0(.in_data(bb_1_active_in_state_0_in_data), .out_data(bb_1_active_in_state_0_out_data));

	reg [31:0] bb_1_predecessor_in_state_0_in_data;
	wire [31:0] bb_1_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_0(.in_data(bb_1_predecessor_in_state_0_in_data), .out_data(bb_1_predecessor_in_state_0_out_data));

	reg [0:0] br_1_happened_in_state_0_in_data;
	wire [0:0] br_1_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened_in_state_0(.in_data(br_1_happened_in_state_0_in_data), .out_data(br_1_happened_in_state_0_out_data));

	reg [0:0] bb_4_active_in_state_1_in_data;
	wire [0:0] bb_4_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_1(.in_data(bb_4_active_in_state_1_in_data), .out_data(bb_4_active_in_state_1_out_data));

	reg [31:0] bb_4_predecessor_in_state_1_in_data;
	wire [31:0] bb_4_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_1(.in_data(bb_4_predecessor_in_state_1_in_data), .out_data(bb_4_predecessor_in_state_1_out_data));

	reg [0:0] br_4_happened_in_state_1_in_data;
	wire [0:0] br_4_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_1(.in_data(br_4_happened_in_state_1_in_data), .out_data(br_4_happened_in_state_1_out_data));

	reg [0:0] bb_3_active_in_state_1_in_data;
	wire [0:0] bb_3_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_1(.in_data(bb_3_active_in_state_1_in_data), .out_data(bb_3_active_in_state_1_out_data));

	reg [31:0] bb_3_predecessor_in_state_1_in_data;
	wire [31:0] bb_3_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_1(.in_data(bb_3_predecessor_in_state_1_in_data), .out_data(bb_3_predecessor_in_state_1_out_data));

	reg [0:0] br_3_happened_in_state_1_in_data;
	wire [0:0] br_3_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_1(.in_data(br_3_happened_in_state_1_in_data), .out_data(br_3_happened_in_state_1_out_data));

	reg [0:0] bb_3_active_in_state_2_in_data;
	wire [0:0] bb_3_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_2(.in_data(bb_3_active_in_state_2_in_data), .out_data(bb_3_active_in_state_2_out_data));

	reg [31:0] bb_3_predecessor_in_state_2_in_data;
	wire [31:0] bb_3_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_2(.in_data(bb_3_predecessor_in_state_2_in_data), .out_data(bb_3_predecessor_in_state_2_out_data));

	reg [0:0] br_3_happened_in_state_2_in_data;
	wire [0:0] br_3_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_2(.in_data(br_3_happened_in_state_2_in_data), .out_data(br_3_happened_in_state_2_out_data));

	reg [0:0] bb_3_active_in_state_3_in_data;
	wire [0:0] bb_3_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_3(.in_data(bb_3_active_in_state_3_in_data), .out_data(bb_3_active_in_state_3_out_data));

	reg [31:0] bb_3_predecessor_in_state_3_in_data;
	wire [31:0] bb_3_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_3(.in_data(bb_3_predecessor_in_state_3_in_data), .out_data(bb_3_predecessor_in_state_3_out_data));

	reg [0:0] br_3_happened_in_state_3_in_data;
	wire [0:0] br_3_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_3(.in_data(br_3_happened_in_state_3_in_data), .out_data(br_3_happened_in_state_3_out_data));

	reg [0:0] bb_2_active_in_state_4_in_data;
	wire [0:0] bb_2_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_4(.in_data(bb_2_active_in_state_4_in_data), .out_data(bb_2_active_in_state_4_out_data));

	reg [31:0] bb_2_predecessor_in_state_4_in_data;
	wire [31:0] bb_2_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_4(.in_data(bb_2_predecessor_in_state_4_in_data), .out_data(bb_2_predecessor_in_state_4_out_data));

	reg [0:0] bb_3_active_in_state_4_in_data;
	wire [0:0] bb_3_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_4(.in_data(bb_3_active_in_state_4_in_data), .out_data(bb_3_active_in_state_4_out_data));

	reg [31:0] bb_3_predecessor_in_state_4_in_data;
	wire [31:0] bb_3_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_4(.in_data(bb_3_predecessor_in_state_4_in_data), .out_data(bb_3_predecessor_in_state_4_out_data));

	reg [0:0] br_3_happened_in_state_4_in_data;
	wire [0:0] br_3_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_4(.in_data(br_3_happened_in_state_4_in_data), .out_data(br_3_happened_in_state_4_out_data));

	reg [31:0] data_in_0_2_in_data;
	wire [31:0] data_in_0_2_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_2(.in_data(data_in_0_2_in_data), .out_data(data_in_0_2_out_data));

	reg [31:0] data_in_0_4_in_data;
	wire [31:0] data_in_0_4_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_4(.in_data(data_in_0_4_in_data), .out_data(data_in_0_4_out_data));

	reg [0:0] data_in_0_6_in_data;
	wire [0:0] data_in_0_6_out_data;
	hls_wire #(.WIDTH(1)) data_in_0_6(.in_data(data_in_0_6_in_data), .out_data(data_in_0_6_out_data));

	reg [31:0] data_in_0_9_in_data;
	wire [31:0] data_in_0_9_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_9(.in_data(data_in_0_9_in_data), .out_data(data_in_0_9_out_data));

	reg [31:0] data_in_0_10_in_data;
	wire [31:0] data_in_0_10_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_10(.in_data(data_in_0_10_in_data), .out_data(data_in_0_10_out_data));

	reg [31:0] data_in_0_12_in_data;
	wire [31:0] data_in_0_12_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_12(.in_data(data_in_0_12_in_data), .out_data(data_in_0_12_out_data));

	reg [0:0] data_in_1_13_in_data;
	wire [0:0] data_in_1_13_out_data;
	hls_wire #(.WIDTH(1)) data_in_1_13(.in_data(data_in_1_13_in_data), .out_data(data_in_1_13_out_data));

	reg [31:0] data_in_1_15_in_data;
	wire [31:0] data_in_1_15_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_15(.in_data(data_in_1_15_in_data), .out_data(data_in_1_15_out_data));

	reg [31:0] data_in_1_17_in_data;
	wire [31:0] data_in_1_17_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_17(.in_data(data_in_1_17_in_data), .out_data(data_in_1_17_out_data));

	reg [0:0] data_in_1_19_in_data;
	wire [0:0] data_in_1_19_out_data;
	hls_wire #(.WIDTH(1)) data_in_1_19(.in_data(data_in_1_19_in_data), .out_data(data_in_1_19_out_data));

	reg [31:0] data_in_1_20_in_data;
	wire [31:0] data_in_1_20_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_20(.in_data(data_in_1_20_in_data), .out_data(data_in_1_20_out_data));

	reg [31:0] data_in_1_22_in_data;
	wire [31:0] data_in_1_22_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_22(.in_data(data_in_1_22_in_data), .out_data(data_in_1_22_out_data));

	reg [31:0] data_in_1_25_in_data;
	wire [31:0] data_in_1_25_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_25(.in_data(data_in_1_25_in_data), .out_data(data_in_1_25_out_data));

	reg [31:0] data_in_2_27_in_data;
	wire [31:0] data_in_2_27_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_27(.in_data(data_in_2_27_in_data), .out_data(data_in_2_27_out_data));

	reg [31:0] data_in_2_29_in_data;
	wire [31:0] data_in_2_29_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_29(.in_data(data_in_2_29_in_data), .out_data(data_in_2_29_out_data));

	reg [0:0] data_in_2_31_in_data;
	wire [0:0] data_in_2_31_out_data;
	hls_wire #(.WIDTH(1)) data_in_2_31(.in_data(data_in_2_31_in_data), .out_data(data_in_2_31_out_data));

	reg [31:0] data_in_2_33_in_data;
	wire [31:0] data_in_2_33_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_33(.in_data(data_in_2_33_in_data), .out_data(data_in_2_33_out_data));

	reg [31:0] data_in_2_35_in_data;
	wire [31:0] data_in_2_35_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_35(.in_data(data_in_2_35_in_data), .out_data(data_in_2_35_out_data));

	reg [31:0] data_in_2_37_in_data;
	wire [31:0] data_in_2_37_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_37(.in_data(data_in_2_37_in_data), .out_data(data_in_2_37_out_data));

	reg [31:0] data_in_3_39_in_data;
	wire [31:0] data_in_3_39_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_39(.in_data(data_in_3_39_in_data), .out_data(data_in_3_39_out_data));

	reg [31:0] data_in_3_41_in_data;
	wire [31:0] data_in_3_41_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_41(.in_data(data_in_3_41_in_data), .out_data(data_in_3_41_out_data));

	reg [0:0] data_in_3_43_in_data;
	wire [0:0] data_in_3_43_out_data;
	hls_wire #(.WIDTH(1)) data_in_3_43(.in_data(data_in_3_43_in_data), .out_data(data_in_3_43_out_data));

	reg [31:0] data_in_3_45_in_data;
	wire [31:0] data_in_3_45_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_45(.in_data(data_in_3_45_in_data), .out_data(data_in_3_45_out_data));

	reg [31:0] data_in_3_47_in_data;
	wire [31:0] data_in_3_47_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_47(.in_data(data_in_3_47_in_data), .out_data(data_in_3_47_out_data));

	reg [31:0] data_in_3_49_in_data;
	wire [31:0] data_in_3_49_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_49(.in_data(data_in_3_49_in_data), .out_data(data_in_3_49_out_data));

	reg [31:0] data_in_4_51_in_data;
	wire [31:0] data_in_4_51_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_51(.in_data(data_in_4_51_in_data), .out_data(data_in_4_51_out_data));

	reg [31:0] data_in_4_53_in_data;
	wire [31:0] data_in_4_53_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_53(.in_data(data_in_4_53_in_data), .out_data(data_in_4_53_out_data));

	reg [0:0] data_in_4_55_in_data;
	wire [0:0] data_in_4_55_out_data;
	hls_wire #(.WIDTH(1)) data_in_4_55(.in_data(data_in_4_55_in_data), .out_data(data_in_4_55_out_data));

	reg [31:0] data_in_4_57_in_data;
	wire [31:0] data_in_4_57_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_57(.in_data(data_in_4_57_in_data), .out_data(data_in_4_57_out_data));

	reg [31:0] data_in_4_59_in_data;
	wire [31:0] data_in_4_59_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_59(.in_data(data_in_4_59_in_data), .out_data(data_in_4_59_out_data));

	reg [31:0] data_in_4_61_in_data;
	wire [31:0] data_in_4_61_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_61(.in_data(data_in_4_61_in_data), .out_data(data_in_4_61_out_data));

	wire [0:0] andOp_62_in0;
	wire [0:0] andOp_62_in1;
	wire [0:0] andOp_62_out;
	andOp #(.WIDTH(1)) andOp_62(.in0(andOp_62_in0), .in1(andOp_62_in1), .out(andOp_62_out));

	wire [0:0] notOp_63_in0;
	wire [0:0] notOp_63_out;
	notOp #(.WIDTH(1)) notOp_63(.in(notOp_63_in0), .out(notOp_63_out));

	wire [0:0] andOp_64_in0;
	wire [0:0] andOp_64_in1;
	wire [0:0] andOp_64_out;
	andOp #(.WIDTH(1)) andOp_64(.in0(andOp_64_in0), .in1(andOp_64_in1), .out(andOp_64_out));

	wire [0:0] notOp_65_in0;
	wire [0:0] notOp_65_out;
	notOp #(.WIDTH(1)) notOp_65(.in(notOp_65_in0), .out(notOp_65_out));

	wire [0:0] andOp_66_in0;
	wire [0:0] andOp_66_in1;
	wire [0:0] andOp_66_out;
	andOp #(.WIDTH(1)) andOp_66(.in0(andOp_66_in0), .in1(andOp_66_in1), .out(andOp_66_out));

	wire [0:0] andOp_67_in0;
	wire [0:0] andOp_67_in1;
	wire [0:0] andOp_67_out;
	andOp #(.WIDTH(1)) andOp_67(.in0(andOp_67_in0), .in1(andOp_67_in1), .out(andOp_67_out));

	wire [0:0] notOp_68_in0;
	wire [0:0] notOp_68_out;
	notOp #(.WIDTH(1)) notOp_68(.in(notOp_68_in0), .out(notOp_68_out));

	wire [0:0] andOp_69_in0;
	wire [0:0] andOp_69_in1;
	wire [0:0] andOp_69_out;
	andOp #(.WIDTH(1)) andOp_69(.in0(andOp_69_in0), .in1(andOp_69_in1), .out(andOp_69_out));

	wire [0:0] notOp_70_in0;
	wire [0:0] notOp_70_out;
	notOp #(.WIDTH(1)) notOp_70(.in(notOp_70_in0), .out(notOp_70_out));

	wire [0:0] andOp_71_in0;
	wire [0:0] andOp_71_in1;
	wire [0:0] andOp_71_out;
	andOp #(.WIDTH(1)) andOp_71(.in0(andOp_71_in0), .in1(andOp_71_in1), .out(andOp_71_out));

	wire [0:0] notOp_72_in0;
	wire [0:0] notOp_72_out;
	notOp #(.WIDTH(1)) notOp_72(.in(notOp_72_in0), .out(notOp_72_out));

	wire [0:0] andOp_73_in0;
	wire [0:0] andOp_73_in1;
	wire [0:0] andOp_73_out;
	andOp #(.WIDTH(1)) andOp_73(.in0(andOp_73_in0), .in1(andOp_73_in1), .out(andOp_73_out));

	wire [0:0] notOp_74_in0;
	wire [0:0] notOp_74_out;
	notOp #(.WIDTH(1)) notOp_74(.in(notOp_74_in0), .out(notOp_74_out));

	wire [0:0] andOp_75_in0;
	wire [0:0] andOp_75_in1;
	wire [0:0] andOp_75_out;
	andOp #(.WIDTH(1)) andOp_75(.in0(andOp_75_in0), .in1(andOp_75_in1), .out(andOp_75_out));

	wire [0:0] andOp_76_in0;
	wire [0:0] andOp_76_in1;
	wire [0:0] andOp_76_out;
	andOp #(.WIDTH(1)) andOp_76(.in0(andOp_76_in0), .in1(andOp_76_in1), .out(andOp_76_out));

	wire [0:0] notOp_77_in0;
	wire [0:0] notOp_77_out;
	notOp #(.WIDTH(1)) notOp_77(.in(notOp_77_in0), .out(notOp_77_out));

	wire [0:0] andOp_78_in0;
	wire [0:0] andOp_78_in1;
	wire [0:0] andOp_78_out;
	andOp #(.WIDTH(1)) andOp_78(.in0(andOp_78_in0), .in1(andOp_78_in1), .out(andOp_78_out));

	wire [0:0] notOp_79_in0;
	wire [0:0] notOp_79_out;
	notOp #(.WIDTH(1)) notOp_79(.in(notOp_79_in0), .out(notOp_79_out));

	wire [0:0] andOp_80_in0;
	wire [0:0] andOp_80_in1;
	wire [0:0] andOp_80_out;
	andOp #(.WIDTH(1)) andOp_80(.in0(andOp_80_in0), .in1(andOp_80_in1), .out(andOp_80_out));

	wire [0:0] andOp_81_in0;
	wire [0:0] andOp_81_in1;
	wire [0:0] andOp_81_out;
	andOp #(.WIDTH(1)) andOp_81(.in0(andOp_81_in0), .in1(andOp_81_in1), .out(andOp_81_out));

	wire [0:0] notOp_82_in0;
	wire [0:0] notOp_82_out;
	notOp #(.WIDTH(1)) notOp_82(.in(notOp_82_in0), .out(notOp_82_out));

	wire [0:0] andOp_83_in0;
	wire [0:0] andOp_83_in1;
	wire [0:0] andOp_83_out;
	andOp #(.WIDTH(1)) andOp_83(.in0(andOp_83_in0), .in1(andOp_83_in1), .out(andOp_83_out));

	wire [0:0] notOp_84_in0;
	wire [0:0] notOp_84_out;
	notOp #(.WIDTH(1)) notOp_84(.in(notOp_84_in0), .out(notOp_84_out));

	wire [0:0] andOp_85_in0;
	wire [0:0] andOp_85_in1;
	wire [0:0] andOp_85_out;
	andOp #(.WIDTH(1)) andOp_85(.in0(andOp_85_in0), .in1(andOp_85_in1), .out(andOp_85_out));

	wire [0:0] andOp_86_in0;
	wire [0:0] andOp_86_in1;
	wire [0:0] andOp_86_out;
	andOp #(.WIDTH(1)) andOp_86(.in0(andOp_86_in0), .in1(andOp_86_in1), .out(andOp_86_out));

	wire [0:0] notOp_87_in0;
	wire [0:0] notOp_87_out;
	notOp #(.WIDTH(1)) notOp_87(.in(notOp_87_in0), .out(notOp_87_out));

	wire [0:0] andOp_88_in0;
	wire [0:0] andOp_88_in1;
	wire [0:0] andOp_88_out;
	andOp #(.WIDTH(1)) andOp_88(.in0(andOp_88_in0), .in1(andOp_88_in1), .out(andOp_88_out));

	wire [0:0] notOp_89_in0;
	wire [0:0] notOp_89_out;
	notOp #(.WIDTH(1)) notOp_89(.in(notOp_89_in0), .out(notOp_89_out));

	wire [0:0] andOp_90_in0;
	wire [0:0] andOp_90_in1;
	wire [0:0] andOp_90_out;
	andOp #(.WIDTH(1)) andOp_90(.in0(andOp_90_in0), .in1(andOp_90_in1), .out(andOp_90_out));

	wire [0:0] andOp_91_in0;
	wire [0:0] andOp_91_in1;
	wire [0:0] andOp_91_out;
	andOp #(.WIDTH(1)) andOp_91(.in0(andOp_91_in0), .in1(andOp_91_in1), .out(andOp_91_out));

	wire [0:0] notOp_92_in0;
	wire [0:0] notOp_92_out;
	notOp #(.WIDTH(1)) notOp_92(.in(notOp_92_in0), .out(notOp_92_out));

	wire [0:0] andOp_93_in0;
	wire [0:0] andOp_93_in1;
	wire [0:0] andOp_93_out;
	andOp #(.WIDTH(1)) andOp_93(.in0(andOp_93_in0), .in1(andOp_93_in1), .out(andOp_93_out));

	wire [0:0] notOp_94_in0;
	wire [0:0] notOp_94_out;
	notOp #(.WIDTH(1)) notOp_94(.in(notOp_94_in0), .out(notOp_94_out));

	wire [0:0] andOp_95_in0;
	wire [0:0] andOp_95_in1;
	wire [0:0] andOp_95_out;
	andOp #(.WIDTH(1)) andOp_95(.in0(andOp_95_in0), .in1(andOp_95_in1), .out(andOp_95_out));

	wire [31:0] eq_96_in0;
	wire [31:0] eq_96_in1;
	wire [0:0] eq_96_out;
	eq #(.WIDTH(32)) eq_96(.in0(eq_96_in0), .in1(eq_96_in1), .out(eq_96_out));

	wire [0:0] orOp_97_in0;
	wire [0:0] orOp_97_in1;
	wire [0:0] orOp_97_out;
	orOp #(.WIDTH(1)) orOp_97(.in0(orOp_97_in0), .in1(orOp_97_in1), .out(orOp_97_out));

	wire [31:0] eq_98_in0;
	wire [31:0] eq_98_in1;
	wire [0:0] eq_98_out;
	eq #(.WIDTH(32)) eq_98(.in0(eq_98_in0), .in1(eq_98_in1), .out(eq_98_out));

	wire [31:0] eq_99_in0;
	wire [31:0] eq_99_in1;
	wire [0:0] eq_99_out;
	eq #(.WIDTH(32)) eq_99(.in0(eq_99_in0), .in1(eq_99_in1), .out(eq_99_out));

	wire [0:0] orOp_100_in0;
	wire [0:0] orOp_100_in1;
	wire [0:0] orOp_100_out;
	orOp #(.WIDTH(1)) orOp_100(.in0(orOp_100_in0), .in1(orOp_100_in1), .out(orOp_100_out));

	wire [31:0] eq_101_in0;
	wire [31:0] eq_101_in1;
	wire [0:0] eq_101_out;
	eq #(.WIDTH(32)) eq_101(.in0(eq_101_in0), .in1(eq_101_in1), .out(eq_101_out));

	wire [31:0] eq_102_in0;
	wire [31:0] eq_102_in1;
	wire [0:0] eq_102_out;
	eq #(.WIDTH(32)) eq_102(.in0(eq_102_in0), .in1(eq_102_in1), .out(eq_102_out));

	wire [0:0] orOp_103_in0;
	wire [0:0] orOp_103_in1;
	wire [0:0] orOp_103_out;
	orOp #(.WIDTH(1)) orOp_103(.in0(orOp_103_in0), .in1(orOp_103_in1), .out(orOp_103_out));

	wire [31:0] eq_104_in0;
	wire [31:0] eq_104_in1;
	wire [0:0] eq_104_out;
	eq #(.WIDTH(32)) eq_104(.in0(eq_104_in0), .in1(eq_104_in1), .out(eq_104_out));

	wire [31:0] eq_105_in0;
	wire [31:0] eq_105_in1;
	wire [0:0] eq_105_out;
	eq #(.WIDTH(32)) eq_105(.in0(eq_105_in0), .in1(eq_105_in1), .out(eq_105_out));

	wire [31:0] eq_106_in0;
	wire [31:0] eq_106_in1;
	wire [0:0] eq_106_out;
	eq #(.WIDTH(32)) eq_106(.in0(eq_106_in0), .in1(eq_106_in1), .out(eq_106_out));

	wire [0:0] orOp_107_in0;
	wire [0:0] orOp_107_in1;
	wire [0:0] orOp_107_out;
	orOp #(.WIDTH(1)) orOp_107(.in0(orOp_107_in0), .in1(orOp_107_in1), .out(orOp_107_out));

	wire [31:0] eq_108_in0;
	wire [31:0] eq_108_in1;
	wire [0:0] eq_108_out;
	eq #(.WIDTH(32)) eq_108(.in0(eq_108_in0), .in1(eq_108_in1), .out(eq_108_out));

	wire [31:0] eq_109_in0;
	wire [31:0] eq_109_in1;
	wire [0:0] eq_109_out;
	eq #(.WIDTH(32)) eq_109(.in0(eq_109_in0), .in1(eq_109_in1), .out(eq_109_out));

	wire [0:0] notOp_110_in0;
	wire [0:0] notOp_110_out;
	notOp #(.WIDTH(1)) notOp_110(.in(notOp_110_in0), .out(notOp_110_out));

	wire [0:0] andOp_111_in0;
	wire [0:0] andOp_111_in1;
	wire [0:0] andOp_111_out;
	andOp #(.WIDTH(1)) andOp_111(.in0(andOp_111_in0), .in1(andOp_111_in1), .out(andOp_111_out));

	wire [31:0] eq_112_in0;
	wire [31:0] eq_112_in1;
	wire [0:0] eq_112_out;
	eq #(.WIDTH(32)) eq_112(.in0(eq_112_in0), .in1(eq_112_in1), .out(eq_112_out));

	wire [31:0] eq_113_in0;
	wire [31:0] eq_113_in1;
	wire [0:0] eq_113_out;
	eq #(.WIDTH(32)) eq_113(.in0(eq_113_in0), .in1(eq_113_in1), .out(eq_113_out));

	wire [0:0] notOp_114_in0;
	wire [0:0] notOp_114_out;
	notOp #(.WIDTH(1)) notOp_114(.in(notOp_114_in0), .out(notOp_114_out));

	wire [0:0] andOp_115_in0;
	wire [0:0] andOp_115_in1;
	wire [0:0] andOp_115_out;
	andOp #(.WIDTH(1)) andOp_115(.in0(andOp_115_in0), .in1(andOp_115_in1), .out(andOp_115_out));

	wire [31:0] eq_116_in0;
	wire [31:0] eq_116_in1;
	wire [0:0] eq_116_out;
	eq #(.WIDTH(32)) eq_116(.in0(eq_116_in0), .in1(eq_116_in1), .out(eq_116_out));

	wire [31:0] eq_117_in0;
	wire [31:0] eq_117_in1;
	wire [0:0] eq_117_out;
	eq #(.WIDTH(32)) eq_117(.in0(eq_117_in0), .in1(eq_117_in1), .out(eq_117_out));

	wire [0:0] notOp_118_in0;
	wire [0:0] notOp_118_out;
	notOp #(.WIDTH(1)) notOp_118(.in(notOp_118_in0), .out(notOp_118_out));

	wire [0:0] andOp_119_in0;
	wire [0:0] andOp_119_in1;
	wire [0:0] andOp_119_out;
	andOp #(.WIDTH(1)) andOp_119(.in0(andOp_119_in0), .in1(andOp_119_in1), .out(andOp_119_out));

	wire [31:0] eq_120_in0;
	wire [31:0] eq_120_in1;
	wire [0:0] eq_120_out;
	eq #(.WIDTH(32)) eq_120(.in0(eq_120_in0), .in1(eq_120_in1), .out(eq_120_out));

	wire [31:0] eq_121_in0;
	wire [31:0] eq_121_in1;
	wire [0:0] eq_121_out;
	eq #(.WIDTH(32)) eq_121(.in0(eq_121_in0), .in1(eq_121_in1), .out(eq_121_out));

	wire [31:0] eq_122_in0;
	wire [31:0] eq_122_in1;
	wire [0:0] eq_122_out;
	eq #(.WIDTH(32)) eq_122(.in0(eq_122_in0), .in1(eq_122_in1), .out(eq_122_out));

	wire [0:0] notOp_123_in0;
	wire [0:0] notOp_123_out;
	notOp #(.WIDTH(1)) notOp_123(.in(notOp_123_in0), .out(notOp_123_out));

	wire [0:0] andOp_124_in0;
	wire [0:0] andOp_124_in1;
	wire [0:0] andOp_124_out;
	andOp #(.WIDTH(1)) andOp_124(.in0(andOp_124_in0), .in1(andOp_124_in1), .out(andOp_124_out));

	wire [31:0] eq_125_in0;
	wire [31:0] eq_125_in1;
	wire [0:0] eq_125_out;
	eq #(.WIDTH(32)) eq_125(.in0(eq_125_in0), .in1(eq_125_in1), .out(eq_125_out));

	wire [0:0] andOp_126_in0;
	wire [0:0] andOp_126_in1;
	wire [0:0] andOp_126_out;
	andOp #(.WIDTH(1)) andOp_126(.in0(andOp_126_in0), .in1(andOp_126_in1), .out(andOp_126_out));

	wire [0:0] andOp_127_in0;
	wire [0:0] andOp_127_in1;
	wire [0:0] andOp_127_out;
	andOp #(.WIDTH(1)) andOp_127(.in0(andOp_127_in0), .in1(andOp_127_in1), .out(andOp_127_out));

	wire [0:0] andOp_128_in0;
	wire [0:0] andOp_128_in1;
	wire [0:0] andOp_128_out;
	andOp #(.WIDTH(1)) andOp_128(.in0(andOp_128_in0), .in1(andOp_128_in1), .out(andOp_128_out));

	wire [0:0] andOp_129_in0;
	wire [0:0] andOp_129_in1;
	wire [0:0] andOp_129_out;
	andOp #(.WIDTH(1)) andOp_129(.in0(andOp_129_in0), .in1(andOp_129_in1), .out(andOp_129_out));

	wire [0:0] andOp_130_in0;
	wire [0:0] andOp_130_in1;
	wire [0:0] andOp_130_out;
	andOp #(.WIDTH(1)) andOp_130(.in0(andOp_130_in0), .in1(andOp_130_in1), .out(andOp_130_out));

	wire [0:0] andOp_131_in0;
	wire [0:0] andOp_131_in1;
	wire [0:0] andOp_131_out;
	andOp #(.WIDTH(1)) andOp_131(.in0(andOp_131_in0), .in1(andOp_131_in1), .out(andOp_131_out));

	wire [0:0] andOp_132_in0;
	wire [0:0] andOp_132_in1;
	wire [0:0] andOp_132_out;
	andOp #(.WIDTH(1)) andOp_132(.in0(andOp_132_in0), .in1(andOp_132_in1), .out(andOp_132_out));

	reg [31:0] tmp_output_133_in_data;
	wire [31:0] tmp_output_133_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_133(.in_data(tmp_output_133_in_data), .out_data(tmp_output_133_out_data));

	wire [31:0] eq_134_in0;
	wire [31:0] eq_134_in1;
	wire [0:0] eq_134_out;
	eq #(.WIDTH(32)) eq_134(.in0(eq_134_in0), .in1(eq_134_in1), .out(eq_134_out));

	wire [0:0] andOp_135_in0;
	wire [0:0] andOp_135_in1;
	wire [0:0] andOp_135_out;
	andOp #(.WIDTH(1)) andOp_135(.in0(andOp_135_in0), .in1(andOp_135_in1), .out(andOp_135_out));

	wire [0:0] andOp_136_in0;
	wire [0:0] andOp_136_in1;
	wire [0:0] andOp_136_out;
	andOp #(.WIDTH(1)) andOp_136(.in0(andOp_136_in0), .in1(andOp_136_in1), .out(andOp_136_out));

	wire [0:0] andOp_137_in0;
	wire [0:0] andOp_137_in1;
	wire [0:0] andOp_137_out;
	andOp #(.WIDTH(1)) andOp_137(.in0(andOp_137_in0), .in1(andOp_137_in1), .out(andOp_137_out));

	wire [0:0] andOp_138_in0;
	wire [0:0] andOp_138_in1;
	wire [0:0] andOp_138_out;
	andOp #(.WIDTH(1)) andOp_138(.in0(andOp_138_in0), .in1(andOp_138_in1), .out(andOp_138_out));

	wire [31:0] concat_139_in0;
	wire [31:0] concat_139_in1;
	wire [63:0] concat_139_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_139(.in0(concat_139_in0), .in1(concat_139_in1), .out(concat_139_out));

	wire [31:0] concat_140_in0;
	wire [31:0] concat_140_in1;
	wire [63:0] concat_140_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_140(.in0(concat_140_in0), .in1(concat_140_in1), .out(concat_140_out));

	wire [0:0] andOp_141_in0;
	wire [0:0] andOp_141_in1;
	wire [0:0] andOp_141_out;
	andOp #(.WIDTH(1)) andOp_141(.in0(andOp_141_in0), .in1(andOp_141_in1), .out(andOp_141_out));

	wire [31:0] concat_142_in0;
	wire [31:0] concat_142_in1;
	wire [63:0] concat_142_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_142(.in0(concat_142_in0), .in1(concat_142_in1), .out(concat_142_out));

	wire [31:0] concat_143_in0;
	wire [31:0] concat_143_in1;
	wire [63:0] concat_143_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_143(.in0(concat_143_in0), .in1(concat_143_in1), .out(concat_143_out));

	wire [0:0] andOp_144_in0;
	wire [0:0] andOp_144_in1;
	wire [0:0] andOp_144_out;
	andOp #(.WIDTH(1)) andOp_144(.in0(andOp_144_in0), .in1(andOp_144_in1), .out(andOp_144_out));

	wire [31:0] concat_145_in0;
	wire [31:0] concat_145_in1;
	wire [63:0] concat_145_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_145(.in0(concat_145_in0), .in1(concat_145_in1), .out(concat_145_out));

	wire [31:0] concat_146_in0;
	wire [31:0] concat_146_in1;
	wire [63:0] concat_146_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_146(.in0(concat_146_in0), .in1(concat_146_in1), .out(concat_146_out));

	wire [0:0] andOp_147_in0;
	wire [0:0] andOp_147_in1;
	wire [0:0] andOp_147_out;
	andOp #(.WIDTH(1)) andOp_147(.in0(andOp_147_in0), .in1(andOp_147_in1), .out(andOp_147_out));

	reg [31:0] tmp_output_148_in_data;
	wire [31:0] tmp_output_148_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_148(.in_data(tmp_output_148_in_data), .out_data(tmp_output_148_out_data));

	wire [31:0] eq_149_in0;
	wire [31:0] eq_149_in1;
	wire [0:0] eq_149_out;
	eq #(.WIDTH(32)) eq_149(.in0(eq_149_in0), .in1(eq_149_in1), .out(eq_149_out));

	wire [31:0] eq_150_in0;
	wire [31:0] eq_150_in1;
	wire [0:0] eq_150_out;
	eq #(.WIDTH(32)) eq_150(.in0(eq_150_in0), .in1(eq_150_in1), .out(eq_150_out));

	wire [31:0] eq_151_in0;
	wire [31:0] eq_151_in1;
	wire [0:0] eq_151_out;
	eq #(.WIDTH(32)) eq_151(.in0(eq_151_in0), .in1(eq_151_in1), .out(eq_151_out));

	wire [0:0] andOp_152_in0;
	wire [0:0] andOp_152_in1;
	wire [0:0] andOp_152_out;
	andOp #(.WIDTH(1)) andOp_152(.in0(andOp_152_in0), .in1(andOp_152_in1), .out(andOp_152_out));

	wire [0:0] andOp_153_in0;
	wire [0:0] andOp_153_in1;
	wire [0:0] andOp_153_out;
	andOp #(.WIDTH(1)) andOp_153(.in0(andOp_153_in0), .in1(andOp_153_in1), .out(andOp_153_out));

	wire [0:0] andOp_154_in0;
	wire [0:0] andOp_154_in1;
	wire [0:0] andOp_154_out;
	andOp #(.WIDTH(1)) andOp_154(.in0(andOp_154_in0), .in1(andOp_154_in1), .out(andOp_154_out));

	wire [0:0] andOp_155_in0;
	wire [0:0] andOp_155_in1;
	wire [0:0] andOp_155_out;
	andOp #(.WIDTH(1)) andOp_155(.in0(andOp_155_in0), .in1(andOp_155_in1), .out(andOp_155_out));

	wire [0:0] andOp_156_in0;
	wire [0:0] andOp_156_in1;
	wire [0:0] andOp_156_out;
	andOp #(.WIDTH(1)) andOp_156(.in0(andOp_156_in0), .in1(andOp_156_in1), .out(andOp_156_out));

	wire [0:0] andOp_157_in0;
	wire [0:0] andOp_157_in1;
	wire [0:0] andOp_157_out;
	andOp #(.WIDTH(1)) andOp_157(.in0(andOp_157_in0), .in1(andOp_157_in1), .out(andOp_157_out));

	wire [0:0] andOp_158_in0;
	wire [0:0] andOp_158_in1;
	wire [0:0] andOp_158_out;
	andOp #(.WIDTH(1)) andOp_158(.in0(andOp_158_in0), .in1(andOp_158_in1), .out(andOp_158_out));

	wire [0:0] andOp_159_in0;
	wire [0:0] andOp_159_in1;
	wire [0:0] andOp_159_out;
	andOp #(.WIDTH(1)) andOp_159(.in0(andOp_159_in0), .in1(andOp_159_in1), .out(andOp_159_out));

	wire [0:0] andOp_160_in0;
	wire [0:0] andOp_160_in1;
	wire [0:0] andOp_160_out;
	andOp #(.WIDTH(1)) andOp_160(.in0(andOp_160_in0), .in1(andOp_160_in1), .out(andOp_160_out));

	wire [0:0] andOp_161_in0;
	wire [0:0] andOp_161_in1;
	wire [0:0] andOp_161_out;
	andOp #(.WIDTH(1)) andOp_161(.in0(andOp_161_in0), .in1(andOp_161_in1), .out(andOp_161_out));

	wire [0:0] andOp_162_in0;
	wire [0:0] andOp_162_in1;
	wire [0:0] andOp_162_out;
	andOp #(.WIDTH(1)) andOp_162(.in0(andOp_162_in0), .in1(andOp_162_in1), .out(andOp_162_out));

	wire [0:0] andOp_163_in0;
	wire [0:0] andOp_163_in1;
	wire [0:0] andOp_163_out;
	andOp #(.WIDTH(1)) andOp_163(.in0(andOp_163_in0), .in1(andOp_163_in1), .out(andOp_163_out));

	wire [0:0] notOp_164_in0;
	wire [0:0] notOp_164_out;
	notOp #(.WIDTH(1)) notOp_164(.in(notOp_164_in0), .out(notOp_164_out));

	wire [0:0] andOp_165_in0;
	wire [0:0] andOp_165_in1;
	wire [0:0] andOp_165_out;
	andOp #(.WIDTH(1)) andOp_165(.in0(andOp_165_in0), .in1(andOp_165_in1), .out(andOp_165_out));

	wire [0:0] notOp_166_in0;
	wire [0:0] notOp_166_out;
	notOp #(.WIDTH(1)) notOp_166(.in(notOp_166_in0), .out(notOp_166_out));

	wire [0:0] andOp_167_in0;
	wire [0:0] andOp_167_in1;
	wire [0:0] andOp_167_out;
	andOp #(.WIDTH(1)) andOp_167(.in0(andOp_167_in0), .in1(andOp_167_in1), .out(andOp_167_out));

	wire [0:0] notOp_168_in0;
	wire [0:0] notOp_168_out;
	notOp #(.WIDTH(1)) notOp_168(.in(notOp_168_in0), .out(notOp_168_out));

	wire [0:0] andOp_169_in0;
	wire [0:0] andOp_169_in1;
	wire [0:0] andOp_169_out;
	andOp #(.WIDTH(1)) andOp_169(.in0(andOp_169_in0), .in1(andOp_169_in1), .out(andOp_169_out));

	wire [0:0] notOp_170_in0;
	wire [0:0] notOp_170_out;
	notOp #(.WIDTH(1)) notOp_170(.in(notOp_170_in0), .out(notOp_170_out));

	wire [0:0] andOp_171_in0;
	wire [0:0] andOp_171_in1;
	wire [0:0] andOp_171_out;
	andOp #(.WIDTH(1)) andOp_171(.in0(andOp_171_in0), .in1(andOp_171_in1), .out(andOp_171_out));

	wire [0:0] notOp_172_in0;
	wire [0:0] notOp_172_out;
	notOp #(.WIDTH(1)) notOp_172(.in(notOp_172_in0), .out(notOp_172_out));

	wire [0:0] andOp_173_in0;
	wire [0:0] andOp_173_in1;
	wire [0:0] andOp_173_out;
	andOp #(.WIDTH(1)) andOp_173(.in0(andOp_173_in0), .in1(andOp_173_in1), .out(andOp_173_out));

	wire [0:0] notOp_174_in0;
	wire [0:0] notOp_174_out;
	notOp #(.WIDTH(1)) notOp_174(.in(notOp_174_in0), .out(notOp_174_out));

	wire [0:0] andOp_175_in0;
	wire [0:0] andOp_175_in1;
	wire [0:0] andOp_175_out;
	andOp #(.WIDTH(1)) andOp_175(.in0(andOp_175_in0), .in1(andOp_175_in1), .out(andOp_175_out));

	wire [0:0] notOp_176_in0;
	wire [0:0] notOp_176_out;
	notOp #(.WIDTH(1)) notOp_176(.in(notOp_176_in0), .out(notOp_176_out));

	wire [0:0] andOp_177_in0;
	wire [0:0] andOp_177_in1;
	wire [0:0] andOp_177_out;
	andOp #(.WIDTH(1)) andOp_177(.in0(andOp_177_in0), .in1(andOp_177_in1), .out(andOp_177_out));

	wire [31:0] eq_178_in0;
	wire [31:0] eq_178_in1;
	wire [0:0] eq_178_out;
	eq #(.WIDTH(32)) eq_178(.in0(eq_178_in0), .in1(eq_178_in1), .out(eq_178_out));

	wire [31:0] eq_179_in0;
	wire [31:0] eq_179_in1;
	wire [0:0] eq_179_out;
	eq #(.WIDTH(32)) eq_179(.in0(eq_179_in0), .in1(eq_179_in1), .out(eq_179_out));

	wire [31:0] eq_180_in0;
	wire [31:0] eq_180_in1;
	wire [0:0] eq_180_out;
	eq #(.WIDTH(32)) eq_180(.in0(eq_180_in0), .in1(eq_180_in1), .out(eq_180_out));

	wire [0:0] andOp_181_in0;
	wire [0:0] andOp_181_in1;
	wire [0:0] andOp_181_out;
	andOp #(.WIDTH(1)) andOp_181(.in0(andOp_181_in0), .in1(andOp_181_in1), .out(andOp_181_out));

	wire [0:0] andOp_182_in0;
	wire [0:0] andOp_182_in1;
	wire [0:0] andOp_182_out;
	andOp #(.WIDTH(1)) andOp_182(.in0(andOp_182_in0), .in1(andOp_182_in1), .out(andOp_182_out));

	wire [0:0] andOp_183_in0;
	wire [0:0] andOp_183_in1;
	wire [0:0] andOp_183_out;
	andOp #(.WIDTH(1)) andOp_183(.in0(andOp_183_in0), .in1(andOp_183_in1), .out(andOp_183_out));

	wire [0:0] andOp_184_in0;
	wire [0:0] andOp_184_in1;
	wire [0:0] andOp_184_out;
	andOp #(.WIDTH(1)) andOp_184(.in0(andOp_184_in0), .in1(andOp_184_in1), .out(andOp_184_out));

	wire [0:0] andOp_185_in0;
	wire [0:0] andOp_185_in1;
	wire [0:0] andOp_185_out;
	andOp #(.WIDTH(1)) andOp_185(.in0(andOp_185_in0), .in1(andOp_185_in1), .out(andOp_185_out));

	wire [31:0] eq_186_in0;
	wire [31:0] eq_186_in1;
	wire [0:0] eq_186_out;
	eq #(.WIDTH(32)) eq_186(.in0(eq_186_in0), .in1(eq_186_in1), .out(eq_186_out));

	wire [31:0] eq_187_in0;
	wire [31:0] eq_187_in1;
	wire [0:0] eq_187_out;
	eq #(.WIDTH(32)) eq_187(.in0(eq_187_in0), .in1(eq_187_in1), .out(eq_187_out));

	wire [0:0] andOp_188_in0;
	wire [0:0] andOp_188_in1;
	wire [0:0] andOp_188_out;
	andOp #(.WIDTH(1)) andOp_188(.in0(andOp_188_in0), .in1(andOp_188_in1), .out(andOp_188_out));

	wire [0:0] andOp_189_in0;
	wire [0:0] andOp_189_in1;
	wire [0:0] andOp_189_out;
	andOp #(.WIDTH(1)) andOp_189(.in0(andOp_189_in0), .in1(andOp_189_in1), .out(andOp_189_out));

	wire [0:0] andOp_190_in0;
	wire [0:0] andOp_190_in1;
	wire [0:0] andOp_190_out;
	andOp #(.WIDTH(1)) andOp_190(.in0(andOp_190_in0), .in1(andOp_190_in1), .out(andOp_190_out));

	wire [31:0] eq_191_in0;
	wire [31:0] eq_191_in1;
	wire [0:0] eq_191_out;
	eq #(.WIDTH(32)) eq_191(.in0(eq_191_in0), .in1(eq_191_in1), .out(eq_191_out));

	wire [31:0] eq_192_in0;
	wire [31:0] eq_192_in1;
	wire [0:0] eq_192_out;
	eq #(.WIDTH(32)) eq_192(.in0(eq_192_in0), .in1(eq_192_in1), .out(eq_192_out));

	wire [31:0] eq_193_in0;
	wire [31:0] eq_193_in1;
	wire [0:0] eq_193_out;
	eq #(.WIDTH(32)) eq_193(.in0(eq_193_in0), .in1(eq_193_in1), .out(eq_193_out));

	wire [31:0] eq_194_in0;
	wire [31:0] eq_194_in1;
	wire [0:0] eq_194_out;
	eq #(.WIDTH(32)) eq_194(.in0(eq_194_in0), .in1(eq_194_in1), .out(eq_194_out));

	wire [31:0] eq_195_in0;
	wire [31:0] eq_195_in1;
	wire [0:0] eq_195_out;
	eq #(.WIDTH(32)) eq_195(.in0(eq_195_in0), .in1(eq_195_in1), .out(eq_195_out));

	wire [31:0] eq_196_in0;
	wire [31:0] eq_196_in1;
	wire [0:0] eq_196_out;
	eq #(.WIDTH(32)) eq_196(.in0(eq_196_in0), .in1(eq_196_in1), .out(eq_196_out));

	// End Functional Units

	reg [0:0] data_store_0_0;
	reg [31:0] data_store_0_1;
	reg [31:0] data_store_0_11;
	reg [31:0] data_store_0_3;
	reg [0:0] data_store_0_5;
	reg [31:0] data_store_0_7;
	reg [31:0] data_store_0_8;
	reg [31:0] data_store_1_14;
	reg [31:0] data_store_1_16;
	reg [0:0] data_store_1_18;
	reg [31:0] data_store_1_21;
	reg [31:0] data_store_1_23;
	reg [31:0] data_store_1_24;
	reg [31:0] data_store_2_26;
	reg [31:0] data_store_2_28;
	reg [0:0] data_store_2_30;
	reg [31:0] data_store_2_32;
	reg [31:0] data_store_2_34;
	reg [31:0] data_store_2_36;
	reg [31:0] data_store_3_38;
	reg [31:0] data_store_3_40;
	reg [0:0] data_store_3_42;
	reg [31:0] data_store_3_44;
	reg [31:0] data_store_3_46;
	reg [31:0] data_store_3_48;
	reg [31:0] data_store_4_50;
	reg [31:0] data_store_4_52;
	reg [0:0] data_store_4_54;
	reg [31:0] data_store_4_56;
	reg [31:0] data_store_4_58;
	reg [31:0] data_store_4_60;
	reg [31:0] global_state;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_3_last_state;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;
	reg [31:0] state_4_last_state;

	// controller for add_add10.add_add10_in0
	// controller for add_add10.add_add10_in1
	// Insensitive connections
	assign add_add10_in0 = phi_phi6_out;
	assign add_add10_in1 = 32'd1;
	// controller for add_add12.add_add12_in0
	// controller for add_add12.add_add12_in1
	// Insensitive connections
	assign add_add12_in0 = data_in_1_17_out_data;
	assign add_add12_in1 = 32'd12;
	// controller for add_add17.add_add17_in0
	// controller for add_add17.add_add17_in1
	// Insensitive connections
	assign add_add17_in0 = data_in_1_17_out_data;
	assign add_add17_in1 = 32'd1;
	// controller for add_add21.add_add21_in0
	// controller for add_add21.add_add21_in1
	// Insensitive connections
	assign add_add21_in0 = mul_mul14_out;
	assign add_add21_in1 = data_in_1_20_out_data;
	// controller for add_add3.add_add3_in0
	// controller for add_add3.add_add3_in1
	// Insensitive connections
	assign add_add3_in0 = phi_phi6_out;
	assign add_add3_in1 = 32'd9;
	// controller for add_add8.add_add8_in0
	// controller for add_add8.add_add8_in1
	// Insensitive connections
	assign add_add8_in0 = phi_phi6_out;
	assign add_add8_in1 = tmp_output_148_out_data;
	// controller for andOp_111.andOp_111_in0
	// controller for andOp_111.andOp_111_in1
	// Insensitive connections
	assign andOp_111_in0 = notOp_110_out;
	assign andOp_111_in1 = andOp_69_out;
	// controller for andOp_115.andOp_115_in0
	// controller for andOp_115.andOp_115_in1
	// Insensitive connections
	assign andOp_115_in0 = notOp_114_out;
	assign andOp_115_in1 = andOp_67_out;
	// controller for andOp_119.andOp_119_in0
	// controller for andOp_119.andOp_119_in1
	// Insensitive connections
	assign andOp_119_in0 = notOp_118_out;
	assign andOp_119_in1 = andOp_64_out;
	// controller for andOp_124.andOp_124_in0
	// controller for andOp_124.andOp_124_in1
	// Insensitive connections
	assign andOp_124_in0 = notOp_123_out;
	assign andOp_124_in1 = andOp_78_out;
	// controller for andOp_126.andOp_126_in0
	// controller for andOp_126.andOp_126_in1
	// Insensitive connections
	assign andOp_126_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_126_in1 = state_0_is_active;
	// controller for andOp_127.andOp_127_in0
	// controller for andOp_127.andOp_127_in1
	// Insensitive connections
	assign andOp_127_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_127_in1 = state_0_is_active;
	// controller for andOp_128.andOp_128_in0
	// controller for andOp_128.andOp_128_in1
	// Insensitive connections
	assign andOp_128_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_128_in1 = state_0_is_active;
	// controller for andOp_129.andOp_129_in0
	// controller for andOp_129.andOp_129_in1
	// Insensitive connections
	assign andOp_129_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_129_in1 = state_0_is_active;
	// controller for andOp_130.andOp_130_in0
	// controller for andOp_130.andOp_130_in1
	// Insensitive connections
	assign andOp_130_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_130_in1 = state_1_is_active;
	// controller for andOp_131.andOp_131_in0
	// controller for andOp_131.andOp_131_in1
	// Insensitive connections
	assign andOp_131_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_131_in1 = state_1_is_active;
	// controller for andOp_132.andOp_132_in0
	// controller for andOp_132.andOp_132_in1
	// Insensitive connections
	assign andOp_132_in0 = bb_3_active_in_state_1_out_data;
	assign andOp_132_in1 = state_1_is_active;
	// controller for andOp_135.andOp_135_in0
	// controller for andOp_135.andOp_135_in1
	// Insensitive connections
	assign andOp_135_in0 = bb_3_active_in_state_1_out_data;
	assign andOp_135_in1 = state_1_is_active;
	// controller for andOp_136.andOp_136_in0
	// controller for andOp_136.andOp_136_in1
	// Insensitive connections
	assign andOp_136_in0 = bb_3_active_in_state_1_out_data;
	assign andOp_136_in1 = state_1_is_active;
	// controller for andOp_137.andOp_137_in0
	// controller for andOp_137.andOp_137_in1
	// Insensitive connections
	assign andOp_137_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_137_in1 = state_0_is_active;
	// controller for andOp_138.andOp_138_in0
	// controller for andOp_138.andOp_138_in1
	// Insensitive connections
	assign andOp_138_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_138_in1 = state_0_is_active;
	// controller for andOp_141.andOp_141_in0
	// controller for andOp_141.andOp_141_in1
	// Insensitive connections
	assign andOp_141_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_141_in1 = state_0_is_active;
	// controller for andOp_144.andOp_144_in0
	// controller for andOp_144.andOp_144_in1
	// Insensitive connections
	assign andOp_144_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_144_in1 = state_0_is_active;
	// controller for andOp_147.andOp_147_in0
	// controller for andOp_147.andOp_147_in1
	// Insensitive connections
	assign andOp_147_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_147_in1 = state_0_is_active;
	// controller for andOp_152.andOp_152_in0
	// controller for andOp_152.andOp_152_in1
	// Insensitive connections
	assign andOp_152_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_152_in1 = state_0_is_active;
	// controller for andOp_153.andOp_153_in0
	// controller for andOp_153.andOp_153_in1
	// Insensitive connections
	assign andOp_153_in0 = bb_3_active_in_state_1_out_data;
	assign andOp_153_in1 = state_1_is_active;
	// controller for andOp_154.andOp_154_in0
	// controller for andOp_154.andOp_154_in1
	// Insensitive connections
	assign andOp_154_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_154_in1 = state_1_is_active;
	// controller for andOp_155.andOp_155_in0
	// controller for andOp_155.andOp_155_in1
	// Insensitive connections
	assign andOp_155_in0 = bb_3_active_in_state_1_out_data;
	assign andOp_155_in1 = state_1_is_active;
	// controller for andOp_156.andOp_156_in0
	// controller for andOp_156.andOp_156_in1
	// Insensitive connections
	assign andOp_156_in0 = bb_3_active_in_state_1_out_data;
	assign andOp_156_in1 = state_1_is_active;
	// controller for andOp_157.andOp_157_in0
	// controller for andOp_157.andOp_157_in1
	// Insensitive connections
	assign andOp_157_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_157_in1 = state_1_is_active;
	// controller for andOp_158.andOp_158_in0
	// controller for andOp_158.andOp_158_in1
	// Insensitive connections
	assign andOp_158_in0 = bb_2_active_in_state_4_out_data;
	assign andOp_158_in1 = state_4_is_active;
	// controller for andOp_159.andOp_159_in0
	// controller for andOp_159.andOp_159_in1
	// Insensitive connections
	assign andOp_159_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_159_in1 = state_0_is_active;
	// controller for andOp_160.andOp_160_in0
	// controller for andOp_160.andOp_160_in1
	// Insensitive connections
	assign andOp_160_in0 = bb_3_active_in_state_1_out_data;
	assign andOp_160_in1 = state_1_is_active;
	// controller for andOp_161.andOp_161_in0
	// controller for andOp_161.andOp_161_in1
	// Insensitive connections
	assign andOp_161_in0 = bb_3_active_in_state_2_out_data;
	assign andOp_161_in1 = state_2_is_active;
	// controller for andOp_162.andOp_162_in0
	// controller for andOp_162.andOp_162_in1
	// Insensitive connections
	assign andOp_162_in0 = bb_3_active_in_state_3_out_data;
	assign andOp_162_in1 = state_3_is_active;
	// controller for andOp_163.andOp_163_in0
	// controller for andOp_163.andOp_163_in1
	// Insensitive connections
	assign andOp_163_in0 = bb_2_active_in_state_4_out_data;
	assign andOp_163_in1 = state_4_is_active;
	// controller for andOp_165.andOp_165_in0
	// controller for andOp_165.andOp_165_in1
	// Insensitive connections
	assign andOp_165_in0 = notOp_164_out;
	assign andOp_165_in1 = 1'd1;
	// controller for andOp_167.andOp_167_in0
	// controller for andOp_167.andOp_167_in1
	// Insensitive connections
	assign andOp_167_in0 = notOp_166_out;
	assign andOp_167_in1 = andOp_165_out;
	// controller for andOp_169.andOp_169_in0
	// controller for andOp_169.andOp_169_in1
	// Insensitive connections
	assign andOp_169_in0 = notOp_168_out;
	assign andOp_169_in1 = 1'd1;
	// controller for andOp_171.andOp_171_in0
	// controller for andOp_171.andOp_171_in1
	// Insensitive connections
	assign andOp_171_in0 = notOp_170_out;
	assign andOp_171_in1 = 1'd1;
	// controller for andOp_173.andOp_173_in0
	// controller for andOp_173.andOp_173_in1
	// Insensitive connections
	assign andOp_173_in0 = notOp_172_out;
	assign andOp_173_in1 = 1'd1;
	// controller for andOp_175.andOp_175_in0
	// controller for andOp_175.andOp_175_in1
	// Insensitive connections
	assign andOp_175_in0 = notOp_174_out;
	assign andOp_175_in1 = 1'd1;
	// controller for andOp_177.andOp_177_in0
	// controller for andOp_177.andOp_177_in1
	// Insensitive connections
	assign andOp_177_in0 = notOp_176_out;
	assign andOp_177_in1 = andOp_175_out;
	// controller for andOp_181.andOp_181_in0
	// controller for andOp_181.andOp_181_in1
	// Insensitive connections
	assign andOp_181_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_181_in1 = state_0_is_active;
	// controller for andOp_182.andOp_182_in0
	// controller for andOp_182.andOp_182_in1
	// Insensitive connections
	assign andOp_182_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_182_in1 = state_0_is_active;
	// controller for andOp_183.andOp_183_in0
	// controller for andOp_183.andOp_183_in1
	// Insensitive connections
	assign andOp_183_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_183_in1 = state_0_is_active;
	// controller for andOp_184.andOp_184_in0
	// controller for andOp_184.andOp_184_in1
	// Insensitive connections
	assign andOp_184_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_184_in1 = state_0_is_active;
	// controller for andOp_185.andOp_185_in0
	// controller for andOp_185.andOp_185_in1
	// Insensitive connections
	assign andOp_185_in0 = bb_4_active_in_state_0_out_data;
	assign andOp_185_in1 = state_0_is_active;
	// controller for andOp_188.andOp_188_in0
	// controller for andOp_188.andOp_188_in1
	// Insensitive connections
	assign andOp_188_in0 = bb_3_active_in_state_1_out_data;
	assign andOp_188_in1 = state_1_is_active;
	// controller for andOp_189.andOp_189_in0
	// controller for andOp_189.andOp_189_in1
	// Insensitive connections
	assign andOp_189_in0 = bb_3_active_in_state_1_out_data;
	assign andOp_189_in1 = state_1_is_active;
	// controller for andOp_190.andOp_190_in0
	// controller for andOp_190.andOp_190_in1
	// Insensitive connections
	assign andOp_190_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_190_in1 = state_1_is_active;
	// controller for andOp_62.andOp_62_in0
	// controller for andOp_62.andOp_62_in1
	// Insensitive connections
	assign andOp_62_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_62_in1 = state_1_is_active;
	// controller for andOp_64.andOp_64_in0
	// controller for andOp_64.andOp_64_in1
	// Insensitive connections
	assign andOp_64_in0 = andOp_62_out;
	assign andOp_64_in1 = data_in_1_13_out_data;
	// controller for andOp_66.andOp_66_in0
	// controller for andOp_66.andOp_66_in1
	// Insensitive connections
	assign andOp_66_in0 = andOp_62_out;
	assign andOp_66_in1 = notOp_65_out;
	// controller for andOp_67.andOp_67_in0
	// controller for andOp_67.andOp_67_in1
	// Insensitive connections
	assign andOp_67_in0 = bb_0_active_in_state_0_out_data;
	assign andOp_67_in1 = state_0_is_active;
	// controller for andOp_69.andOp_69_in0
	// controller for andOp_69.andOp_69_in1
	// Insensitive connections
	assign andOp_69_in0 = bb_1_active_in_state_0_out_data;
	assign andOp_69_in1 = state_0_is_active;
	// controller for andOp_71.andOp_71_in0
	// controller for andOp_71.andOp_71_in1
	// Insensitive connections
	assign andOp_71_in0 = bb_4_active_in_state_1_out_data;
	assign andOp_71_in1 = state_1_is_active;
	// controller for andOp_73.andOp_73_in0
	// controller for andOp_73.andOp_73_in1
	// Insensitive connections
	assign andOp_73_in0 = andOp_71_out;
	assign andOp_73_in1 = data_in_1_13_out_data;
	// controller for andOp_75.andOp_75_in0
	// controller for andOp_75.andOp_75_in1
	// Insensitive connections
	assign andOp_75_in0 = andOp_71_out;
	assign andOp_75_in1 = notOp_74_out;
	// controller for andOp_76.andOp_76_in0
	// controller for andOp_76.andOp_76_in1
	// Insensitive connections
	assign andOp_76_in0 = bb_3_active_in_state_4_out_data;
	assign andOp_76_in1 = state_4_is_active;
	// controller for andOp_78.andOp_78_in0
	// controller for andOp_78.andOp_78_in1
	// Insensitive connections
	assign andOp_78_in0 = andOp_76_out;
	assign andOp_78_in1 = data_in_4_55_out_data;
	// controller for andOp_80.andOp_80_in0
	// controller for andOp_80.andOp_80_in1
	// Insensitive connections
	assign andOp_80_in0 = andOp_76_out;
	assign andOp_80_in1 = notOp_79_out;
	// controller for andOp_81.andOp_81_in0
	// controller for andOp_81.andOp_81_in1
	// Insensitive connections
	assign andOp_81_in0 = bb_3_active_in_state_4_out_data;
	assign andOp_81_in1 = state_4_is_active;
	// controller for andOp_83.andOp_83_in0
	// controller for andOp_83.andOp_83_in1
	// Insensitive connections
	assign andOp_83_in0 = andOp_81_out;
	assign andOp_83_in1 = data_in_4_55_out_data;
	// controller for andOp_85.andOp_85_in0
	// controller for andOp_85.andOp_85_in1
	// Insensitive connections
	assign andOp_85_in0 = andOp_81_out;
	assign andOp_85_in1 = notOp_84_out;
	// controller for andOp_86.andOp_86_in0
	// controller for andOp_86.andOp_86_in1
	// Insensitive connections
	assign andOp_86_in0 = bb_3_active_in_state_4_out_data;
	assign andOp_86_in1 = state_4_is_active;
	// controller for andOp_88.andOp_88_in0
	// controller for andOp_88.andOp_88_in1
	// Insensitive connections
	assign andOp_88_in0 = andOp_86_out;
	assign andOp_88_in1 = data_in_4_55_out_data;
	// controller for andOp_90.andOp_90_in0
	// controller for andOp_90.andOp_90_in1
	// Insensitive connections
	assign andOp_90_in0 = andOp_86_out;
	assign andOp_90_in1 = notOp_89_out;
	// controller for andOp_91.andOp_91_in0
	// controller for andOp_91.andOp_91_in1
	// Insensitive connections
	assign andOp_91_in0 = bb_3_active_in_state_4_out_data;
	assign andOp_91_in1 = state_4_is_active;
	// controller for andOp_93.andOp_93_in0
	// controller for andOp_93.andOp_93_in1
	// Insensitive connections
	assign andOp_93_in0 = andOp_91_out;
	assign andOp_93_in1 = data_in_4_55_out_data;
	// controller for andOp_95.andOp_95_in0
	// controller for andOp_95.andOp_95_in1
	// Insensitive connections
	assign andOp_95_in0 = andOp_91_out;
	assign andOp_95_in1 = notOp_94_out;
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_98_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_112_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_0.bb_1_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_0_in_data = orOp_100_out;
		end else begin
			bb_1_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_0.bb_1_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_115_out) begin 
			bb_1_predecessor_in_state_0_in_data = 32'd0;
		end else if (eq_113_out) begin 
			bb_1_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_4.bb_2_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_4_in_data = orOp_107_out;
		end else begin
			bb_2_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_4.bb_2_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_124_out) begin 
			bb_2_predecessor_in_state_4_in_data = 32'd3;
		end else if (eq_122_out) begin 
			bb_2_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_1.bb_3_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_1_in_data = orOp_103_out;
		end else begin
			bb_3_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_2.bb_3_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_2_in_data = eq_104_out;
		end else begin
			bb_3_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_3.bb_3_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_3_in_data = eq_105_out;
		end else begin
			bb_3_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_4.bb_3_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_4_in_data = eq_108_out;
		end else begin
			bb_3_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_1.bb_3_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_119_out) begin 
			bb_3_predecessor_in_state_1_in_data = 32'd4;
		end else if (eq_117_out) begin 
			bb_3_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_2.bb_3_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_120_out) begin 
			bb_3_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_3.bb_3_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_121_out) begin 
			bb_3_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_4.bb_3_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_125_out) begin 
			bb_3_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_0.bb_4_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_0_in_data = orOp_97_out;
		end else begin
			bb_4_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_1.bb_4_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_1_in_data = eq_101_out;
		end else begin
			bb_4_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_0.bb_4_predecessor_in_state_0_in_data
	always @(*) begin
		if (andOp_111_out) begin 
			bb_4_predecessor_in_state_0_in_data = 32'd1;
		end else if (eq_109_out) begin 
			bb_4_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_1.bb_4_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_116_out) begin 
			bb_4_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_67_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_68_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_1_happened_in_state_0.br_1_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_69_out) begin 
			br_1_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_70_out) begin 
			br_1_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_1_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_1.br_3_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_76_out) begin 
			br_3_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_77_out) begin 
			br_3_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_2.br_3_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_81_out) begin 
			br_3_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_82_out) begin 
			br_3_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_3.br_3_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_86_out) begin 
			br_3_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_87_out) begin 
			br_3_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_4.br_3_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_91_out) begin 
			br_3_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_92_out) begin 
			br_3_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_0.br_4_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_62_out) begin 
			br_4_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_63_out) begin 
			br_4_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_1.br_4_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_71_out) begin 
			br_4_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_72_out) begin 
			br_4_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_1_in_data = 0;
		end
	end
	// controller for concat_139.concat_139_in0
	// controller for concat_139.concat_139_in1
	// Insensitive connections
	assign concat_139_in0 = data_in_0_9_out_data;
	assign concat_139_in1 = 32'd0;
	// controller for concat_140.concat_140_in0
	// controller for concat_140.concat_140_in1
	// Insensitive connections
	assign concat_140_in0 = 32'd3;
	assign concat_140_in1 = 32'd0;
	// controller for concat_142.concat_142_in0
	// controller for concat_142.concat_142_in1
	// Insensitive connections
	assign concat_142_in0 = data_in_0_12_out_data;
	assign concat_142_in1 = 32'd0;
	// controller for concat_143.concat_143_in0
	// controller for concat_143.concat_143_in1
	// Insensitive connections
	assign concat_143_in0 = 32'd4;
	assign concat_143_in1 = 32'd1;
	// controller for concat_145.concat_145_in0
	// controller for concat_145.concat_145_in1
	// Insensitive connections
	assign concat_145_in0 = data_in_0_10_out_data;
	assign concat_145_in1 = 32'd0;
	// controller for concat_146.concat_146_in0
	// controller for concat_146.concat_146_in1
	// Insensitive connections
	assign concat_146_in0 = 32'd4;
	assign concat_146_in1 = 32'd1;
	// controller for data_in_0_10.data_in_0_10_in_data
	always @(*) begin
		if (eq_178_out) begin 
			data_in_0_10_in_data = 32'd0;
		end else if (eq_179_out) begin 
			data_in_0_10_in_data = data_store_1_23;
		end else if (eq_180_out) begin 
			data_in_0_10_in_data = data_store_4_58;
		end else begin
			data_in_0_10_in_data = 0;
		end
	end
	// controller for data_in_0_12.data_in_0_12_in_data
	always @(*) begin
		if (eq_178_out) begin 
			data_in_0_12_in_data = data_store_0_11;
		end else if (eq_179_out) begin 
			data_in_0_12_in_data = data_store_1_24;
		end else if (eq_180_out) begin 
			data_in_0_12_in_data = data_store_4_60;
		end else begin
			data_in_0_12_in_data = 0;
		end
	end
	// controller for data_in_0_2.data_in_0_2_in_data
	always @(*) begin
		if (eq_178_out) begin 
			data_in_0_2_in_data = data_store_0_1;
		end else if (eq_179_out) begin 
			data_in_0_2_in_data = data_store_1_14;
		end else if (eq_180_out) begin 
			data_in_0_2_in_data = data_store_4_50;
		end else begin
			data_in_0_2_in_data = 0;
		end
	end
	// controller for data_in_0_4.data_in_0_4_in_data
	always @(*) begin
		if (eq_178_out) begin 
			data_in_0_4_in_data = data_store_0_3;
		end else if (eq_179_out) begin 
			data_in_0_4_in_data = data_store_1_16;
		end else if (eq_180_out) begin 
			data_in_0_4_in_data = data_store_4_52;
		end else begin
			data_in_0_4_in_data = 0;
		end
	end
	// controller for data_in_0_6.data_in_0_6_in_data
	always @(*) begin
		if (eq_178_out) begin 
			data_in_0_6_in_data = data_store_0_5;
		end else if (eq_179_out) begin 
			data_in_0_6_in_data = data_store_1_18;
		end else if (eq_180_out) begin 
			data_in_0_6_in_data = data_store_4_54;
		end else begin
			data_in_0_6_in_data = 0;
		end
	end
	// controller for data_in_0_9.data_in_0_9_in_data
	always @(*) begin
		if (eq_178_out) begin 
			data_in_0_9_in_data = data_store_0_8;
		end else if (eq_179_out) begin 
			data_in_0_9_in_data = data_store_1_21;
		end else if (eq_180_out) begin 
			data_in_0_9_in_data = data_store_4_56;
		end else begin
			data_in_0_9_in_data = 0;
		end
	end
	// controller for data_in_1_13.data_in_1_13_in_data
	always @(*) begin
		if (eq_186_out) begin 
			data_in_1_13_in_data = data_store_0_0;
		end else if (eq_187_out) begin 
			data_in_1_13_in_data = 1'd0;
		end else begin
			data_in_1_13_in_data = 0;
		end
	end
	// controller for data_in_1_15.data_in_1_15_in_data
	always @(*) begin
		if (eq_186_out) begin 
			data_in_1_15_in_data = data_store_0_1;
		end else if (eq_187_out) begin 
			data_in_1_15_in_data = data_store_1_14;
		end else begin
			data_in_1_15_in_data = 0;
		end
	end
	// controller for data_in_1_17.data_in_1_17_in_data
	always @(*) begin
		if (eq_186_out) begin 
			data_in_1_17_in_data = data_store_0_3;
		end else if (eq_187_out) begin 
			data_in_1_17_in_data = data_store_1_16;
		end else begin
			data_in_1_17_in_data = 0;
		end
	end
	// controller for data_in_1_19.data_in_1_19_in_data
	always @(*) begin
		if (eq_186_out) begin 
			data_in_1_19_in_data = data_store_0_5;
		end else if (eq_187_out) begin 
			data_in_1_19_in_data = data_store_1_18;
		end else begin
			data_in_1_19_in_data = 0;
		end
	end
	// controller for data_in_1_20.data_in_1_20_in_data
	always @(*) begin
		if (eq_186_out) begin 
			data_in_1_20_in_data = data_store_0_7;
		end else if (eq_187_out) begin 
			data_in_1_20_in_data = 32'd0;
		end else begin
			data_in_1_20_in_data = 0;
		end
	end
	// controller for data_in_1_22.data_in_1_22_in_data
	always @(*) begin
		if (eq_186_out) begin 
			data_in_1_22_in_data = data_store_0_8;
		end else if (eq_187_out) begin 
			data_in_1_22_in_data = data_store_1_21;
		end else begin
			data_in_1_22_in_data = 0;
		end
	end
	// controller for data_in_1_25.data_in_1_25_in_data
	always @(*) begin
		if (eq_186_out) begin 
			data_in_1_25_in_data = data_store_0_11;
		end else if (eq_187_out) begin 
			data_in_1_25_in_data = data_store_1_24;
		end else begin
			data_in_1_25_in_data = 0;
		end
	end
	// controller for data_in_2_27.data_in_2_27_in_data
	always @(*) begin
		if (eq_191_out) begin 
			data_in_2_27_in_data = data_store_1_14;
		end else if (eq_192_out) begin 
			data_in_2_27_in_data = data_store_2_26;
		end else begin
			data_in_2_27_in_data = 0;
		end
	end
	// controller for data_in_2_29.data_in_2_29_in_data
	always @(*) begin
		if (eq_191_out) begin 
			data_in_2_29_in_data = data_store_1_16;
		end else if (eq_192_out) begin 
			data_in_2_29_in_data = data_store_2_28;
		end else begin
			data_in_2_29_in_data = 0;
		end
	end
	// controller for data_in_2_31.data_in_2_31_in_data
	always @(*) begin
		if (eq_191_out) begin 
			data_in_2_31_in_data = data_store_1_18;
		end else if (eq_192_out) begin 
			data_in_2_31_in_data = data_store_2_30;
		end else begin
			data_in_2_31_in_data = 0;
		end
	end
	// controller for data_in_2_33.data_in_2_33_in_data
	always @(*) begin
		if (eq_191_out) begin 
			data_in_2_33_in_data = data_store_1_21;
		end else if (eq_192_out) begin 
			data_in_2_33_in_data = data_store_2_32;
		end else begin
			data_in_2_33_in_data = 0;
		end
	end
	// controller for data_in_2_35.data_in_2_35_in_data
	always @(*) begin
		if (eq_191_out) begin 
			data_in_2_35_in_data = data_store_1_23;
		end else if (eq_192_out) begin 
			data_in_2_35_in_data = data_store_2_34;
		end else begin
			data_in_2_35_in_data = 0;
		end
	end
	// controller for data_in_2_37.data_in_2_37_in_data
	always @(*) begin
		if (eq_191_out) begin 
			data_in_2_37_in_data = data_store_1_24;
		end else if (eq_192_out) begin 
			data_in_2_37_in_data = data_store_2_36;
		end else begin
			data_in_2_37_in_data = 0;
		end
	end
	// controller for data_in_3_39.data_in_3_39_in_data
	always @(*) begin
		if (eq_193_out) begin 
			data_in_3_39_in_data = data_store_2_26;
		end else if (eq_194_out) begin 
			data_in_3_39_in_data = data_store_3_38;
		end else begin
			data_in_3_39_in_data = 0;
		end
	end
	// controller for data_in_3_41.data_in_3_41_in_data
	always @(*) begin
		if (eq_193_out) begin 
			data_in_3_41_in_data = data_store_2_28;
		end else if (eq_194_out) begin 
			data_in_3_41_in_data = data_store_3_40;
		end else begin
			data_in_3_41_in_data = 0;
		end
	end
	// controller for data_in_3_43.data_in_3_43_in_data
	always @(*) begin
		if (eq_193_out) begin 
			data_in_3_43_in_data = data_store_2_30;
		end else if (eq_194_out) begin 
			data_in_3_43_in_data = data_store_3_42;
		end else begin
			data_in_3_43_in_data = 0;
		end
	end
	// controller for data_in_3_45.data_in_3_45_in_data
	always @(*) begin
		if (eq_193_out) begin 
			data_in_3_45_in_data = data_store_2_32;
		end else if (eq_194_out) begin 
			data_in_3_45_in_data = data_store_3_44;
		end else begin
			data_in_3_45_in_data = 0;
		end
	end
	// controller for data_in_3_47.data_in_3_47_in_data
	always @(*) begin
		if (eq_193_out) begin 
			data_in_3_47_in_data = data_store_2_34;
		end else if (eq_194_out) begin 
			data_in_3_47_in_data = data_store_3_46;
		end else begin
			data_in_3_47_in_data = 0;
		end
	end
	// controller for data_in_3_49.data_in_3_49_in_data
	always @(*) begin
		if (eq_193_out) begin 
			data_in_3_49_in_data = data_store_2_36;
		end else if (eq_194_out) begin 
			data_in_3_49_in_data = data_store_3_48;
		end else begin
			data_in_3_49_in_data = 0;
		end
	end
	// controller for data_in_4_51.data_in_4_51_in_data
	always @(*) begin
		if (eq_195_out) begin 
			data_in_4_51_in_data = data_store_3_38;
		end else if (eq_196_out) begin 
			data_in_4_51_in_data = data_store_4_50;
		end else begin
			data_in_4_51_in_data = 0;
		end
	end
	// controller for data_in_4_53.data_in_4_53_in_data
	always @(*) begin
		if (eq_195_out) begin 
			data_in_4_53_in_data = data_store_3_40;
		end else if (eq_196_out) begin 
			data_in_4_53_in_data = data_store_4_52;
		end else begin
			data_in_4_53_in_data = 0;
		end
	end
	// controller for data_in_4_55.data_in_4_55_in_data
	always @(*) begin
		if (eq_195_out) begin 
			data_in_4_55_in_data = data_store_3_42;
		end else if (eq_196_out) begin 
			data_in_4_55_in_data = data_store_4_54;
		end else begin
			data_in_4_55_in_data = 0;
		end
	end
	// controller for data_in_4_57.data_in_4_57_in_data
	always @(*) begin
		if (eq_195_out) begin 
			data_in_4_57_in_data = data_store_3_44;
		end else if (eq_196_out) begin 
			data_in_4_57_in_data = data_store_4_56;
		end else begin
			data_in_4_57_in_data = 0;
		end
	end
	// controller for data_in_4_59.data_in_4_59_in_data
	always @(*) begin
		if (eq_195_out) begin 
			data_in_4_59_in_data = data_store_3_46;
		end else if (eq_196_out) begin 
			data_in_4_59_in_data = data_store_4_58;
		end else begin
			data_in_4_59_in_data = 0;
		end
	end
	// controller for data_in_4_61.data_in_4_61_in_data
	always @(*) begin
		if (eq_195_out) begin 
			data_in_4_61_in_data = data_store_3_48;
		end else if (eq_196_out) begin 
			data_in_4_61_in_data = data_store_4_60;
		end else begin
			data_in_4_61_in_data = 0;
		end
	end
	// controller for eq_101.eq_101_in0
	// controller for eq_101.eq_101_in1
	// Insensitive connections
	assign eq_101_in0 = 32'd4;
	assign eq_101_in1 = state_1_entry_BB_reg;
	// controller for eq_102.eq_102_in0
	// controller for eq_102.eq_102_in1
	// Insensitive connections
	assign eq_102_in0 = 32'd3;
	assign eq_102_in1 = state_1_entry_BB_reg;
	// controller for eq_104.eq_104_in0
	// controller for eq_104.eq_104_in1
	// Insensitive connections
	assign eq_104_in0 = 32'd3;
	assign eq_104_in1 = state_2_entry_BB_reg;
	// controller for eq_105.eq_105_in0
	// controller for eq_105.eq_105_in1
	// Insensitive connections
	assign eq_105_in0 = 32'd3;
	assign eq_105_in1 = state_3_entry_BB_reg;
	// controller for eq_106.eq_106_in0
	// controller for eq_106.eq_106_in1
	// Insensitive connections
	assign eq_106_in0 = 32'd2;
	assign eq_106_in1 = state_4_entry_BB_reg;
	// controller for eq_108.eq_108_in0
	// controller for eq_108.eq_108_in1
	// Insensitive connections
	assign eq_108_in0 = 32'd3;
	assign eq_108_in1 = state_4_entry_BB_reg;
	// controller for eq_109.eq_109_in0
	// controller for eq_109.eq_109_in1
	// Insensitive connections
	assign eq_109_in0 = 32'd4;
	assign eq_109_in1 = state_0_entry_BB_reg;
	// controller for eq_112.eq_112_in0
	// controller for eq_112.eq_112_in1
	// Insensitive connections
	assign eq_112_in0 = 32'd0;
	assign eq_112_in1 = state_0_entry_BB_reg;
	// controller for eq_113.eq_113_in0
	// controller for eq_113.eq_113_in1
	// Insensitive connections
	assign eq_113_in0 = 32'd1;
	assign eq_113_in1 = state_0_entry_BB_reg;
	// controller for eq_116.eq_116_in0
	// controller for eq_116.eq_116_in1
	// Insensitive connections
	assign eq_116_in0 = 32'd4;
	assign eq_116_in1 = state_1_entry_BB_reg;
	// controller for eq_117.eq_117_in0
	// controller for eq_117.eq_117_in1
	// Insensitive connections
	assign eq_117_in0 = 32'd3;
	assign eq_117_in1 = state_1_entry_BB_reg;
	// controller for eq_120.eq_120_in0
	// controller for eq_120.eq_120_in1
	// Insensitive connections
	assign eq_120_in0 = 32'd3;
	assign eq_120_in1 = state_2_entry_BB_reg;
	// controller for eq_121.eq_121_in0
	// controller for eq_121.eq_121_in1
	// Insensitive connections
	assign eq_121_in0 = 32'd3;
	assign eq_121_in1 = state_3_entry_BB_reg;
	// controller for eq_122.eq_122_in0
	// controller for eq_122.eq_122_in1
	// Insensitive connections
	assign eq_122_in0 = 32'd2;
	assign eq_122_in1 = state_4_entry_BB_reg;
	// controller for eq_125.eq_125_in0
	// controller for eq_125.eq_125_in1
	// Insensitive connections
	assign eq_125_in0 = 32'd3;
	assign eq_125_in1 = state_4_entry_BB_reg;
	// controller for eq_134.eq_134_in0
	// controller for eq_134.eq_134_in1
	// Insensitive connections
	assign eq_134_in0 = 32'd4;
	assign eq_134_in1 = state_1_entry_BB_reg;
	// controller for eq_149.eq_149_in0
	// controller for eq_149.eq_149_in1
	// Insensitive connections
	assign eq_149_in0 = 32'd4;
	assign eq_149_in1 = state_0_entry_BB_reg;
	// controller for eq_150.eq_150_in0
	// controller for eq_150.eq_150_in1
	// Insensitive connections
	assign eq_150_in0 = 32'd0;
	assign eq_150_in1 = state_0_entry_BB_reg;
	// controller for eq_151.eq_151_in0
	// controller for eq_151.eq_151_in1
	// Insensitive connections
	assign eq_151_in0 = 32'd1;
	assign eq_151_in1 = state_0_entry_BB_reg;
	// controller for eq_178.eq_178_in0
	// controller for eq_178.eq_178_in1
	// Insensitive connections
	assign eq_178_in0 = 32'd0;
	assign eq_178_in1 = state_0_last_state;
	// controller for eq_179.eq_179_in0
	// controller for eq_179.eq_179_in1
	// Insensitive connections
	assign eq_179_in0 = 32'd1;
	assign eq_179_in1 = state_0_last_state;
	// controller for eq_180.eq_180_in0
	// controller for eq_180.eq_180_in1
	// Insensitive connections
	assign eq_180_in0 = 32'd4;
	assign eq_180_in1 = state_0_last_state;
	// controller for eq_186.eq_186_in0
	// controller for eq_186.eq_186_in1
	// Insensitive connections
	assign eq_186_in0 = 32'd0;
	assign eq_186_in1 = state_1_last_state;
	// controller for eq_187.eq_187_in0
	// controller for eq_187.eq_187_in1
	// Insensitive connections
	assign eq_187_in0 = 32'd1;
	assign eq_187_in1 = state_1_last_state;
	// controller for eq_191.eq_191_in0
	// controller for eq_191.eq_191_in1
	// Insensitive connections
	assign eq_191_in0 = 32'd1;
	assign eq_191_in1 = state_2_last_state;
	// controller for eq_192.eq_192_in0
	// controller for eq_192.eq_192_in1
	// Insensitive connections
	assign eq_192_in0 = 32'd2;
	assign eq_192_in1 = state_2_last_state;
	// controller for eq_193.eq_193_in0
	// controller for eq_193.eq_193_in1
	// Insensitive connections
	assign eq_193_in0 = 32'd2;
	assign eq_193_in1 = state_3_last_state;
	// controller for eq_194.eq_194_in0
	// controller for eq_194.eq_194_in1
	// Insensitive connections
	assign eq_194_in0 = 32'd3;
	assign eq_194_in1 = state_3_last_state;
	// controller for eq_195.eq_195_in0
	// controller for eq_195.eq_195_in1
	// Insensitive connections
	assign eq_195_in0 = 32'd3;
	assign eq_195_in1 = state_4_last_state;
	// controller for eq_196.eq_196_in0
	// controller for eq_196.eq_196_in1
	// Insensitive connections
	assign eq_196_in0 = 32'd4;
	assign eq_196_in1 = state_4_last_state;
	// controller for eq_96.eq_96_in0
	// controller for eq_96.eq_96_in1
	// Insensitive connections
	assign eq_96_in0 = 32'd4;
	assign eq_96_in1 = state_0_entry_BB_reg;
	// controller for eq_98.eq_98_in0
	// controller for eq_98.eq_98_in1
	// Insensitive connections
	assign eq_98_in0 = 32'd0;
	assign eq_98_in1 = state_0_entry_BB_reg;
	// controller for eq_99.eq_99_in0
	// controller for eq_99.eq_99_in1
	// Insensitive connections
	assign eq_99_in0 = 32'd1;
	assign eq_99_in1 = state_0_entry_BB_reg;
	// controller for icmp_icmp0.icmp_icmp0_in0
	// controller for icmp_icmp0.icmp_icmp0_in1
	// Insensitive connections
	assign icmp_icmp0_in0 = add_add10_out;
	assign icmp_icmp0_in1 = 32'd3;
	// controller for icmp_icmp16.icmp_icmp16_in0
	// controller for icmp_icmp16.icmp_icmp16_in1
	// Insensitive connections
	assign icmp_icmp16_in0 = add_add17_out;
	assign icmp_icmp16_in1 = 32'd3;
	// controller for mul_mul1.mul_mul1_in0
	// controller for mul_mul1.mul_mul1_in1
	// Insensitive connections
	assign mul_mul1_in0 = phi_phi5_out;
	assign mul_mul1_in1 = 32'd3;
	// controller for mul_mul14.mul_mul14_in0
	// controller for mul_mul14.mul_mul14_in1
	// Insensitive connections
	assign mul_mul14_in0 = ram_rdata_2;
	assign mul_mul14_in1 = ram_rdata_1;
	// controller for notOp_110.notOp_110_in0
	// Insensitive connections
	assign notOp_110_in0 = eq_109_out;
	// controller for notOp_114.notOp_114_in0
	// Insensitive connections
	assign notOp_114_in0 = eq_113_out;
	// controller for notOp_118.notOp_118_in0
	// Insensitive connections
	assign notOp_118_in0 = eq_117_out;
	// controller for notOp_123.notOp_123_in0
	// Insensitive connections
	assign notOp_123_in0 = eq_122_out;
	// controller for notOp_164.notOp_164_in0
	// Insensitive connections
	assign notOp_164_in0 = andOp_66_out;
	// controller for notOp_166.notOp_166_in0
	// Insensitive connections
	assign notOp_166_in0 = andOp_80_out;
	// controller for notOp_168.notOp_168_in0
	// Insensitive connections
	assign notOp_168_in0 = andOp_159_out;
	// controller for notOp_170.notOp_170_in0
	// Insensitive connections
	assign notOp_170_in0 = andOp_160_out;
	// controller for notOp_172.notOp_172_in0
	// Insensitive connections
	assign notOp_172_in0 = andOp_161_out;
	// controller for notOp_174.notOp_174_in0
	// Insensitive connections
	assign notOp_174_in0 = andOp_162_out;
	// controller for notOp_176.notOp_176_in0
	// Insensitive connections
	assign notOp_176_in0 = andOp_163_out;
	// controller for notOp_63.notOp_63_in0
	// Insensitive connections
	assign notOp_63_in0 = andOp_62_out;
	// controller for notOp_65.notOp_65_in0
	// Insensitive connections
	assign notOp_65_in0 = data_in_1_13_out_data;
	// controller for notOp_68.notOp_68_in0
	// Insensitive connections
	assign notOp_68_in0 = andOp_67_out;
	// controller for notOp_70.notOp_70_in0
	// Insensitive connections
	assign notOp_70_in0 = andOp_69_out;
	// controller for notOp_72.notOp_72_in0
	// Insensitive connections
	assign notOp_72_in0 = andOp_71_out;
	// controller for notOp_74.notOp_74_in0
	// Insensitive connections
	assign notOp_74_in0 = data_in_1_13_out_data;
	// controller for notOp_77.notOp_77_in0
	// Insensitive connections
	assign notOp_77_in0 = andOp_76_out;
	// controller for notOp_79.notOp_79_in0
	// Insensitive connections
	assign notOp_79_in0 = data_in_4_55_out_data;
	// controller for notOp_82.notOp_82_in0
	// Insensitive connections
	assign notOp_82_in0 = andOp_81_out;
	// controller for notOp_84.notOp_84_in0
	// Insensitive connections
	assign notOp_84_in0 = data_in_4_55_out_data;
	// controller for notOp_87.notOp_87_in0
	// Insensitive connections
	assign notOp_87_in0 = andOp_86_out;
	// controller for notOp_89.notOp_89_in0
	// Insensitive connections
	assign notOp_89_in0 = data_in_4_55_out_data;
	// controller for notOp_92.notOp_92_in0
	// Insensitive connections
	assign notOp_92_in0 = andOp_91_out;
	// controller for notOp_94.notOp_94_in0
	// Insensitive connections
	assign notOp_94_in0 = data_in_4_55_out_data;
	// controller for orOp_100.orOp_100_in0
	// controller for orOp_100.orOp_100_in1
	// Insensitive connections
	assign orOp_100_in0 = eq_99_out;
	assign orOp_100_in1 = andOp_67_out;
	// controller for orOp_103.orOp_103_in0
	// controller for orOp_103.orOp_103_in1
	// Insensitive connections
	assign orOp_103_in0 = eq_102_out;
	assign orOp_103_in1 = andOp_64_out;
	// controller for orOp_107.orOp_107_in0
	// controller for orOp_107.orOp_107_in1
	// Insensitive connections
	assign orOp_107_in0 = eq_106_out;
	assign orOp_107_in1 = andOp_78_out;
	// controller for orOp_97.orOp_97_in0
	// controller for orOp_97.orOp_97_in1
	// Insensitive connections
	assign orOp_97_in0 = eq_96_out;
	assign orOp_97_in1 = andOp_69_out;
	// controller for phi_phi5.phi_phi5_in
	// controller for phi_phi5.phi_phi5_last_block
	// controller for phi_phi5.phi_phi5_s
	// Insensitive connections
	assign phi_phi5_in = concat_139_out;
	assign phi_phi5_last_block = bb_1_predecessor_in_state_0_out_data;
	assign phi_phi5_s = concat_140_out;
	// controller for phi_phi6.phi_phi6_in
	// controller for phi_phi6.phi_phi6_last_block
	// controller for phi_phi6.phi_phi6_s
	// Insensitive connections
	assign phi_phi6_in = concat_142_out;
	assign phi_phi6_last_block = bb_4_predecessor_in_state_0_out_data;
	assign phi_phi6_s = concat_143_out;
	// controller for phi_phi7.phi_phi7_in
	// controller for phi_phi7.phi_phi7_last_block
	// controller for phi_phi7.phi_phi7_s
	// Insensitive connections
	assign phi_phi7_in = concat_145_out;
	assign phi_phi7_last_block = bb_4_predecessor_in_state_0_out_data;
	assign phi_phi7_s = concat_146_out;
	// controller for ram.ram_raddr_1_reg
	always @(*) begin
		if (andOp_128_out) begin 
			ram_raddr_1_reg = add_add8_out;
		end else begin
			ram_raddr_1_reg = 0;
		end
	end
	// controller for ram.ram_raddr_2_reg
	always @(*) begin
		if (andOp_129_out) begin 
			ram_raddr_2_reg = add_add3_out;
		end else begin
			ram_raddr_2_reg = 0;
		end
	end
	// controller for ram.ram_waddr_0_reg
	always @(*) begin
		if (andOp_136_out) begin 
			ram_waddr_0_reg = add_add12_out;
		end else begin
			ram_waddr_0_reg = 0;
		end
	end
	// controller for ram.ram_wdata_0_reg
	always @(*) begin
		if (andOp_132_out) begin 
			ram_wdata_0_reg = tmp_output_133_out_data;
		end else begin
			ram_wdata_0_reg = 0;
		end
	end
	// controller for ram.ram_wen_0_reg
	always @(*) begin
		if (andOp_135_out) begin 
			ram_wen_0_reg = -(1'd1);
		end else begin
			ram_wen_0_reg = 0;
		end
	end
	// controller for ret23.valid_reg
	always @(*) begin
		if (andOp_158_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// controller for tmp_output_133.tmp_output_133_in_data
	always @(*) begin
		if (eq_134_out) begin 
			tmp_output_133_in_data = add_add21_out;
		end else begin
			tmp_output_133_in_data = 0;
		end
	end
	// controller for tmp_output_148.tmp_output_148_in_data
	always @(*) begin
		if (eq_149_out) begin 
			tmp_output_148_in_data = data_in_0_2_out_data;
		end else if (eq_150_out) begin 
			tmp_output_148_in_data = mul_mul1_out;
		end else if (eq_151_out) begin 
			tmp_output_148_in_data = mul_mul1_out;
		end else begin
			tmp_output_148_in_data = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			data_store_0_0 <= 0;
		end else begin
			if (andOp_181_out) begin
				data_store_0_0 <= icmp_icmp0_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_1 <= 0;
		end else begin
			if (andOp_182_out) begin
				data_store_0_1 <= mul_mul1_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_11 <= 0;
		end else begin
			if (andOp_185_out) begin
				data_store_0_11 <= add_add10_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_3 <= 0;
		end else begin
			if (andOp_183_out) begin
				data_store_0_3 <= phi_phi5_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_5 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_5 <= data_in_0_6_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_7 <= 0;
		end else begin
			if (andOp_184_out) begin
				data_store_0_7 <= phi_phi7_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_8 <= 0;
		end else begin
			if (state_0_is_active) begin
				data_store_0_8 <= data_in_0_9_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_14 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_14 <= data_in_1_15_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_16 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_16 <= data_in_1_17_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_18 <= 0;
		end else begin
			if (andOp_188_out) begin
				data_store_1_18 <= icmp_icmp16_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_21 <= 0;
		end else begin
			if (andOp_189_out) begin
				data_store_1_21 <= add_add17_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_23 <= 0;
		end else begin
			if (andOp_190_out) begin
				data_store_1_23 <= add_add21_out;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_24 <= 0;
		end else begin
			if (state_1_is_active) begin
				data_store_1_24 <= data_in_1_25_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_26 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_26 <= data_in_2_27_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_28 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_28 <= data_in_2_29_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_30 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_30 <= data_in_2_31_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_32 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_32 <= data_in_2_33_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_34 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_34 <= data_in_2_35_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_36 <= 0;
		end else begin
			if (state_2_is_active) begin
				data_store_2_36 <= data_in_2_37_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_38 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_38 <= data_in_3_39_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_40 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_40 <= data_in_3_41_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_42 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_42 <= data_in_3_43_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_44 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_44 <= data_in_3_45_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_46 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_46 <= data_in_3_47_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_48 <= 0;
		end else begin
			if (state_3_is_active) begin
				data_store_3_48 <= data_in_3_49_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_50 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_50 <= data_in_4_51_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_52 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_52 <= data_in_4_53_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_54 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_54 <= data_in_4_55_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_56 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_56 <= data_in_4_57_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_58 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_58 <= data_in_4_59_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_60 <= 0;
		end else begin
			if (state_4_is_active) begin
				data_store_4_60 <= data_in_4_61_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_159_out) begin
				global_state <= 32'd1;
			end
			if (andOp_160_out) begin
				global_state <= 32'd2;
			end
			if (andOp_161_out) begin
				global_state <= 32'd3;
			end
			if (andOp_162_out) begin
				global_state <= 32'd4;
			end
			if (andOp_163_out) begin
				global_state <= 32'd4;
			end
			if (andOp_66_out) begin
				global_state <= 32'd0;
			end
			if (andOp_80_out) begin
				global_state <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
			if (andOp_66_out) begin
				state_0_entry_BB_reg <= 32'd4;
			end
			if (andOp_80_out) begin
				state_0_entry_BB_reg <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (andOp_167_out) begin
				state_0_is_active <= 1'd0;
			end
			if (andOp_66_out) begin
				state_0_is_active <= 1'd1;
			end
			if (andOp_80_out) begin
				state_0_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
			if (andOp_66_out) begin
				state_0_last_BB_reg <= 32'd4;
			end
			if (andOp_80_out) begin
				state_0_last_BB_reg <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
			if (andOp_66_out) begin
				state_0_last_state <= 32'd1;
			end
			if (andOp_80_out) begin
				state_0_last_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_159_out) begin
				state_1_entry_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_159_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_169_out) begin
				state_1_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_159_out) begin
				state_1_last_BB_reg <= bb_4_predecessor_in_state_0_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_159_out) begin
				state_1_last_state <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_160_out) begin
				state_2_entry_BB_reg <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_160_out) begin
				state_2_is_active <= 1'd1;
			end
			if (andOp_171_out) begin
				state_2_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_160_out) begin
				state_2_last_BB_reg <= bb_3_predecessor_in_state_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_160_out) begin
				state_2_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_161_out) begin
				state_3_entry_BB_reg <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_161_out) begin
				state_3_is_active <= 1'd1;
			end
			if (andOp_173_out) begin
				state_3_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_161_out) begin
				state_3_last_BB_reg <= bb_3_predecessor_in_state_2_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_state <= 0;
		end else begin
			if (andOp_161_out) begin
				state_3_last_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_162_out) begin
				state_4_entry_BB_reg <= 32'd3;
			end
			if (andOp_163_out) begin
				state_4_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_162_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_163_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_177_out) begin
				state_4_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_162_out) begin
				state_4_last_BB_reg <= bb_3_predecessor_in_state_3_out_data;
			end
			if (andOp_163_out) begin
				state_4_last_BB_reg <= bb_2_predecessor_in_state_4_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_state <= 0;
		end else begin
			if (andOp_162_out) begin
				state_4_last_state <= 32'd3;
			end
			if (andOp_163_out) begin
				state_4_last_state <= 32'd4;
			end
		end
	end

endmodule

