module channel_reduce_4_inner(input [0:0] clk, input [0:0] rst, output [31:0] out_in_data, output [0:0] out_read_valid, output [0:0] out_rst, output [31:0] out_write_valid, input [31:0] out_out_data, input [0:0] out_read_ready, input [0:0] out_write_ready, output [0:0] valid, output [31:0] in_in_data, output [0:0] in_read_valid, output [0:0] in_rst, output [31:0] in_write_valid, input [31:0] in_out_data, input [0:0] in_read_ready, input [0:0] in_write_ready);

	reg [31:0] out_in_data_reg;
	reg [0:0] out_read_valid_reg;
	reg [0:0] out_rst_reg;
	reg [31:0] out_write_valid_reg;
	reg [0:0] valid_reg;
	reg [31:0] in_in_data_reg;
	reg [0:0] in_read_valid_reg;
	reg [0:0] in_rst_reg;
	reg [31:0] in_write_valid_reg;

	assign out_in_data = out_in_data_reg;
	assign out_read_valid = out_read_valid_reg;
	assign out_rst = out_rst_reg;
	assign out_write_valid = out_write_valid_reg;
	assign valid = valid_reg;
	assign in_in_data = in_in_data_reg;
	assign in_read_valid = in_read_valid_reg;
	assign in_rst = in_rst_reg;
	assign in_write_valid = in_write_valid_reg;

	// Start debug wires and ports

	initial begin
	end





	// End debug wires and ports

	// Start Functional Units
	add call_18();

	reg [31:0] raddr_ram_0_reg;
	reg [31:0] waddr_ram_0_reg;
	reg [31:0] wdata_ram_0_reg;
	reg [0:0] wen_ram_0_reg;
	wire [31:0] rdata_ram_0;
	register #(.WIDTH(32)) ram_0(.clk(clk), .raddr(raddr_ram_0_reg), .rdata(rdata_ram_0), .rst(rst), .waddr(waddr_ram_0_reg), .wdata(wdata_ram_0_reg), .wen(wen_ram_0_reg));

	add alloca_0();

	add bitcast_1();

	add call_2();

	br_dummy br_unit();

	add call_19();

	reg [63:0] phi_in_phi_5;
	reg [31:0] phi_last_block_phi_5;
	reg [63:0] phi_s_phi_5;
	wire [31:0] phi_out_phi_5;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_5(.in(phi_in_phi_5), .last_block(phi_last_block_phi_5), .out(phi_out_phi_5), .s(phi_s_phi_5));

	reg [31:0] add_in0_add_12;
	reg [31:0] add_in1_add_12;
	wire [31:0] add_out_add_12;
	add #(.WIDTH(32)) add_add_12(.in0(add_in0_add_12), .in1(add_in1_add_12), .out(add_out_add_12));

	reg [31:0] add_in0_add_7;
	reg [31:0] add_in1_add_7;
	wire [31:0] add_out_add_7;
	add #(.WIDTH(32)) add_add_7(.in0(add_in0_add_7), .in1(add_in1_add_7), .out(add_out_add_7));

	reg [31:0] cmp_in0_icmp_8;
	reg [31:0] cmp_in1_icmp_8;
	wire [0:0] cmp_out_icmp_8;
	eq #(.WIDTH(32)) icmp_8(.in0(cmp_in0_icmp_8), .in1(cmp_in1_icmp_8), .out(cmp_out_icmp_8));

	add call_10();

	// End Functional Units

	// Start instruction result storage
	reg [31:0] load_tmp_1;
	reg [31:0] add_tmp_2;
	reg [0:0] icmp_tmp_3;
	// End instruction result storage

	// Start pipeline variables
	// End pipeline variables

	reg [31:0] global_state;
	reg [31:0] last_BB_reg;
	// Start pipeline reset block
	always @(posedge clk) begin
		if (rst) begin
		end
	end
	// End pipeline reset block

	// Start pipeline valid chain block
	always @(posedge clk) begin

		if (!rst) begin
		end
	end
	// End pipeline valid chain block

	always @(posedge clk) begin
	end
	// Start pipeline initiation block
	always @(posedge clk) begin
	end
	// End pipeline initiation block

	always @(posedge clk) begin
		if (rst) begin
			last_BB_reg <= 0;
		end else begin
			if ((global_state == 0)) begin
			end
			if ((global_state == 1)) begin
					last_BB_reg <= 0;
			end
			if ((global_state == 2)) begin
			end
			if ((global_state == 3)) begin
			end
			if ((global_state == 4)) begin
			end
			if ((global_state == 5)) begin
					last_BB_reg <= 2;
			end
			if ((global_state == 6)) begin
			end
			if ((global_state == 7)) begin
			end
			if ((global_state == 8)) begin
					last_BB_reg <= 1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			// Control code
			if ((global_state == 0)) begin 
				// Next state transition logic
				// Condition = True

				if (1) begin
					global_state <= 1;
				end
			end
			if ((global_state == 1)) begin 
				// Next state transition logic
				// Condition = True

				if (1) begin
					global_state <= 2;
				end
			end
			if ((global_state == 2)) begin 
				// Next state transition logic
				// Condition = True

				if (1) begin
				if (in_read_ready) begin 
					global_state <= 3;
				end
				end
			end
			if ((global_state == 3)) begin 
				// Next state transition logic
				// Condition = True

				if (1) begin
					global_state <= 4;
				end
			end
			if ((global_state == 4)) begin 
				// Next state transition logic
				// Condition = True

				if (1) begin
					global_state <= 5;
				end
			end
			if ((global_state == 5)) begin 
				// Next state transition logic
				// Condition = (  %exitcond = icmp eq i32 %10, 4)
				if ((icmp_tmp_3)) begin
					global_state <= 6;
				end
				// Condition = (!(  %exitcond = icmp eq i32 %10, 4))
				if (!(icmp_tmp_3)) begin
					global_state <= 2;
				end
			end
			if ((global_state == 6)) begin 
				// Next state transition logic
				// Condition = True

				if (1) begin
				if (out_write_ready) begin 
					global_state <= 7;
				end
				end
			end
			if ((global_state == 7)) begin 
				// Next state transition logic
				// Condition = True

				if (1) begin
					global_state <= 8;
				end
			end
			if ((global_state == 8)) begin 
				// Next state transition logic
				// Condition = True

				if (1) begin
					global_state <= 8;
				end
			end

			// Temporary storage code
			if ((global_state == 0)) begin 
				// Temporary storage
				// Store data computed at the stage
			end
			if ((global_state == 1)) begin 
				// Temporary storage
				// Store data computed at the stage
			end
			if ((global_state == 2)) begin 
				// Temporary storage
				if (in_read_ready) begin
				// Store data computed at the stage
					load_tmp_1 <= rdata_ram_0;
					add_tmp_2 <= add_out_add_7;
					icmp_tmp_3 <= cmp_out_icmp_8;
				end
			end
			if ((global_state == 3)) begin 
				// Temporary storage
				// Store data computed at the stage
			end
			if ((global_state == 4)) begin 
				// Temporary storage
				// Store data computed at the stage
			end
			if ((global_state == 5)) begin 
				// Temporary storage
				// Store data computed at the stage
			end
			if ((global_state == 6)) begin 
				// Temporary storage
				if (out_write_ready) begin
				// Store data computed at the stage
				end
			end
			if ((global_state == 7)) begin 
				// Temporary storage
				// Store data computed at the stage
			end
			if ((global_state == 8)) begin 
				// Temporary storage
				// Store data computed at the stage
			end
		end
	end


	// Start pipeline instruction code
	// Start pipeline stages
	// End pipeline instruction code

	// controller for ram_0.raddr_ram_0_reg
	always @(*) begin
		if ((global_state == 2)) begin 
				if (in_read_ready) begin
					raddr_ram_0_reg = 0;
				end
		end
		if ((global_state == 7)) begin 
				if (1) begin
					raddr_ram_0_reg = 0;
				end
		end
		else
		end
	// controller for ram_0.waddr_ram_0_reg
	always @(*) begin
		if ((global_state == 0)) begin 
				if (1) begin
					waddr_ram_0_reg = 0;
				end
		end
		if ((global_state == 4)) begin 
				if (1) begin
					waddr_ram_0_reg = 0;
				end
		end
		else
		end
	// controller for ram_0.wdata_ram_0_reg
	always @(*) begin
		if ((global_state == 0)) begin 
				if (1) begin
					wdata_ram_0_reg = (32'd0);
				end
		end
		if ((global_state == 4)) begin 
				if (1) begin
					wdata_ram_0_reg = add_out_add_12;
				end
		end
		else
		end
	// controller for ram_0.wen_ram_0_reg
	always @(*) begin
		if ((global_state == 0)) begin 
				if (1) begin
					wen_ram_0_reg = 1;
				end
		end
		if ((global_state == 4)) begin 
				if (1) begin
					wen_ram_0_reg = 1;
				end
		end
		else
		end
	// controller for phi_5.phi_in_phi_5
	always @(*) begin
		if ((global_state == 2)) begin 
				if (in_read_ready) begin
					phi_in_phi_5 = {(32'd0), add_tmp_2};
				end
		end
		else
		end
	// controller for phi_5.phi_last_block_phi_5
	always @(*) begin
		if ((global_state == 2)) begin 
				if (in_read_ready) begin
					phi_last_block_phi_5 = last_BB_reg;
				end
		end
		else
		end
	// controller for phi_5.phi_s_phi_5
	always @(*) begin
		if ((global_state == 2)) begin 
				if (in_read_ready) begin
					phi_s_phi_5 = {32'd0, 32'd2};
				end
		end
		else
		end
	// controller for add_add_7.add_in0_add_7
	always @(*) begin
		if ((global_state == 2)) begin 
				if (in_read_ready) begin
					add_in0_add_7 = phi_out_phi_5;
				end
		end
		else
		end
	// controller for add_add_7.add_in1_add_7
	always @(*) begin
		if ((global_state == 2)) begin 
				if (in_read_ready) begin
					add_in1_add_7 = (32'd1);
				end
		end
		else
		end
	// controller for icmp_8.cmp_in0_icmp_8
	always @(*) begin
		if ((global_state == 2)) begin 
				if (in_read_ready) begin
					cmp_in0_icmp_8 = add_out_add_7;
				end
		end
		else
		end
	// controller for icmp_8.cmp_in1_icmp_8
	always @(*) begin
		if ((global_state == 2)) begin 
				if (in_read_ready) begin
					cmp_in1_icmp_8 = (32'd4);
				end
		end
		else
		end
	// controller for in.in_read_valid_reg
	always @(*) begin
		if ((global_state == 3)) begin 
				if (1) begin
					in_read_valid_reg = -(1'd1);
				end
		end
		if ((global_state == 4)) begin 
				if (1) begin
					in_read_valid_reg = (1'd0);
				end
		end
		else
			in_read_valid_reg = 0;
		end
	// controller for add_add_12.add_in0_add_12
	always @(*) begin
		if ((global_state == 4)) begin 
				if (1) begin
					add_in0_add_12 = load_tmp_1;
				end
		end
		else
		end
	// controller for add_add_12.add_in1_add_12
	always @(*) begin
		if ((global_state == 4)) begin 
				if (1) begin
					add_in1_add_12 = in_out_data;
				end
		end
		else
		end
	// controller for out.out_in_data_reg
	always @(*) begin
		if ((global_state == 7)) begin 
				if (1) begin
					out_in_data_reg = rdata_ram_0;
				end
		end
		else
			out_in_data_reg = 0;
		end
	// controller for out.out_write_valid_reg
	always @(*) begin
		if ((global_state == 7)) begin 
				if (1) begin
					out_write_valid_reg = -(1'd1);
				end
		end
		if ((global_state == 8)) begin 
				if (1) begin
					out_write_valid_reg = (1'd0);
				end
		end
		else
			out_write_valid_reg = 0;
		end
	// controller for ret_24.valid_reg
	always @(*) begin
		if ((global_state == 8)) begin 
				if (1) begin
					valid_reg = 1;
				end
		end
		else
			valid_reg = 0;
		end
endmodule

module channel_reduce_4(input [0:0] clk, input [0:0] rst, output [31:0] out_in_data, output [0:0] out_read_valid, output [0:0] out_rst, output [31:0] out_write_valid, input [31:0] out_out_data, input [0:0] out_read_ready, input [0:0] out_write_ready, output [0:0] valid, output [31:0] in_in_data, output [0:0] in_read_valid, output [0:0] in_rst, output [31:0] in_write_valid, input [31:0] in_out_data, input [0:0] in_read_ready, input [0:0] in_write_ready);


	initial begin
	end




	channel_reduce_4_inner inner(.clk(clk), .in_in_data(in_in_data), .in_out_data(in_out_data), .in_read_ready(in_read_ready), .in_read_valid(in_read_valid), .in_rst(in_rst), .in_write_ready(in_write_ready), .in_write_valid(in_write_valid), .out_in_data(out_in_data), .out_out_data(out_out_data), .out_read_ready(out_read_ready), .out_read_valid(out_read_valid), .out_rst(out_rst), .out_write_ready(out_write_ready), .out_write_valid(out_write_valid), .rst(rst), .valid(valid));

endmodule
