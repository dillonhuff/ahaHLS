module channel_reduce_4(input [0:0] clk, input [0:0] rst, output [31:0] in_in_data, output [0:0] in_read_valid, output [0:0] in_rst, output [0:0] in_write_valid, input [31:0] in_out_data, input [0:0] in_read_ready, input [0:0] in_write_ready, output [0:0] valid, output [31:0] out_in_data, output [0:0] out_read_valid, output [0:0] out_rst, output [0:0] out_write_valid, input [31:0] out_out_data, input [0:0] out_read_ready, input [0:0] out_write_ready);

	reg [31:0] in_in_data_reg;
	reg [0:0] in_read_valid_reg;
	reg [0:0] in_rst_reg;
	reg [0:0] in_write_valid_reg;
	reg [0:0] valid_reg;
	reg [31:0] out_in_data_reg;
	reg [0:0] out_read_valid_reg;
	reg [0:0] out_rst_reg;
	reg [0:0] out_write_valid_reg;

	assign in_in_data = in_in_data_reg;
	assign in_read_valid = in_read_valid_reg;
	assign in_rst = in_rst_reg;
	assign in_write_valid = in_write_valid_reg;
	assign valid = valid_reg;
	assign out_in_data = out_in_data_reg;
	assign out_read_valid = out_read_valid_reg;
	assign out_rst = out_rst_reg;
	assign out_write_valid = out_write_valid_reg;

	// Start debug wires and ports

	initial begin
	end





	// End debug wires and ports

	// Start Functional Units
	br_dummy br_unit();

	add alloca_0();

	add bitcast_1();

	add call_2();

	reg [31:0] raddr_ram_0_reg;
	reg [31:0] waddr_ram_0_reg;
	reg [31:0] wdata_ram_0_reg;
	reg [0:0] wen_ram_0_reg;
	wire [31:0] rdata_ram_0;
	register #(.WIDTH(32)) ram_0(.clk(clk), .raddr(raddr_ram_0_reg), .rdata(rdata_ram_0), .rst(rst), .waddr(waddr_ram_0_reg), .wdata(wdata_ram_0_reg), .wen(wen_ram_0_reg));

	add call_20();

	reg [63:0] phi_in_phi_7;
	reg [31:0] phi_last_block_phi_7;
	reg [63:0] phi_s_phi_7;
	wire [31:0] phi_out_phi_7;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_7(.in(phi_in_phi_7), .last_block(phi_last_block_phi_7), .out(phi_out_phi_7), .s(phi_s_phi_7));

	reg [31:0] add_in0_add_13;
	reg [31:0] add_in1_add_13;
	wire [31:0] add_out_add_13;
	add #(.WIDTH(32)) add_add_13(.in0(add_in0_add_13), .in1(add_in1_add_13), .out(add_out_add_13));

	reg [31:0] add_in0_add_15;
	reg [31:0] add_in1_add_15;
	wire [31:0] add_out_add_15;
	add #(.WIDTH(32)) add_add_15(.in0(add_in0_add_15), .in1(add_in1_add_15), .out(add_out_add_15));

	reg [31:0] cmp_in0_icmp_16;
	reg [31:0] cmp_in1_icmp_16;
	wire [0:0] cmp_out_icmp_16;
	eq #(.WIDTH(32)) icmp_16(.in0(cmp_in0_icmp_16), .in1(cmp_in1_icmp_16), .out(cmp_out_icmp_16));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] bb_8_active_in_state_1_in_data;
	wire [0:0] bb_8_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active_in_state_1(.in_data(bb_8_active_in_state_1_in_data), .out_data(bb_8_active_in_state_1_out_data));

	reg [31:0] bb_8_predecessor_in_state_1_in_data;
	wire [31:0] bb_8_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor_in_state_1(.in_data(bb_8_predecessor_in_state_1_in_data), .out_data(bb_8_predecessor_in_state_1_out_data));

	reg [0:0] bb_0_active_in_state_1_in_data;
	wire [0:0] bb_0_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_1(.in_data(bb_0_active_in_state_1_in_data), .out_data(bb_0_active_in_state_1_out_data));

	reg [31:0] bb_0_predecessor_in_state_1_in_data;
	wire [31:0] bb_0_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_1(.in_data(bb_0_predecessor_in_state_1_in_data), .out_data(bb_0_predecessor_in_state_1_out_data));

	reg [0:0] bb_3_active_in_state_1_in_data;
	wire [0:0] bb_3_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_1(.in_data(bb_3_active_in_state_1_in_data), .out_data(bb_3_active_in_state_1_out_data));

	reg [31:0] bb_3_predecessor_in_state_1_in_data;
	wire [31:0] bb_3_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_1(.in_data(bb_3_predecessor_in_state_1_in_data), .out_data(bb_3_predecessor_in_state_1_out_data));

	reg [0:0] bb_9_active_in_state_1_in_data;
	wire [0:0] bb_9_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_9_active_in_state_1(.in_data(bb_9_active_in_state_1_in_data), .out_data(bb_9_active_in_state_1_out_data));

	reg [31:0] bb_9_predecessor_in_state_1_in_data;
	wire [31:0] bb_9_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_9_predecessor_in_state_1(.in_data(bb_9_predecessor_in_state_1_in_data), .out_data(bb_9_predecessor_in_state_1_out_data));

	reg [0:0] bb_10_active_in_state_2_in_data;
	wire [0:0] bb_10_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_2(.in_data(bb_10_active_in_state_2_in_data), .out_data(bb_10_active_in_state_2_out_data));

	reg [31:0] bb_10_predecessor_in_state_2_in_data;
	wire [31:0] bb_10_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_2(.in_data(bb_10_predecessor_in_state_2_in_data), .out_data(bb_10_predecessor_in_state_2_out_data));

	reg [0:0] bb_4_active_in_state_3_in_data;
	wire [0:0] bb_4_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_3(.in_data(bb_4_active_in_state_3_in_data), .out_data(bb_4_active_in_state_3_out_data));

	reg [31:0] bb_4_predecessor_in_state_3_in_data;
	wire [31:0] bb_4_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_3(.in_data(bb_4_predecessor_in_state_3_in_data), .out_data(bb_4_predecessor_in_state_3_out_data));

	reg [0:0] bb_10_active_in_state_3_in_data;
	wire [0:0] bb_10_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_3(.in_data(bb_10_active_in_state_3_in_data), .out_data(bb_10_active_in_state_3_out_data));

	reg [31:0] bb_10_predecessor_in_state_3_in_data;
	wire [31:0] bb_10_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_3(.in_data(bb_10_predecessor_in_state_3_in_data), .out_data(bb_10_predecessor_in_state_3_out_data));

	reg [0:0] bb_5_active_in_state_4_in_data;
	wire [0:0] bb_5_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_5_active_in_state_4(.in_data(bb_5_active_in_state_4_in_data), .out_data(bb_5_active_in_state_4_out_data));

	reg [31:0] bb_5_predecessor_in_state_4_in_data;
	wire [31:0] bb_5_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_5_predecessor_in_state_4(.in_data(bb_5_predecessor_in_state_4_in_data), .out_data(bb_5_predecessor_in_state_4_out_data));

	reg [0:0] bb_6_active_in_state_4_in_data;
	wire [0:0] bb_6_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_6_active_in_state_4(.in_data(bb_6_active_in_state_4_in_data), .out_data(bb_6_active_in_state_4_out_data));

	reg [31:0] bb_6_predecessor_in_state_4_in_data;
	wire [31:0] bb_6_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_6_predecessor_in_state_4(.in_data(bb_6_predecessor_in_state_4_in_data), .out_data(bb_6_predecessor_in_state_4_out_data));

	reg [0:0] bb_7_active_in_state_4_in_data;
	wire [0:0] bb_7_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_7_active_in_state_4(.in_data(bb_7_active_in_state_4_in_data), .out_data(bb_7_active_in_state_4_out_data));

	reg [31:0] bb_7_predecessor_in_state_4_in_data;
	wire [31:0] bb_7_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_7_predecessor_in_state_4(.in_data(bb_7_predecessor_in_state_4_in_data), .out_data(bb_7_predecessor_in_state_4_out_data));

	reg [0:0] bb_4_active_in_state_4_in_data;
	wire [0:0] bb_4_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_4(.in_data(bb_4_active_in_state_4_in_data), .out_data(bb_4_active_in_state_4_out_data));

	reg [31:0] bb_4_predecessor_in_state_4_in_data;
	wire [31:0] bb_4_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_4(.in_data(bb_4_predecessor_in_state_4_in_data), .out_data(bb_4_predecessor_in_state_4_out_data));

	reg [0:0] bb_2_active_in_state_4_in_data;
	wire [0:0] bb_2_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_4(.in_data(bb_2_active_in_state_4_in_data), .out_data(bb_2_active_in_state_4_out_data));

	reg [31:0] bb_2_predecessor_in_state_4_in_data;
	wire [31:0] bb_2_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_4(.in_data(bb_2_predecessor_in_state_4_in_data), .out_data(bb_2_predecessor_in_state_4_out_data));

	reg [0:0] bb_1_active_in_state_4_in_data;
	wire [0:0] bb_1_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_4(.in_data(bb_1_active_in_state_4_in_data), .out_data(bb_1_active_in_state_4_out_data));

	reg [31:0] bb_1_predecessor_in_state_4_in_data;
	wire [31:0] bb_1_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_4(.in_data(bb_1_predecessor_in_state_4_in_data), .out_data(bb_1_predecessor_in_state_4_out_data));

	reg [0:0] andOp_45_in0;
	reg [0:0] andOp_45_in1;
	wire [0:0] andOp_45_out;
	andOp #(.WIDTH(1)) andOp_45(.in0(andOp_45_in0), .in1(andOp_45_in1), .out(andOp_45_out));

	reg [0:0] andOp_46_in0;
	reg [0:0] andOp_46_in1;
	wire [0:0] andOp_46_out;
	andOp #(.WIDTH(1)) andOp_46(.in0(andOp_46_in0), .in1(andOp_46_in1), .out(andOp_46_out));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] notOp_47_in0;
	wire [0:0] notOp_47_out;
	notOp #(.WIDTH(1)) notOp_47(.in(notOp_47_in0), .out(notOp_47_out));

	reg [0:0] andOp_48_in0;
	reg [0:0] andOp_48_in1;
	wire [0:0] andOp_48_out;
	andOp #(.WIDTH(1)) andOp_48(.in0(andOp_48_in0), .in1(andOp_48_in1), .out(andOp_48_out));

	reg [0:0] andOp_49_in0;
	reg [0:0] andOp_49_in1;
	wire [0:0] andOp_49_out;
	andOp #(.WIDTH(1)) andOp_49(.in0(andOp_49_in0), .in1(andOp_49_in1), .out(andOp_49_out));

	reg [0:0] br_8_happened_in_state_1_in_data;
	wire [0:0] br_8_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_8_happened_in_state_1(.in_data(br_8_happened_in_state_1_in_data), .out_data(br_8_happened_in_state_1_out_data));

	reg [0:0] notOp_50_in0;
	wire [0:0] notOp_50_out;
	notOp #(.WIDTH(1)) notOp_50(.in(notOp_50_in0), .out(notOp_50_out));

	reg [0:0] andOp_51_in0;
	reg [0:0] andOp_51_in1;
	wire [0:0] andOp_51_out;
	andOp #(.WIDTH(1)) andOp_51(.in0(andOp_51_in0), .in1(andOp_51_in1), .out(andOp_51_out));

	reg [0:0] andOp_52_in0;
	reg [0:0] andOp_52_in1;
	wire [0:0] andOp_52_out;
	andOp #(.WIDTH(1)) andOp_52(.in0(andOp_52_in0), .in1(andOp_52_in1), .out(andOp_52_out));

	reg [0:0] br_0_happened_in_state_1_in_data;
	wire [0:0] br_0_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_1(.in_data(br_0_happened_in_state_1_in_data), .out_data(br_0_happened_in_state_1_out_data));

	reg [0:0] notOp_53_in0;
	wire [0:0] notOp_53_out;
	notOp #(.WIDTH(1)) notOp_53(.in(notOp_53_in0), .out(notOp_53_out));

	reg [0:0] andOp_54_in0;
	reg [0:0] andOp_54_in1;
	wire [0:0] andOp_54_out;
	andOp #(.WIDTH(1)) andOp_54(.in0(andOp_54_in0), .in1(andOp_54_in1), .out(andOp_54_out));

	reg [0:0] andOp_55_in0;
	reg [0:0] andOp_55_in1;
	wire [0:0] andOp_55_out;
	andOp #(.WIDTH(1)) andOp_55(.in0(andOp_55_in0), .in1(andOp_55_in1), .out(andOp_55_out));

	reg [0:0] br_3_happened_in_state_1_in_data;
	wire [0:0] br_3_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_1(.in_data(br_3_happened_in_state_1_in_data), .out_data(br_3_happened_in_state_1_out_data));

	reg [0:0] notOp_56_in0;
	wire [0:0] notOp_56_out;
	notOp #(.WIDTH(1)) notOp_56(.in(notOp_56_in0), .out(notOp_56_out));

	reg [0:0] andOp_57_in0;
	reg [0:0] andOp_57_in1;
	wire [0:0] andOp_57_out;
	andOp #(.WIDTH(1)) andOp_57(.in0(andOp_57_in0), .in1(andOp_57_in1), .out(andOp_57_out));

	reg [0:0] andOp_58_in0;
	reg [0:0] andOp_58_in1;
	wire [0:0] andOp_58_out;
	andOp #(.WIDTH(1)) andOp_58(.in0(andOp_58_in0), .in1(andOp_58_in1), .out(andOp_58_out));

	reg [0:0] br_9_happened_in_state_1_in_data;
	wire [0:0] br_9_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_9_happened_in_state_1(.in_data(br_9_happened_in_state_1_in_data), .out_data(br_9_happened_in_state_1_out_data));

	reg [0:0] notOp_59_in0;
	wire [0:0] notOp_59_out;
	notOp #(.WIDTH(1)) notOp_59(.in(notOp_59_in0), .out(notOp_59_out));

	reg [0:0] andOp_60_in0;
	reg [0:0] andOp_60_in1;
	wire [0:0] andOp_60_out;
	andOp #(.WIDTH(1)) andOp_60(.in0(andOp_60_in0), .in1(andOp_60_in1), .out(andOp_60_out));

	reg [0:0] notOp_61_in0;
	wire [0:0] notOp_61_out;
	notOp #(.WIDTH(1)) notOp_61(.in(notOp_61_in0), .out(notOp_61_out));

	reg [0:0] andOp_62_in0;
	reg [0:0] andOp_62_in1;
	wire [0:0] andOp_62_out;
	andOp #(.WIDTH(1)) andOp_62(.in0(andOp_62_in0), .in1(andOp_62_in1), .out(andOp_62_out));

	reg [0:0] andOp_63_in0;
	reg [0:0] andOp_63_in1;
	wire [0:0] andOp_63_out;
	andOp #(.WIDTH(1)) andOp_63(.in0(andOp_63_in0), .in1(andOp_63_in1), .out(andOp_63_out));

	reg [0:0] andOp_64_in0;
	reg [0:0] andOp_64_in1;
	wire [0:0] andOp_64_out;
	andOp #(.WIDTH(1)) andOp_64(.in0(andOp_64_in0), .in1(andOp_64_in1), .out(andOp_64_out));

	reg [0:0] br_10_happened_in_state_2_in_data;
	wire [0:0] br_10_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_2(.in_data(br_10_happened_in_state_2_in_data), .out_data(br_10_happened_in_state_2_out_data));

	reg [0:0] notOp_65_in0;
	wire [0:0] notOp_65_out;
	notOp #(.WIDTH(1)) notOp_65(.in(notOp_65_in0), .out(notOp_65_out));

	reg [0:0] andOp_66_in0;
	reg [0:0] andOp_66_in1;
	wire [0:0] andOp_66_out;
	andOp #(.WIDTH(1)) andOp_66(.in0(andOp_66_in0), .in1(andOp_66_in1), .out(andOp_66_out));

	reg [0:0] andOp_67_in0;
	reg [0:0] andOp_67_in1;
	wire [0:0] andOp_67_out;
	andOp #(.WIDTH(1)) andOp_67(.in0(andOp_67_in0), .in1(andOp_67_in1), .out(andOp_67_out));

	reg [0:0] br_4_happened_in_state_3_in_data;
	wire [0:0] br_4_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_3(.in_data(br_4_happened_in_state_3_in_data), .out_data(br_4_happened_in_state_3_out_data));

	reg [0:0] notOp_68_in0;
	wire [0:0] notOp_68_out;
	notOp #(.WIDTH(1)) notOp_68(.in(notOp_68_in0), .out(notOp_68_out));

	reg [0:0] andOp_69_in0;
	reg [0:0] andOp_69_in1;
	wire [0:0] andOp_69_out;
	andOp #(.WIDTH(1)) andOp_69(.in0(andOp_69_in0), .in1(andOp_69_in1), .out(andOp_69_out));

	reg [0:0] notOp_70_in0;
	wire [0:0] notOp_70_out;
	notOp #(.WIDTH(1)) notOp_70(.in(notOp_70_in0), .out(notOp_70_out));

	reg [0:0] andOp_71_in0;
	reg [0:0] andOp_71_in1;
	wire [0:0] andOp_71_out;
	andOp #(.WIDTH(1)) andOp_71(.in0(andOp_71_in0), .in1(andOp_71_in1), .out(andOp_71_out));

	reg [0:0] andOp_72_in0;
	reg [0:0] andOp_72_in1;
	wire [0:0] andOp_72_out;
	andOp #(.WIDTH(1)) andOp_72(.in0(andOp_72_in0), .in1(andOp_72_in1), .out(andOp_72_out));

	reg [0:0] andOp_73_in0;
	reg [0:0] andOp_73_in1;
	wire [0:0] andOp_73_out;
	andOp #(.WIDTH(1)) andOp_73(.in0(andOp_73_in0), .in1(andOp_73_in1), .out(andOp_73_out));

	reg [0:0] br_10_happened_in_state_3_in_data;
	wire [0:0] br_10_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_3(.in_data(br_10_happened_in_state_3_in_data), .out_data(br_10_happened_in_state_3_out_data));

	reg [0:0] notOp_74_in0;
	wire [0:0] notOp_74_out;
	notOp #(.WIDTH(1)) notOp_74(.in(notOp_74_in0), .out(notOp_74_out));

	reg [0:0] andOp_75_in0;
	reg [0:0] andOp_75_in1;
	wire [0:0] andOp_75_out;
	andOp #(.WIDTH(1)) andOp_75(.in0(andOp_75_in0), .in1(andOp_75_in1), .out(andOp_75_out));

	reg [0:0] andOp_76_in0;
	reg [0:0] andOp_76_in1;
	wire [0:0] andOp_76_out;
	andOp #(.WIDTH(1)) andOp_76(.in0(andOp_76_in0), .in1(andOp_76_in1), .out(andOp_76_out));

	reg [0:0] br_5_happened_in_state_4_in_data;
	wire [0:0] br_5_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_5_happened_in_state_4(.in_data(br_5_happened_in_state_4_in_data), .out_data(br_5_happened_in_state_4_out_data));

	reg [0:0] notOp_77_in0;
	wire [0:0] notOp_77_out;
	notOp #(.WIDTH(1)) notOp_77(.in(notOp_77_in0), .out(notOp_77_out));

	reg [0:0] andOp_78_in0;
	reg [0:0] andOp_78_in1;
	wire [0:0] andOp_78_out;
	andOp #(.WIDTH(1)) andOp_78(.in0(andOp_78_in0), .in1(andOp_78_in1), .out(andOp_78_out));

	reg [0:0] andOp_79_in0;
	reg [0:0] andOp_79_in1;
	wire [0:0] andOp_79_out;
	andOp #(.WIDTH(1)) andOp_79(.in0(andOp_79_in0), .in1(andOp_79_in1), .out(andOp_79_out));

	reg [0:0] br_6_happened_in_state_4_in_data;
	wire [0:0] br_6_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_6_happened_in_state_4(.in_data(br_6_happened_in_state_4_in_data), .out_data(br_6_happened_in_state_4_out_data));

	reg [0:0] notOp_80_in0;
	wire [0:0] notOp_80_out;
	notOp #(.WIDTH(1)) notOp_80(.in(notOp_80_in0), .out(notOp_80_out));

	reg [0:0] andOp_81_in0;
	reg [0:0] andOp_81_in1;
	wire [0:0] andOp_81_out;
	andOp #(.WIDTH(1)) andOp_81(.in0(andOp_81_in0), .in1(andOp_81_in1), .out(andOp_81_out));

	reg [0:0] notOp_82_in0;
	wire [0:0] notOp_82_out;
	notOp #(.WIDTH(1)) notOp_82(.in(notOp_82_in0), .out(notOp_82_out));

	reg [0:0] andOp_83_in0;
	reg [0:0] andOp_83_in1;
	wire [0:0] andOp_83_out;
	andOp #(.WIDTH(1)) andOp_83(.in0(andOp_83_in0), .in1(andOp_83_in1), .out(andOp_83_out));

	reg [0:0] andOp_84_in0;
	reg [0:0] andOp_84_in1;
	wire [0:0] andOp_84_out;
	andOp #(.WIDTH(1)) andOp_84(.in0(andOp_84_in0), .in1(andOp_84_in1), .out(andOp_84_out));

	reg [0:0] andOp_85_in0;
	reg [0:0] andOp_85_in1;
	wire [0:0] andOp_85_out;
	andOp #(.WIDTH(1)) andOp_85(.in0(andOp_85_in0), .in1(andOp_85_in1), .out(andOp_85_out));

	reg [0:0] br_7_happened_in_state_4_in_data;
	wire [0:0] br_7_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_7_happened_in_state_4(.in_data(br_7_happened_in_state_4_in_data), .out_data(br_7_happened_in_state_4_out_data));

	reg [0:0] notOp_86_in0;
	wire [0:0] notOp_86_out;
	notOp #(.WIDTH(1)) notOp_86(.in(notOp_86_in0), .out(notOp_86_out));

	reg [0:0] andOp_87_in0;
	reg [0:0] andOp_87_in1;
	wire [0:0] andOp_87_out;
	andOp #(.WIDTH(1)) andOp_87(.in0(andOp_87_in0), .in1(andOp_87_in1), .out(andOp_87_out));

	reg [0:0] andOp_88_in0;
	reg [0:0] andOp_88_in1;
	wire [0:0] andOp_88_out;
	andOp #(.WIDTH(1)) andOp_88(.in0(andOp_88_in0), .in1(andOp_88_in1), .out(andOp_88_out));

	reg [0:0] br_4_happened_in_state_4_in_data;
	wire [0:0] br_4_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_4(.in_data(br_4_happened_in_state_4_in_data), .out_data(br_4_happened_in_state_4_out_data));

	reg [0:0] notOp_89_in0;
	wire [0:0] notOp_89_out;
	notOp #(.WIDTH(1)) notOp_89(.in(notOp_89_in0), .out(notOp_89_out));

	reg [0:0] andOp_90_in0;
	reg [0:0] andOp_90_in1;
	wire [0:0] andOp_90_out;
	andOp #(.WIDTH(1)) andOp_90(.in0(andOp_90_in0), .in1(andOp_90_in1), .out(andOp_90_out));

	reg [0:0] notOp_91_in0;
	wire [0:0] notOp_91_out;
	notOp #(.WIDTH(1)) notOp_91(.in(notOp_91_in0), .out(notOp_91_out));

	reg [0:0] andOp_92_in0;
	reg [0:0] andOp_92_in1;
	wire [0:0] andOp_92_out;
	andOp #(.WIDTH(1)) andOp_92(.in0(andOp_92_in0), .in1(andOp_92_in1), .out(andOp_92_out));

	reg [0:0] andOp_93_in0;
	reg [0:0] andOp_93_in1;
	wire [0:0] andOp_93_out;
	andOp #(.WIDTH(1)) andOp_93(.in0(andOp_93_in0), .in1(andOp_93_in1), .out(andOp_93_out));

	reg [0:0] andOp_94_in0;
	reg [0:0] andOp_94_in1;
	wire [0:0] andOp_94_out;
	andOp #(.WIDTH(1)) andOp_94(.in0(andOp_94_in0), .in1(andOp_94_in1), .out(andOp_94_out));

	reg [0:0] br_1_happened_in_state_4_in_data;
	wire [0:0] br_1_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened_in_state_4(.in_data(br_1_happened_in_state_4_in_data), .out_data(br_1_happened_in_state_4_out_data));

	reg [0:0] notOp_95_in0;
	wire [0:0] notOp_95_out;
	notOp #(.WIDTH(1)) notOp_95(.in(notOp_95_in0), .out(notOp_95_out));

	reg [31:0] eq_96_in0;
	reg [31:0] eq_96_in1;
	wire [0:0] eq_96_out;
	eq #(.WIDTH(32)) eq_96(.in0(eq_96_in0), .in1(eq_96_in1), .out(eq_96_out));

	reg [31:0] eq_97_in0;
	reg [31:0] eq_97_in1;
	wire [0:0] eq_97_out;
	eq #(.WIDTH(32)) eq_97(.in0(eq_97_in0), .in1(eq_97_in1), .out(eq_97_out));

	reg [0:0] orOp_98_in0;
	reg [0:0] orOp_98_in1;
	wire [0:0] orOp_98_out;
	orOp #(.WIDTH(1)) orOp_98(.in0(orOp_98_in0), .in1(orOp_98_in1), .out(orOp_98_out));

	reg [31:0] eq_99_in0;
	reg [31:0] eq_99_in1;
	wire [0:0] eq_99_out;
	eq #(.WIDTH(32)) eq_99(.in0(eq_99_in0), .in1(eq_99_in1), .out(eq_99_out));

	reg [31:0] eq_100_in0;
	reg [31:0] eq_100_in1;
	wire [0:0] eq_100_out;
	eq #(.WIDTH(32)) eq_100(.in0(eq_100_in0), .in1(eq_100_in1), .out(eq_100_out));

	reg [0:0] orOp_101_in0;
	reg [0:0] orOp_101_in1;
	wire [0:0] orOp_101_out;
	orOp #(.WIDTH(1)) orOp_101(.in0(orOp_101_in0), .in1(orOp_101_in1), .out(orOp_101_out));

	reg [31:0] eq_102_in0;
	reg [31:0] eq_102_in1;
	wire [0:0] eq_102_out;
	eq #(.WIDTH(32)) eq_102(.in0(eq_102_in0), .in1(eq_102_in1), .out(eq_102_out));

	reg [0:0] orOp_103_in0;
	reg [0:0] orOp_103_in1;
	wire [0:0] orOp_103_out;
	orOp #(.WIDTH(1)) orOp_103(.in0(orOp_103_in0), .in1(orOp_103_in1), .out(orOp_103_out));

	reg [31:0] eq_104_in0;
	reg [31:0] eq_104_in1;
	wire [0:0] eq_104_out;
	eq #(.WIDTH(32)) eq_104(.in0(eq_104_in0), .in1(eq_104_in1), .out(eq_104_out));

	reg [31:0] eq_105_in0;
	reg [31:0] eq_105_in1;
	wire [0:0] eq_105_out;
	eq #(.WIDTH(32)) eq_105(.in0(eq_105_in0), .in1(eq_105_in1), .out(eq_105_out));

	reg [0:0] orOp_106_in0;
	reg [0:0] orOp_106_in1;
	wire [0:0] orOp_106_out;
	orOp #(.WIDTH(1)) orOp_106(.in0(orOp_106_in0), .in1(orOp_106_in1), .out(orOp_106_out));

	reg [31:0] eq_107_in0;
	reg [31:0] eq_107_in1;
	wire [0:0] eq_107_out;
	eq #(.WIDTH(32)) eq_107(.in0(eq_107_in0), .in1(eq_107_in1), .out(eq_107_out));

	reg [31:0] eq_108_in0;
	reg [31:0] eq_108_in1;
	wire [0:0] eq_108_out;
	eq #(.WIDTH(32)) eq_108(.in0(eq_108_in0), .in1(eq_108_in1), .out(eq_108_out));

	reg [0:0] orOp_109_in0;
	reg [0:0] orOp_109_in1;
	wire [0:0] orOp_109_out;
	orOp #(.WIDTH(1)) orOp_109(.in0(orOp_109_in0), .in1(orOp_109_in1), .out(orOp_109_out));

	reg [31:0] eq_110_in0;
	reg [31:0] eq_110_in1;
	wire [0:0] eq_110_out;
	eq #(.WIDTH(32)) eq_110(.in0(eq_110_in0), .in1(eq_110_in1), .out(eq_110_out));

	reg [0:0] orOp_111_in0;
	reg [0:0] orOp_111_in1;
	wire [0:0] orOp_111_out;
	orOp #(.WIDTH(1)) orOp_111(.in0(orOp_111_in0), .in1(orOp_111_in1), .out(orOp_111_out));

	reg [31:0] eq_112_in0;
	reg [31:0] eq_112_in1;
	wire [0:0] eq_112_out;
	eq #(.WIDTH(32)) eq_112(.in0(eq_112_in0), .in1(eq_112_in1), .out(eq_112_out));

	reg [0:0] orOp_113_in0;
	reg [0:0] orOp_113_in1;
	wire [0:0] orOp_113_out;
	orOp #(.WIDTH(1)) orOp_113(.in0(orOp_113_in0), .in1(orOp_113_in1), .out(orOp_113_out));

	reg [31:0] eq_114_in0;
	reg [31:0] eq_114_in1;
	wire [0:0] eq_114_out;
	eq #(.WIDTH(32)) eq_114(.in0(eq_114_in0), .in1(eq_114_in1), .out(eq_114_out));

	reg [31:0] eq_115_in0;
	reg [31:0] eq_115_in1;
	wire [0:0] eq_115_out;
	eq #(.WIDTH(32)) eq_115(.in0(eq_115_in0), .in1(eq_115_in1), .out(eq_115_out));

	reg [0:0] orOp_116_in0;
	reg [0:0] orOp_116_in1;
	wire [0:0] orOp_116_out;
	orOp #(.WIDTH(1)) orOp_116(.in0(orOp_116_in0), .in1(orOp_116_in1), .out(orOp_116_out));

	reg [31:0] eq_117_in0;
	reg [31:0] eq_117_in1;
	wire [0:0] eq_117_out;
	eq #(.WIDTH(32)) eq_117(.in0(eq_117_in0), .in1(eq_117_in1), .out(eq_117_out));

	reg [0:0] orOp_118_in0;
	reg [0:0] orOp_118_in1;
	wire [0:0] orOp_118_out;
	orOp #(.WIDTH(1)) orOp_118(.in0(orOp_118_in0), .in1(orOp_118_in1), .out(orOp_118_out));

	reg [31:0] eq_119_in0;
	reg [31:0] eq_119_in1;
	wire [0:0] eq_119_out;
	eq #(.WIDTH(32)) eq_119(.in0(eq_119_in0), .in1(eq_119_in1), .out(eq_119_out));

	reg [31:0] eq_120_in0;
	reg [31:0] eq_120_in1;
	wire [0:0] eq_120_out;
	eq #(.WIDTH(32)) eq_120(.in0(eq_120_in0), .in1(eq_120_in1), .out(eq_120_out));

	reg [0:0] notOp_121_in0;
	wire [0:0] notOp_121_out;
	notOp #(.WIDTH(1)) notOp_121(.in(notOp_121_in0), .out(notOp_121_out));

	reg [0:0] andOp_122_in0;
	reg [0:0] andOp_122_in1;
	wire [0:0] andOp_122_out;
	andOp #(.WIDTH(1)) andOp_122(.in0(andOp_122_in0), .in1(andOp_122_in1), .out(andOp_122_out));

	reg [31:0] eq_123_in0;
	reg [31:0] eq_123_in1;
	wire [0:0] eq_123_out;
	eq #(.WIDTH(32)) eq_123(.in0(eq_123_in0), .in1(eq_123_in1), .out(eq_123_out));

	reg [31:0] eq_124_in0;
	reg [31:0] eq_124_in1;
	wire [0:0] eq_124_out;
	eq #(.WIDTH(32)) eq_124(.in0(eq_124_in0), .in1(eq_124_in1), .out(eq_124_out));

	reg [0:0] notOp_125_in0;
	wire [0:0] notOp_125_out;
	notOp #(.WIDTH(1)) notOp_125(.in(notOp_125_in0), .out(notOp_125_out));

	reg [0:0] andOp_126_in0;
	reg [0:0] andOp_126_in1;
	wire [0:0] andOp_126_out;
	andOp #(.WIDTH(1)) andOp_126(.in0(andOp_126_in0), .in1(andOp_126_in1), .out(andOp_126_out));

	reg [31:0] eq_127_in0;
	reg [31:0] eq_127_in1;
	wire [0:0] eq_127_out;
	eq #(.WIDTH(32)) eq_127(.in0(eq_127_in0), .in1(eq_127_in1), .out(eq_127_out));

	reg [0:0] notOp_128_in0;
	wire [0:0] notOp_128_out;
	notOp #(.WIDTH(1)) notOp_128(.in(notOp_128_in0), .out(notOp_128_out));

	reg [0:0] andOp_129_in0;
	reg [0:0] andOp_129_in1;
	wire [0:0] andOp_129_out;
	andOp #(.WIDTH(1)) andOp_129(.in0(andOp_129_in0), .in1(andOp_129_in1), .out(andOp_129_out));

	reg [31:0] eq_130_in0;
	reg [31:0] eq_130_in1;
	wire [0:0] eq_130_out;
	eq #(.WIDTH(32)) eq_130(.in0(eq_130_in0), .in1(eq_130_in1), .out(eq_130_out));

	reg [31:0] eq_131_in0;
	reg [31:0] eq_131_in1;
	wire [0:0] eq_131_out;
	eq #(.WIDTH(32)) eq_131(.in0(eq_131_in0), .in1(eq_131_in1), .out(eq_131_out));

	reg [0:0] notOp_132_in0;
	wire [0:0] notOp_132_out;
	notOp #(.WIDTH(1)) notOp_132(.in(notOp_132_in0), .out(notOp_132_out));

	reg [0:0] andOp_133_in0;
	reg [0:0] andOp_133_in1;
	wire [0:0] andOp_133_out;
	andOp #(.WIDTH(1)) andOp_133(.in0(andOp_133_in0), .in1(andOp_133_in1), .out(andOp_133_out));

	reg [31:0] eq_134_in0;
	reg [31:0] eq_134_in1;
	wire [0:0] eq_134_out;
	eq #(.WIDTH(32)) eq_134(.in0(eq_134_in0), .in1(eq_134_in1), .out(eq_134_out));

	reg [31:0] eq_135_in0;
	reg [31:0] eq_135_in1;
	wire [0:0] eq_135_out;
	eq #(.WIDTH(32)) eq_135(.in0(eq_135_in0), .in1(eq_135_in1), .out(eq_135_out));

	reg [0:0] notOp_136_in0;
	wire [0:0] notOp_136_out;
	notOp #(.WIDTH(1)) notOp_136(.in(notOp_136_in0), .out(notOp_136_out));

	reg [0:0] andOp_137_in0;
	reg [0:0] andOp_137_in1;
	wire [0:0] andOp_137_out;
	andOp #(.WIDTH(1)) andOp_137(.in0(andOp_137_in0), .in1(andOp_137_in1), .out(andOp_137_out));

	reg [31:0] eq_138_in0;
	reg [31:0] eq_138_in1;
	wire [0:0] eq_138_out;
	eq #(.WIDTH(32)) eq_138(.in0(eq_138_in0), .in1(eq_138_in1), .out(eq_138_out));

	reg [0:0] notOp_139_in0;
	wire [0:0] notOp_139_out;
	notOp #(.WIDTH(1)) notOp_139(.in(notOp_139_in0), .out(notOp_139_out));

	reg [0:0] andOp_140_in0;
	reg [0:0] andOp_140_in1;
	wire [0:0] andOp_140_out;
	andOp #(.WIDTH(1)) andOp_140(.in0(andOp_140_in0), .in1(andOp_140_in1), .out(andOp_140_out));

	reg [31:0] eq_141_in0;
	reg [31:0] eq_141_in1;
	wire [0:0] eq_141_out;
	eq #(.WIDTH(32)) eq_141(.in0(eq_141_in0), .in1(eq_141_in1), .out(eq_141_out));

	reg [0:0] notOp_142_in0;
	wire [0:0] notOp_142_out;
	notOp #(.WIDTH(1)) notOp_142(.in(notOp_142_in0), .out(notOp_142_out));

	reg [0:0] andOp_143_in0;
	reg [0:0] andOp_143_in1;
	wire [0:0] andOp_143_out;
	andOp #(.WIDTH(1)) andOp_143(.in0(andOp_143_in0), .in1(andOp_143_in1), .out(andOp_143_out));

	reg [31:0] eq_144_in0;
	reg [31:0] eq_144_in1;
	wire [0:0] eq_144_out;
	eq #(.WIDTH(32)) eq_144(.in0(eq_144_in0), .in1(eq_144_in1), .out(eq_144_out));

	reg [31:0] eq_145_in0;
	reg [31:0] eq_145_in1;
	wire [0:0] eq_145_out;
	eq #(.WIDTH(32)) eq_145(.in0(eq_145_in0), .in1(eq_145_in1), .out(eq_145_out));

	reg [0:0] notOp_146_in0;
	wire [0:0] notOp_146_out;
	notOp #(.WIDTH(1)) notOp_146(.in(notOp_146_in0), .out(notOp_146_out));

	reg [0:0] andOp_147_in0;
	reg [0:0] andOp_147_in1;
	wire [0:0] andOp_147_out;
	andOp #(.WIDTH(1)) andOp_147(.in0(andOp_147_in0), .in1(andOp_147_in1), .out(andOp_147_out));

	reg [31:0] eq_148_in0;
	reg [31:0] eq_148_in1;
	wire [0:0] eq_148_out;
	eq #(.WIDTH(32)) eq_148(.in0(eq_148_in0), .in1(eq_148_in1), .out(eq_148_out));

	reg [0:0] notOp_149_in0;
	wire [0:0] notOp_149_out;
	notOp #(.WIDTH(1)) notOp_149(.in(notOp_149_in0), .out(notOp_149_out));

	reg [0:0] andOp_150_in0;
	reg [0:0] andOp_150_in1;
	wire [0:0] andOp_150_out;
	andOp #(.WIDTH(1)) andOp_150(.in0(andOp_150_in0), .in1(andOp_150_in1), .out(andOp_150_out));

	reg [0:0] andOp_151_in0;
	reg [0:0] andOp_151_in1;
	wire [0:0] andOp_151_out;
	andOp #(.WIDTH(1)) andOp_151(.in0(andOp_151_in0), .in1(andOp_151_in1), .out(andOp_151_out));

	reg [0:0] andOp_152_in0;
	reg [0:0] andOp_152_in1;
	wire [0:0] andOp_152_out;
	andOp #(.WIDTH(1)) andOp_152(.in0(andOp_152_in0), .in1(andOp_152_in1), .out(andOp_152_out));

	reg [0:0] andOp_153_in0;
	reg [0:0] andOp_153_in1;
	wire [0:0] andOp_153_out;
	andOp #(.WIDTH(1)) andOp_153(.in0(andOp_153_in0), .in1(andOp_153_in1), .out(andOp_153_out));

	reg [0:0] andOp_154_in0;
	reg [0:0] andOp_154_in1;
	wire [0:0] andOp_154_out;
	andOp #(.WIDTH(1)) andOp_154(.in0(andOp_154_in0), .in1(andOp_154_in1), .out(andOp_154_out));

	reg [0:0] andOp_155_in0;
	reg [0:0] andOp_155_in1;
	wire [0:0] andOp_155_out;
	andOp #(.WIDTH(1)) andOp_155(.in0(andOp_155_in0), .in1(andOp_155_in1), .out(andOp_155_out));

	reg [0:0] andOp_156_in0;
	reg [0:0] andOp_156_in1;
	wire [0:0] andOp_156_out;
	andOp #(.WIDTH(1)) andOp_156(.in0(andOp_156_in0), .in1(andOp_156_in1), .out(andOp_156_out));

	reg [0:0] andOp_157_in0;
	reg [0:0] andOp_157_in1;
	wire [0:0] andOp_157_out;
	andOp #(.WIDTH(1)) andOp_157(.in0(andOp_157_in0), .in1(andOp_157_in1), .out(andOp_157_out));

	reg [0:0] andOp_158_in0;
	reg [0:0] andOp_158_in1;
	wire [0:0] andOp_158_out;
	andOp #(.WIDTH(1)) andOp_158(.in0(andOp_158_in0), .in1(andOp_158_in1), .out(andOp_158_out));

	reg [0:0] andOp_159_in0;
	reg [0:0] andOp_159_in1;
	wire [0:0] andOp_159_out;
	andOp #(.WIDTH(1)) andOp_159(.in0(andOp_159_in0), .in1(andOp_159_in1), .out(andOp_159_out));

	reg [0:0] andOp_160_in0;
	reg [0:0] andOp_160_in1;
	wire [0:0] andOp_160_out;
	andOp #(.WIDTH(1)) andOp_160(.in0(andOp_160_in0), .in1(andOp_160_in1), .out(andOp_160_out));

	reg [0:0] andOp_161_in0;
	reg [0:0] andOp_161_in1;
	wire [0:0] andOp_161_out;
	andOp #(.WIDTH(1)) andOp_161(.in0(andOp_161_in0), .in1(andOp_161_in1), .out(andOp_161_out));

	reg [31:0] concat_162_in0;
	reg [31:0] concat_162_in1;
	wire [63:0] concat_162_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_162(.in0(concat_162_in0), .in1(concat_162_in1), .out(concat_162_out));

	reg [31:0] concat_163_in0;
	reg [31:0] concat_163_in1;
	wire [63:0] concat_163_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_163(.in0(concat_163_in0), .in1(concat_163_in1), .out(concat_163_out));

	reg [0:0] andOp_164_in0;
	reg [0:0] andOp_164_in1;
	wire [0:0] andOp_164_out;
	andOp #(.WIDTH(1)) andOp_164(.in0(andOp_164_in0), .in1(andOp_164_in1), .out(andOp_164_out));

	reg [31:0] tmp_output_165_in_data;
	wire [31:0] tmp_output_165_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_165(.in_data(tmp_output_165_in_data), .out_data(tmp_output_165_out_data));

	reg [31:0] eq_166_in0;
	reg [31:0] eq_166_in1;
	wire [0:0] eq_166_out;
	eq #(.WIDTH(32)) eq_166(.in0(eq_166_in0), .in1(eq_166_in1), .out(eq_166_out));

	reg [0:0] andOp_167_in0;
	reg [0:0] andOp_167_in1;
	wire [0:0] andOp_167_out;
	andOp #(.WIDTH(1)) andOp_167(.in0(andOp_167_in0), .in1(andOp_167_in1), .out(andOp_167_out));

	reg [0:0] andOp_168_in0;
	reg [0:0] andOp_168_in1;
	wire [0:0] andOp_168_out;
	andOp #(.WIDTH(1)) andOp_168(.in0(andOp_168_in0), .in1(andOp_168_in1), .out(andOp_168_out));

	reg [0:0] andOp_169_in0;
	reg [0:0] andOp_169_in1;
	wire [0:0] andOp_169_out;
	andOp #(.WIDTH(1)) andOp_169(.in0(andOp_169_in0), .in1(andOp_169_in1), .out(andOp_169_out));

	reg [0:0] andOp_170_in0;
	reg [0:0] andOp_170_in1;
	wire [0:0] andOp_170_out;
	andOp #(.WIDTH(1)) andOp_170(.in0(andOp_170_in0), .in1(andOp_170_in1), .out(andOp_170_out));

	reg [0:0] andOp_171_in0;
	reg [0:0] andOp_171_in1;
	wire [0:0] andOp_171_out;
	andOp #(.WIDTH(1)) andOp_171(.in0(andOp_171_in0), .in1(andOp_171_in1), .out(andOp_171_out));

	reg [0:0] andOp_172_in0;
	reg [0:0] andOp_172_in1;
	wire [0:0] andOp_172_out;
	andOp #(.WIDTH(1)) andOp_172(.in0(andOp_172_in0), .in1(andOp_172_in1), .out(andOp_172_out));

	reg [0:0] andOp_173_in0;
	reg [0:0] andOp_173_in1;
	wire [0:0] andOp_173_out;
	andOp #(.WIDTH(1)) andOp_173(.in0(andOp_173_in0), .in1(andOp_173_in1), .out(andOp_173_out));

	reg [0:0] andOp_174_in0;
	reg [0:0] andOp_174_in1;
	wire [0:0] andOp_174_out;
	andOp #(.WIDTH(1)) andOp_174(.in0(andOp_174_in0), .in1(andOp_174_in1), .out(andOp_174_out));

	reg [0:0] andOp_175_in0;
	reg [0:0] andOp_175_in1;
	wire [0:0] andOp_175_out;
	andOp #(.WIDTH(1)) andOp_175(.in0(andOp_175_in0), .in1(andOp_175_in1), .out(andOp_175_out));

	reg [0:0] andOp_176_in0;
	reg [0:0] andOp_176_in1;
	wire [0:0] andOp_176_out;
	andOp #(.WIDTH(1)) andOp_176(.in0(andOp_176_in0), .in1(andOp_176_in1), .out(andOp_176_out));

	reg [0:0] andOp_177_in0;
	reg [0:0] andOp_177_in1;
	wire [0:0] andOp_177_out;
	andOp #(.WIDTH(1)) andOp_177(.in0(andOp_177_in0), .in1(andOp_177_in1), .out(andOp_177_out));

	reg [0:0] notOp_178_in0;
	wire [0:0] notOp_178_out;
	notOp #(.WIDTH(1)) notOp_178(.in(notOp_178_in0), .out(notOp_178_out));

	reg [0:0] andOp_179_in0;
	reg [0:0] andOp_179_in1;
	wire [0:0] andOp_179_out;
	andOp #(.WIDTH(1)) andOp_179(.in0(andOp_179_in0), .in1(andOp_179_in1), .out(andOp_179_out));

	reg [0:0] notOp_180_in0;
	wire [0:0] notOp_180_out;
	notOp #(.WIDTH(1)) notOp_180(.in(notOp_180_in0), .out(notOp_180_out));

	reg [0:0] andOp_181_in0;
	reg [0:0] andOp_181_in1;
	wire [0:0] andOp_181_out;
	andOp #(.WIDTH(1)) andOp_181(.in0(andOp_181_in0), .in1(andOp_181_in1), .out(andOp_181_out));

	reg [0:0] notOp_182_in0;
	wire [0:0] notOp_182_out;
	notOp #(.WIDTH(1)) notOp_182(.in(notOp_182_in0), .out(notOp_182_out));

	reg [0:0] andOp_183_in0;
	reg [0:0] andOp_183_in1;
	wire [0:0] andOp_183_out;
	andOp #(.WIDTH(1)) andOp_183(.in0(andOp_183_in0), .in1(andOp_183_in1), .out(andOp_183_out));

	reg [0:0] notOp_184_in0;
	wire [0:0] notOp_184_out;
	notOp #(.WIDTH(1)) notOp_184(.in(notOp_184_in0), .out(notOp_184_out));

	reg [0:0] andOp_185_in0;
	reg [0:0] andOp_185_in1;
	wire [0:0] andOp_185_out;
	andOp #(.WIDTH(1)) andOp_185(.in0(andOp_185_in0), .in1(andOp_185_in1), .out(andOp_185_out));

	reg [0:0] notOp_186_in0;
	wire [0:0] notOp_186_out;
	notOp #(.WIDTH(1)) notOp_186(.in(notOp_186_in0), .out(notOp_186_out));

	reg [0:0] andOp_187_in0;
	reg [0:0] andOp_187_in1;
	wire [0:0] andOp_187_out;
	andOp #(.WIDTH(1)) andOp_187(.in0(andOp_187_in0), .in1(andOp_187_in1), .out(andOp_187_out));

	reg [0:0] notOp_188_in0;
	wire [0:0] notOp_188_out;
	notOp #(.WIDTH(1)) notOp_188(.in(notOp_188_in0), .out(notOp_188_out));

	reg [0:0] andOp_189_in0;
	reg [0:0] andOp_189_in1;
	wire [0:0] andOp_189_out;
	andOp #(.WIDTH(1)) andOp_189(.in0(andOp_189_in0), .in1(andOp_189_in1), .out(andOp_189_out));

	reg [0:0] notOp_190_in0;
	wire [0:0] notOp_190_out;
	notOp #(.WIDTH(1)) notOp_190(.in(notOp_190_in0), .out(notOp_190_out));

	reg [0:0] andOp_191_in0;
	reg [0:0] andOp_191_in1;
	wire [0:0] andOp_191_out;
	andOp #(.WIDTH(1)) andOp_191(.in0(andOp_191_in0), .in1(andOp_191_in1), .out(andOp_191_out));

	reg [0:0] notOp_192_in0;
	wire [0:0] notOp_192_out;
	notOp #(.WIDTH(1)) notOp_192(.in(notOp_192_in0), .out(notOp_192_out));

	reg [0:0] andOp_193_in0;
	reg [0:0] andOp_193_in1;
	wire [0:0] andOp_193_out;
	andOp #(.WIDTH(1)) andOp_193(.in0(andOp_193_in0), .in1(andOp_193_in1), .out(andOp_193_out));

	reg [0:0] andOp_194_in0;
	reg [0:0] andOp_194_in1;
	wire [0:0] andOp_194_out;
	andOp #(.WIDTH(1)) andOp_194(.in0(andOp_194_in0), .in1(andOp_194_in1), .out(andOp_194_out));

	reg [0:0] andOp_195_in0;
	reg [0:0] andOp_195_in1;
	wire [0:0] andOp_195_out;
	andOp #(.WIDTH(1)) andOp_195(.in0(andOp_195_in0), .in1(andOp_195_in1), .out(andOp_195_out));

	reg [0:0] andOp_196_in0;
	reg [0:0] andOp_196_in1;
	wire [0:0] andOp_196_out;
	andOp #(.WIDTH(1)) andOp_196(.in0(andOp_196_in0), .in1(andOp_196_in1), .out(andOp_196_out));

	reg [0:0] andOp_197_in0;
	reg [0:0] andOp_197_in1;
	wire [0:0] andOp_197_out;
	andOp #(.WIDTH(1)) andOp_197(.in0(andOp_197_in0), .in1(andOp_197_in1), .out(andOp_197_out));

	reg [0:0] notOp_198_in0;
	wire [0:0] notOp_198_out;
	notOp #(.WIDTH(1)) notOp_198(.in(notOp_198_in0), .out(notOp_198_out));

	reg [0:0] andOp_199_in0;
	reg [0:0] andOp_199_in1;
	wire [0:0] andOp_199_out;
	andOp #(.WIDTH(1)) andOp_199(.in0(andOp_199_in0), .in1(andOp_199_in1), .out(andOp_199_out));

	reg [0:0] andOp_200_in0;
	reg [0:0] andOp_200_in1;
	wire [0:0] andOp_200_out;
	andOp #(.WIDTH(1)) andOp_200(.in0(andOp_200_in0), .in1(andOp_200_in1), .out(andOp_200_out));

	reg [31:0] eq_201_in0;
	reg [31:0] eq_201_in1;
	wire [0:0] eq_201_out;
	eq #(.WIDTH(32)) eq_201(.in0(eq_201_in0), .in1(eq_201_in1), .out(eq_201_out));

	reg [0:0] andOp_202_in0;
	reg [0:0] andOp_202_in1;
	wire [0:0] andOp_202_out;
	andOp #(.WIDTH(1)) andOp_202(.in0(andOp_202_in0), .in1(andOp_202_in1), .out(andOp_202_out));

	reg [0:0] notOp_203_in0;
	wire [0:0] notOp_203_out;
	notOp #(.WIDTH(1)) notOp_203(.in(notOp_203_in0), .out(notOp_203_out));

	reg [0:0] andOp_204_in0;
	reg [0:0] andOp_204_in1;
	wire [0:0] andOp_204_out;
	andOp #(.WIDTH(1)) andOp_204(.in0(andOp_204_in0), .in1(andOp_204_in1), .out(andOp_204_out));

	reg [31:0] eq_205_in0;
	reg [31:0] eq_205_in1;
	wire [0:0] eq_205_out;
	eq #(.WIDTH(32)) eq_205(.in0(eq_205_in0), .in1(eq_205_in1), .out(eq_205_out));

	reg [0:0] andOp_206_in0;
	reg [0:0] andOp_206_in1;
	wire [0:0] andOp_206_out;
	andOp #(.WIDTH(1)) andOp_206(.in0(andOp_206_in0), .in1(andOp_206_in1), .out(andOp_206_out));

	reg [31:0] eq_207_in0;
	reg [31:0] eq_207_in1;
	wire [0:0] eq_207_out;
	eq #(.WIDTH(32)) eq_207(.in0(eq_207_in0), .in1(eq_207_in1), .out(eq_207_out));

	reg [0:0] andOp_208_in0;
	reg [0:0] andOp_208_in1;
	wire [0:0] andOp_208_out;
	andOp #(.WIDTH(1)) andOp_208(.in0(andOp_208_in0), .in1(andOp_208_in1), .out(andOp_208_out));

	reg [0:0] notOp_209_in0;
	wire [0:0] notOp_209_out;
	notOp #(.WIDTH(1)) notOp_209(.in(notOp_209_in0), .out(notOp_209_out));

	reg [0:0] andOp_210_in0;
	reg [0:0] andOp_210_in1;
	wire [0:0] andOp_210_out;
	andOp #(.WIDTH(1)) andOp_210(.in0(andOp_210_in0), .in1(andOp_210_in1), .out(andOp_210_out));

	reg [0:0] andOp_211_in0;
	reg [0:0] andOp_211_in1;
	wire [0:0] andOp_211_out;
	andOp #(.WIDTH(1)) andOp_211(.in0(andOp_211_in0), .in1(andOp_211_in1), .out(andOp_211_out));

	reg [31:0] eq_212_in0;
	reg [31:0] eq_212_in1;
	wire [0:0] eq_212_out;
	eq #(.WIDTH(32)) eq_212(.in0(eq_212_in0), .in1(eq_212_in1), .out(eq_212_out));

	reg [0:0] andOp_213_in0;
	reg [0:0] andOp_213_in1;
	wire [0:0] andOp_213_out;
	andOp #(.WIDTH(1)) andOp_213(.in0(andOp_213_in0), .in1(andOp_213_in1), .out(andOp_213_out));

	reg [0:0] notOp_214_in0;
	wire [0:0] notOp_214_out;
	notOp #(.WIDTH(1)) notOp_214(.in(notOp_214_in0), .out(notOp_214_out));

	reg [0:0] andOp_215_in0;
	reg [0:0] andOp_215_in1;
	wire [0:0] andOp_215_out;
	andOp #(.WIDTH(1)) andOp_215(.in0(andOp_215_in0), .in1(andOp_215_in1), .out(andOp_215_out));

	reg [31:0] eq_216_in0;
	reg [31:0] eq_216_in1;
	wire [0:0] eq_216_out;
	eq #(.WIDTH(32)) eq_216(.in0(eq_216_in0), .in1(eq_216_in1), .out(eq_216_out));

	reg [0:0] andOp_217_in0;
	reg [0:0] andOp_217_in1;
	wire [0:0] andOp_217_out;
	andOp #(.WIDTH(1)) andOp_217(.in0(andOp_217_in0), .in1(andOp_217_in1), .out(andOp_217_out));

	reg [0:0] notOp_218_in0;
	wire [0:0] notOp_218_out;
	notOp #(.WIDTH(1)) notOp_218(.in(notOp_218_in0), .out(notOp_218_out));

	reg [0:0] andOp_219_in0;
	reg [0:0] andOp_219_in1;
	wire [0:0] andOp_219_out;
	andOp #(.WIDTH(1)) andOp_219(.in0(andOp_219_in0), .in1(andOp_219_in1), .out(andOp_219_out));

	reg [0:0] andOp_220_in0;
	reg [0:0] andOp_220_in1;
	wire [0:0] andOp_220_out;
	andOp #(.WIDTH(1)) andOp_220(.in0(andOp_220_in0), .in1(andOp_220_in1), .out(andOp_220_out));

	reg [31:0] eq_221_in0;
	reg [31:0] eq_221_in1;
	wire [0:0] eq_221_out;
	eq #(.WIDTH(32)) eq_221(.in0(eq_221_in0), .in1(eq_221_in1), .out(eq_221_out));

	reg [0:0] andOp_222_in0;
	reg [0:0] andOp_222_in1;
	wire [0:0] andOp_222_out;
	andOp #(.WIDTH(1)) andOp_222(.in0(andOp_222_in0), .in1(andOp_222_in1), .out(andOp_222_out));

	reg [0:0] notOp_223_in0;
	wire [0:0] notOp_223_out;
	notOp #(.WIDTH(1)) notOp_223(.in(notOp_223_in0), .out(notOp_223_out));

	reg [0:0] andOp_224_in0;
	reg [0:0] andOp_224_in1;
	wire [0:0] andOp_224_out;
	andOp #(.WIDTH(1)) andOp_224(.in0(andOp_224_in0), .in1(andOp_224_in1), .out(andOp_224_out));

	reg [31:0] eq_225_in0;
	reg [31:0] eq_225_in1;
	wire [0:0] eq_225_out;
	eq #(.WIDTH(32)) eq_225(.in0(eq_225_in0), .in1(eq_225_in1), .out(eq_225_out));

	reg [0:0] andOp_226_in0;
	reg [0:0] andOp_226_in1;
	wire [0:0] andOp_226_out;
	andOp #(.WIDTH(1)) andOp_226(.in0(andOp_226_in0), .in1(andOp_226_in1), .out(andOp_226_out));

	reg [31:0] eq_227_in0;
	reg [31:0] eq_227_in1;
	wire [0:0] eq_227_out;
	eq #(.WIDTH(32)) eq_227(.in0(eq_227_in0), .in1(eq_227_in1), .out(eq_227_out));

	reg [0:0] andOp_228_in0;
	reg [0:0] andOp_228_in1;
	wire [0:0] andOp_228_out;
	andOp #(.WIDTH(1)) andOp_228(.in0(andOp_228_in0), .in1(andOp_228_in1), .out(andOp_228_out));

	reg [0:0] notOp_229_in0;
	wire [0:0] notOp_229_out;
	notOp #(.WIDTH(1)) notOp_229(.in(notOp_229_in0), .out(notOp_229_out));

	reg [0:0] andOp_230_in0;
	reg [0:0] andOp_230_in1;
	wire [0:0] andOp_230_out;
	andOp #(.WIDTH(1)) andOp_230(.in0(andOp_230_in0), .in1(andOp_230_in1), .out(andOp_230_out));

	reg [0:0] andOp_231_in0;
	reg [0:0] andOp_231_in1;
	wire [0:0] andOp_231_out;
	andOp #(.WIDTH(1)) andOp_231(.in0(andOp_231_in0), .in1(andOp_231_in1), .out(andOp_231_out));

	reg [31:0] eq_232_in0;
	reg [31:0] eq_232_in1;
	wire [0:0] eq_232_out;
	eq #(.WIDTH(32)) eq_232(.in0(eq_232_in0), .in1(eq_232_in1), .out(eq_232_out));

	reg [0:0] andOp_233_in0;
	reg [0:0] andOp_233_in1;
	wire [0:0] andOp_233_out;
	andOp #(.WIDTH(1)) andOp_233(.in0(andOp_233_in0), .in1(andOp_233_in1), .out(andOp_233_out));

	reg [0:0] notOp_234_in0;
	wire [0:0] notOp_234_out;
	notOp #(.WIDTH(1)) notOp_234(.in(notOp_234_in0), .out(notOp_234_out));

	reg [0:0] andOp_235_in0;
	reg [0:0] andOp_235_in1;
	wire [0:0] andOp_235_out;
	andOp #(.WIDTH(1)) andOp_235(.in0(andOp_235_in0), .in1(andOp_235_in1), .out(andOp_235_out));

	reg [31:0] eq_236_in0;
	reg [31:0] eq_236_in1;
	wire [0:0] eq_236_out;
	eq #(.WIDTH(32)) eq_236(.in0(eq_236_in0), .in1(eq_236_in1), .out(eq_236_out));

	reg [0:0] andOp_237_in0;
	reg [0:0] andOp_237_in1;
	wire [0:0] andOp_237_out;
	andOp #(.WIDTH(1)) andOp_237(.in0(andOp_237_in0), .in1(andOp_237_in1), .out(andOp_237_out));

	reg [0:0] notOp_238_in0;
	wire [0:0] notOp_238_out;
	notOp #(.WIDTH(1)) notOp_238(.in(notOp_238_in0), .out(notOp_238_out));

	reg [0:0] andOp_239_in0;
	reg [0:0] andOp_239_in1;
	wire [0:0] andOp_239_out;
	andOp #(.WIDTH(1)) andOp_239(.in0(andOp_239_in0), .in1(andOp_239_in1), .out(andOp_239_out));

	reg [0:0] andOp_240_in0;
	reg [0:0] andOp_240_in1;
	wire [0:0] andOp_240_out;
	andOp #(.WIDTH(1)) andOp_240(.in0(andOp_240_in0), .in1(andOp_240_in1), .out(andOp_240_out));

	reg [31:0] eq_241_in0;
	reg [31:0] eq_241_in1;
	wire [0:0] eq_241_out;
	eq #(.WIDTH(32)) eq_241(.in0(eq_241_in0), .in1(eq_241_in1), .out(eq_241_out));

	reg [0:0] andOp_242_in0;
	reg [0:0] andOp_242_in1;
	wire [0:0] andOp_242_out;
	andOp #(.WIDTH(1)) andOp_242(.in0(andOp_242_in0), .in1(andOp_242_in1), .out(andOp_242_out));

	reg [0:0] notOp_243_in0;
	wire [0:0] notOp_243_out;
	notOp #(.WIDTH(1)) notOp_243(.in(notOp_243_in0), .out(notOp_243_out));

	reg [0:0] andOp_244_in0;
	reg [0:0] andOp_244_in1;
	wire [0:0] andOp_244_out;
	andOp #(.WIDTH(1)) andOp_244(.in0(andOp_244_in0), .in1(andOp_244_in1), .out(andOp_244_out));

	reg [31:0] eq_245_in0;
	reg [31:0] eq_245_in1;
	wire [0:0] eq_245_out;
	eq #(.WIDTH(32)) eq_245(.in0(eq_245_in0), .in1(eq_245_in1), .out(eq_245_out));

	reg [0:0] andOp_246_in0;
	reg [0:0] andOp_246_in1;
	wire [0:0] andOp_246_out;
	andOp #(.WIDTH(1)) andOp_246(.in0(andOp_246_in0), .in1(andOp_246_in1), .out(andOp_246_out));

	reg [0:0] notOp_247_in0;
	wire [0:0] notOp_247_out;
	notOp #(.WIDTH(1)) notOp_247(.in(notOp_247_in0), .out(notOp_247_out));

	reg [0:0] andOp_248_in0;
	reg [0:0] andOp_248_in1;
	wire [0:0] andOp_248_out;
	andOp #(.WIDTH(1)) andOp_248(.in0(andOp_248_in0), .in1(andOp_248_in1), .out(andOp_248_out));

	reg [0:0] andOp_249_in0;
	reg [0:0] andOp_249_in1;
	wire [0:0] andOp_249_out;
	andOp #(.WIDTH(1)) andOp_249(.in0(andOp_249_in0), .in1(andOp_249_in1), .out(andOp_249_out));

	reg [31:0] eq_250_in0;
	reg [31:0] eq_250_in1;
	wire [0:0] eq_250_out;
	eq #(.WIDTH(32)) eq_250(.in0(eq_250_in0), .in1(eq_250_in1), .out(eq_250_out));

	reg [0:0] andOp_251_in0;
	reg [0:0] andOp_251_in1;
	wire [0:0] andOp_251_out;
	andOp #(.WIDTH(1)) andOp_251(.in0(andOp_251_in0), .in1(andOp_251_in1), .out(andOp_251_out));

	reg [0:0] notOp_252_in0;
	wire [0:0] notOp_252_out;
	notOp #(.WIDTH(1)) notOp_252(.in(notOp_252_in0), .out(notOp_252_out));

	reg [0:0] andOp_253_in0;
	reg [0:0] andOp_253_in1;
	wire [0:0] andOp_253_out;
	andOp #(.WIDTH(1)) andOp_253(.in0(andOp_253_in0), .in1(andOp_253_in1), .out(andOp_253_out));

	reg [31:0] eq_254_in0;
	reg [31:0] eq_254_in1;
	wire [0:0] eq_254_out;
	eq #(.WIDTH(32)) eq_254(.in0(eq_254_in0), .in1(eq_254_in1), .out(eq_254_out));

	reg [0:0] andOp_255_in0;
	reg [0:0] andOp_255_in1;
	wire [0:0] andOp_255_out;
	andOp #(.WIDTH(1)) andOp_255(.in0(andOp_255_in0), .in1(andOp_255_in1), .out(andOp_255_out));

	reg [0:0] notOp_256_in0;
	wire [0:0] notOp_256_out;
	notOp #(.WIDTH(1)) notOp_256(.in(notOp_256_in0), .out(notOp_256_out));

	reg [0:0] andOp_257_in0;
	reg [0:0] andOp_257_in1;
	wire [0:0] andOp_257_out;
	andOp #(.WIDTH(1)) andOp_257(.in0(andOp_257_in0), .in1(andOp_257_in1), .out(andOp_257_out));

	reg [0:0] andOp_258_in0;
	reg [0:0] andOp_258_in1;
	wire [0:0] andOp_258_out;
	andOp #(.WIDTH(1)) andOp_258(.in0(andOp_258_in0), .in1(andOp_258_in1), .out(andOp_258_out));

	reg [31:0] eq_259_in0;
	reg [31:0] eq_259_in1;
	wire [0:0] eq_259_out;
	eq #(.WIDTH(32)) eq_259(.in0(eq_259_in0), .in1(eq_259_in1), .out(eq_259_out));

	reg [0:0] andOp_260_in0;
	reg [0:0] andOp_260_in1;
	wire [0:0] andOp_260_out;
	andOp #(.WIDTH(1)) andOp_260(.in0(andOp_260_in0), .in1(andOp_260_in1), .out(andOp_260_out));

	reg [0:0] notOp_261_in0;
	wire [0:0] notOp_261_out;
	notOp #(.WIDTH(1)) notOp_261(.in(notOp_261_in0), .out(notOp_261_out));

	reg [0:0] andOp_262_in0;
	reg [0:0] andOp_262_in1;
	wire [0:0] andOp_262_out;
	andOp #(.WIDTH(1)) andOp_262(.in0(andOp_262_in0), .in1(andOp_262_in1), .out(andOp_262_out));

	reg [31:0] eq_263_in0;
	reg [31:0] eq_263_in1;
	wire [0:0] eq_263_out;
	eq #(.WIDTH(32)) eq_263(.in0(eq_263_in0), .in1(eq_263_in1), .out(eq_263_out));

	reg [0:0] andOp_264_in0;
	reg [0:0] andOp_264_in1;
	wire [0:0] andOp_264_out;
	andOp #(.WIDTH(1)) andOp_264(.in0(andOp_264_in0), .in1(andOp_264_in1), .out(andOp_264_out));

	reg [0:0] notOp_265_in0;
	wire [0:0] notOp_265_out;
	notOp #(.WIDTH(1)) notOp_265(.in(notOp_265_in0), .out(notOp_265_out));

	reg [0:0] andOp_266_in0;
	reg [0:0] andOp_266_in1;
	wire [0:0] andOp_266_out;
	andOp #(.WIDTH(1)) andOp_266(.in0(andOp_266_in0), .in1(andOp_266_in1), .out(andOp_266_out));

	reg [0:0] andOp_267_in0;
	reg [0:0] andOp_267_in1;
	wire [0:0] andOp_267_out;
	andOp #(.WIDTH(1)) andOp_267(.in0(andOp_267_in0), .in1(andOp_267_in1), .out(andOp_267_out));

	reg [31:0] eq_268_in0;
	reg [31:0] eq_268_in1;
	wire [0:0] eq_268_out;
	eq #(.WIDTH(32)) eq_268(.in0(eq_268_in0), .in1(eq_268_in1), .out(eq_268_out));

	reg [0:0] andOp_269_in0;
	reg [0:0] andOp_269_in1;
	wire [0:0] andOp_269_out;
	andOp #(.WIDTH(1)) andOp_269(.in0(andOp_269_in0), .in1(andOp_269_in1), .out(andOp_269_out));

	reg [0:0] notOp_270_in0;
	wire [0:0] notOp_270_out;
	notOp #(.WIDTH(1)) notOp_270(.in(notOp_270_in0), .out(notOp_270_out));

	reg [0:0] andOp_271_in0;
	reg [0:0] andOp_271_in1;
	wire [0:0] andOp_271_out;
	andOp #(.WIDTH(1)) andOp_271(.in0(andOp_271_in0), .in1(andOp_271_in1), .out(andOp_271_out));

	reg [31:0] eq_272_in0;
	reg [31:0] eq_272_in1;
	wire [0:0] eq_272_out;
	eq #(.WIDTH(32)) eq_272(.in0(eq_272_in0), .in1(eq_272_in1), .out(eq_272_out));

	reg [0:0] andOp_273_in0;
	reg [0:0] andOp_273_in1;
	wire [0:0] andOp_273_out;
	andOp #(.WIDTH(1)) andOp_273(.in0(andOp_273_in0), .in1(andOp_273_in1), .out(andOp_273_out));

	reg [0:0] notOp_274_in0;
	wire [0:0] notOp_274_out;
	notOp #(.WIDTH(1)) notOp_274(.in(notOp_274_in0), .out(notOp_274_out));

	reg [0:0] andOp_275_in0;
	reg [0:0] andOp_275_in1;
	wire [0:0] andOp_275_out;
	andOp #(.WIDTH(1)) andOp_275(.in0(andOp_275_in0), .in1(andOp_275_in1), .out(andOp_275_out));

	reg [0:0] andOp_276_in0;
	reg [0:0] andOp_276_in1;
	wire [0:0] andOp_276_out;
	andOp #(.WIDTH(1)) andOp_276(.in0(andOp_276_in0), .in1(andOp_276_in1), .out(andOp_276_out));

	reg [31:0] eq_277_in0;
	reg [31:0] eq_277_in1;
	wire [0:0] eq_277_out;
	eq #(.WIDTH(32)) eq_277(.in0(eq_277_in0), .in1(eq_277_in1), .out(eq_277_out));

	reg [0:0] andOp_278_in0;
	reg [0:0] andOp_278_in1;
	wire [0:0] andOp_278_out;
	andOp #(.WIDTH(1)) andOp_278(.in0(andOp_278_in0), .in1(andOp_278_in1), .out(andOp_278_out));

	reg [0:0] notOp_279_in0;
	wire [0:0] notOp_279_out;
	notOp #(.WIDTH(1)) notOp_279(.in(notOp_279_in0), .out(notOp_279_out));

	reg [0:0] andOp_280_in0;
	reg [0:0] andOp_280_in1;
	wire [0:0] andOp_280_out;
	andOp #(.WIDTH(1)) andOp_280(.in0(andOp_280_in0), .in1(andOp_280_in1), .out(andOp_280_out));

	reg [31:0] eq_281_in0;
	reg [31:0] eq_281_in1;
	wire [0:0] eq_281_out;
	eq #(.WIDTH(32)) eq_281(.in0(eq_281_in0), .in1(eq_281_in1), .out(eq_281_out));

	reg [0:0] andOp_282_in0;
	reg [0:0] andOp_282_in1;
	wire [0:0] andOp_282_out;
	andOp #(.WIDTH(1)) andOp_282(.in0(andOp_282_in0), .in1(andOp_282_in1), .out(andOp_282_out));

	reg [31:0] eq_283_in0;
	reg [31:0] eq_283_in1;
	wire [0:0] eq_283_out;
	eq #(.WIDTH(32)) eq_283(.in0(eq_283_in0), .in1(eq_283_in1), .out(eq_283_out));

	reg [0:0] andOp_284_in0;
	reg [0:0] andOp_284_in1;
	wire [0:0] andOp_284_out;
	andOp #(.WIDTH(1)) andOp_284(.in0(andOp_284_in0), .in1(andOp_284_in1), .out(andOp_284_out));

	reg [0:0] notOp_285_in0;
	wire [0:0] notOp_285_out;
	notOp #(.WIDTH(1)) notOp_285(.in(notOp_285_in0), .out(notOp_285_out));

	reg [0:0] andOp_286_in0;
	reg [0:0] andOp_286_in1;
	wire [0:0] andOp_286_out;
	andOp #(.WIDTH(1)) andOp_286(.in0(andOp_286_in0), .in1(andOp_286_in1), .out(andOp_286_out));

	reg [0:0] andOp_287_in0;
	reg [0:0] andOp_287_in1;
	wire [0:0] andOp_287_out;
	andOp #(.WIDTH(1)) andOp_287(.in0(andOp_287_in0), .in1(andOp_287_in1), .out(andOp_287_out));

	reg [31:0] eq_288_in0;
	reg [31:0] eq_288_in1;
	wire [0:0] eq_288_out;
	eq #(.WIDTH(32)) eq_288(.in0(eq_288_in0), .in1(eq_288_in1), .out(eq_288_out));

	reg [0:0] andOp_289_in0;
	reg [0:0] andOp_289_in1;
	wire [0:0] andOp_289_out;
	andOp #(.WIDTH(1)) andOp_289(.in0(andOp_289_in0), .in1(andOp_289_in1), .out(andOp_289_out));

	reg [0:0] notOp_290_in0;
	wire [0:0] notOp_290_out;
	notOp #(.WIDTH(1)) notOp_290(.in(notOp_290_in0), .out(notOp_290_out));

	reg [0:0] andOp_291_in0;
	reg [0:0] andOp_291_in1;
	wire [0:0] andOp_291_out;
	andOp #(.WIDTH(1)) andOp_291(.in0(andOp_291_in0), .in1(andOp_291_in1), .out(andOp_291_out));

	reg [31:0] eq_292_in0;
	reg [31:0] eq_292_in1;
	wire [0:0] eq_292_out;
	eq #(.WIDTH(32)) eq_292(.in0(eq_292_in0), .in1(eq_292_in1), .out(eq_292_out));

	reg [0:0] andOp_293_in0;
	reg [0:0] andOp_293_in1;
	wire [0:0] andOp_293_out;
	andOp #(.WIDTH(1)) andOp_293(.in0(andOp_293_in0), .in1(andOp_293_in1), .out(andOp_293_out));

	reg [0:0] notOp_294_in0;
	wire [0:0] notOp_294_out;
	notOp #(.WIDTH(1)) notOp_294(.in(notOp_294_in0), .out(notOp_294_out));

	reg [0:0] andOp_295_in0;
	reg [0:0] andOp_295_in1;
	wire [0:0] andOp_295_out;
	andOp #(.WIDTH(1)) andOp_295(.in0(andOp_295_in0), .in1(andOp_295_in1), .out(andOp_295_out));

	reg [0:0] andOp_296_in0;
	reg [0:0] andOp_296_in1;
	wire [0:0] andOp_296_out;
	andOp #(.WIDTH(1)) andOp_296(.in0(andOp_296_in0), .in1(andOp_296_in1), .out(andOp_296_out));

	reg [31:0] eq_297_in0;
	reg [31:0] eq_297_in1;
	wire [0:0] eq_297_out;
	eq #(.WIDTH(32)) eq_297(.in0(eq_297_in0), .in1(eq_297_in1), .out(eq_297_out));

	reg [0:0] andOp_298_in0;
	reg [0:0] andOp_298_in1;
	wire [0:0] andOp_298_out;
	andOp #(.WIDTH(1)) andOp_298(.in0(andOp_298_in0), .in1(andOp_298_in1), .out(andOp_298_out));

	reg [0:0] notOp_299_in0;
	wire [0:0] notOp_299_out;
	notOp #(.WIDTH(1)) notOp_299(.in(notOp_299_in0), .out(notOp_299_out));

	reg [0:0] andOp_300_in0;
	reg [0:0] andOp_300_in1;
	wire [0:0] andOp_300_out;
	andOp #(.WIDTH(1)) andOp_300(.in0(andOp_300_in0), .in1(andOp_300_in1), .out(andOp_300_out));

	reg [31:0] eq_301_in0;
	reg [31:0] eq_301_in1;
	wire [0:0] eq_301_out;
	eq #(.WIDTH(32)) eq_301(.in0(eq_301_in0), .in1(eq_301_in1), .out(eq_301_out));

	reg [0:0] andOp_302_in0;
	reg [0:0] andOp_302_in1;
	wire [0:0] andOp_302_out;
	andOp #(.WIDTH(1)) andOp_302(.in0(andOp_302_in0), .in1(andOp_302_in1), .out(andOp_302_out));

	reg [0:0] notOp_303_in0;
	wire [0:0] notOp_303_out;
	notOp #(.WIDTH(1)) notOp_303(.in(notOp_303_in0), .out(notOp_303_out));

	reg [0:0] andOp_304_in0;
	reg [0:0] andOp_304_in1;
	wire [0:0] andOp_304_out;
	andOp #(.WIDTH(1)) andOp_304(.in0(andOp_304_in0), .in1(andOp_304_in1), .out(andOp_304_out));

	reg [0:0] andOp_305_in0;
	reg [0:0] andOp_305_in1;
	wire [0:0] andOp_305_out;
	andOp #(.WIDTH(1)) andOp_305(.in0(andOp_305_in0), .in1(andOp_305_in1), .out(andOp_305_out));

	reg [31:0] eq_306_in0;
	reg [31:0] eq_306_in1;
	wire [0:0] eq_306_out;
	eq #(.WIDTH(32)) eq_306(.in0(eq_306_in0), .in1(eq_306_in1), .out(eq_306_out));

	reg [0:0] andOp_307_in0;
	reg [0:0] andOp_307_in1;
	wire [0:0] andOp_307_out;
	andOp #(.WIDTH(1)) andOp_307(.in0(andOp_307_in0), .in1(andOp_307_in1), .out(andOp_307_out));

	reg [0:0] notOp_308_in0;
	wire [0:0] notOp_308_out;
	notOp #(.WIDTH(1)) notOp_308(.in(notOp_308_in0), .out(notOp_308_out));

	reg [0:0] andOp_309_in0;
	reg [0:0] andOp_309_in1;
	wire [0:0] andOp_309_out;
	andOp #(.WIDTH(1)) andOp_309(.in0(andOp_309_in0), .in1(andOp_309_in1), .out(andOp_309_out));

	reg [31:0] eq_310_in0;
	reg [31:0] eq_310_in1;
	wire [0:0] eq_310_out;
	eq #(.WIDTH(32)) eq_310(.in0(eq_310_in0), .in1(eq_310_in1), .out(eq_310_out));

	reg [0:0] andOp_311_in0;
	reg [0:0] andOp_311_in1;
	wire [0:0] andOp_311_out;
	andOp #(.WIDTH(1)) andOp_311(.in0(andOp_311_in0), .in1(andOp_311_in1), .out(andOp_311_out));

	reg [0:0] notOp_312_in0;
	wire [0:0] notOp_312_out;
	notOp #(.WIDTH(1)) notOp_312(.in(notOp_312_in0), .out(notOp_312_out));

	reg [0:0] andOp_313_in0;
	reg [0:0] andOp_313_in1;
	wire [0:0] andOp_313_out;
	andOp #(.WIDTH(1)) andOp_313(.in0(andOp_313_in0), .in1(andOp_313_in1), .out(andOp_313_out));

	reg [0:0] andOp_314_in0;
	reg [0:0] andOp_314_in1;
	wire [0:0] andOp_314_out;
	andOp #(.WIDTH(1)) andOp_314(.in0(andOp_314_in0), .in1(andOp_314_in1), .out(andOp_314_out));

	reg [31:0] eq_315_in0;
	reg [31:0] eq_315_in1;
	wire [0:0] eq_315_out;
	eq #(.WIDTH(32)) eq_315(.in0(eq_315_in0), .in1(eq_315_in1), .out(eq_315_out));

	reg [0:0] andOp_316_in0;
	reg [0:0] andOp_316_in1;
	wire [0:0] andOp_316_out;
	andOp #(.WIDTH(1)) andOp_316(.in0(andOp_316_in0), .in1(andOp_316_in1), .out(andOp_316_out));

	reg [0:0] notOp_317_in0;
	wire [0:0] notOp_317_out;
	notOp #(.WIDTH(1)) notOp_317(.in(notOp_317_in0), .out(notOp_317_out));

	reg [0:0] andOp_318_in0;
	reg [0:0] andOp_318_in1;
	wire [0:0] andOp_318_out;
	andOp #(.WIDTH(1)) andOp_318(.in0(andOp_318_in0), .in1(andOp_318_in1), .out(andOp_318_out));

	reg [31:0] eq_319_in0;
	reg [31:0] eq_319_in1;
	wire [0:0] eq_319_out;
	eq #(.WIDTH(32)) eq_319(.in0(eq_319_in0), .in1(eq_319_in1), .out(eq_319_out));

	reg [0:0] andOp_320_in0;
	reg [0:0] andOp_320_in1;
	wire [0:0] andOp_320_out;
	andOp #(.WIDTH(1)) andOp_320(.in0(andOp_320_in0), .in1(andOp_320_in1), .out(andOp_320_out));

	reg [0:0] notOp_321_in0;
	wire [0:0] notOp_321_out;
	notOp #(.WIDTH(1)) notOp_321(.in(notOp_321_in0), .out(notOp_321_out));

	reg [0:0] andOp_322_in0;
	reg [0:0] andOp_322_in1;
	wire [0:0] andOp_322_out;
	andOp #(.WIDTH(1)) andOp_322(.in0(andOp_322_in0), .in1(andOp_322_in1), .out(andOp_322_out));

	reg [0:0] andOp_323_in0;
	reg [0:0] andOp_323_in1;
	wire [0:0] andOp_323_out;
	andOp #(.WIDTH(1)) andOp_323(.in0(andOp_323_in0), .in1(andOp_323_in1), .out(andOp_323_out));

	reg [31:0] eq_324_in0;
	reg [31:0] eq_324_in1;
	wire [0:0] eq_324_out;
	eq #(.WIDTH(32)) eq_324(.in0(eq_324_in0), .in1(eq_324_in1), .out(eq_324_out));

	reg [0:0] andOp_325_in0;
	reg [0:0] andOp_325_in1;
	wire [0:0] andOp_325_out;
	andOp #(.WIDTH(1)) andOp_325(.in0(andOp_325_in0), .in1(andOp_325_in1), .out(andOp_325_out));

	reg [0:0] notOp_326_in0;
	wire [0:0] notOp_326_out;
	notOp #(.WIDTH(1)) notOp_326(.in(notOp_326_in0), .out(notOp_326_out));

	reg [0:0] andOp_327_in0;
	reg [0:0] andOp_327_in1;
	wire [0:0] andOp_327_out;
	andOp #(.WIDTH(1)) andOp_327(.in0(andOp_327_in0), .in1(andOp_327_in1), .out(andOp_327_out));

	reg [31:0] eq_328_in0;
	reg [31:0] eq_328_in1;
	wire [0:0] eq_328_out;
	eq #(.WIDTH(32)) eq_328(.in0(eq_328_in0), .in1(eq_328_in1), .out(eq_328_out));

	reg [0:0] andOp_329_in0;
	reg [0:0] andOp_329_in1;
	wire [0:0] andOp_329_out;
	andOp #(.WIDTH(1)) andOp_329(.in0(andOp_329_in0), .in1(andOp_329_in1), .out(andOp_329_out));

	reg [0:0] notOp_330_in0;
	wire [0:0] notOp_330_out;
	notOp #(.WIDTH(1)) notOp_330(.in(notOp_330_in0), .out(notOp_330_out));

	reg [0:0] andOp_331_in0;
	reg [0:0] andOp_331_in1;
	wire [0:0] andOp_331_out;
	andOp #(.WIDTH(1)) andOp_331(.in0(andOp_331_in0), .in1(andOp_331_in1), .out(andOp_331_out));

	reg [0:0] andOp_332_in0;
	reg [0:0] andOp_332_in1;
	wire [0:0] andOp_332_out;
	andOp #(.WIDTH(1)) andOp_332(.in0(andOp_332_in0), .in1(andOp_332_in1), .out(andOp_332_out));

	reg [31:0] eq_333_in0;
	reg [31:0] eq_333_in1;
	wire [0:0] eq_333_out;
	eq #(.WIDTH(32)) eq_333(.in0(eq_333_in0), .in1(eq_333_in1), .out(eq_333_out));

	reg [0:0] andOp_334_in0;
	reg [0:0] andOp_334_in1;
	wire [0:0] andOp_334_out;
	andOp #(.WIDTH(1)) andOp_334(.in0(andOp_334_in0), .in1(andOp_334_in1), .out(andOp_334_out));

	reg [0:0] notOp_335_in0;
	wire [0:0] notOp_335_out;
	notOp #(.WIDTH(1)) notOp_335(.in(notOp_335_in0), .out(notOp_335_out));

	reg [0:0] andOp_336_in0;
	reg [0:0] andOp_336_in1;
	wire [0:0] andOp_336_out;
	andOp #(.WIDTH(1)) andOp_336(.in0(andOp_336_in0), .in1(andOp_336_in1), .out(andOp_336_out));

	reg [31:0] eq_337_in0;
	reg [31:0] eq_337_in1;
	wire [0:0] eq_337_out;
	eq #(.WIDTH(32)) eq_337(.in0(eq_337_in0), .in1(eq_337_in1), .out(eq_337_out));

	reg [0:0] andOp_338_in0;
	reg [0:0] andOp_338_in1;
	wire [0:0] andOp_338_out;
	andOp #(.WIDTH(1)) andOp_338(.in0(andOp_338_in0), .in1(andOp_338_in1), .out(andOp_338_out));

	reg [0:0] notOp_339_in0;
	wire [0:0] notOp_339_out;
	notOp #(.WIDTH(1)) notOp_339(.in(notOp_339_in0), .out(notOp_339_out));

	reg [0:0] andOp_340_in0;
	reg [0:0] andOp_340_in1;
	wire [0:0] andOp_340_out;
	andOp #(.WIDTH(1)) andOp_340(.in0(andOp_340_in0), .in1(andOp_340_in1), .out(andOp_340_out));

	reg [0:0] andOp_341_in0;
	reg [0:0] andOp_341_in1;
	wire [0:0] andOp_341_out;
	andOp #(.WIDTH(1)) andOp_341(.in0(andOp_341_in0), .in1(andOp_341_in1), .out(andOp_341_out));

	reg [31:0] eq_342_in0;
	reg [31:0] eq_342_in1;
	wire [0:0] eq_342_out;
	eq #(.WIDTH(32)) eq_342(.in0(eq_342_in0), .in1(eq_342_in1), .out(eq_342_out));

	reg [0:0] andOp_343_in0;
	reg [0:0] andOp_343_in1;
	wire [0:0] andOp_343_out;
	andOp #(.WIDTH(1)) andOp_343(.in0(andOp_343_in0), .in1(andOp_343_in1), .out(andOp_343_out));

	reg [0:0] notOp_344_in0;
	wire [0:0] notOp_344_out;
	notOp #(.WIDTH(1)) notOp_344(.in(notOp_344_in0), .out(notOp_344_out));

	reg [0:0] andOp_345_in0;
	reg [0:0] andOp_345_in1;
	wire [0:0] andOp_345_out;
	andOp #(.WIDTH(1)) andOp_345(.in0(andOp_345_in0), .in1(andOp_345_in1), .out(andOp_345_out));

	reg [31:0] eq_346_in0;
	reg [31:0] eq_346_in1;
	wire [0:0] eq_346_out;
	eq #(.WIDTH(32)) eq_346(.in0(eq_346_in0), .in1(eq_346_in1), .out(eq_346_out));

	reg [0:0] andOp_347_in0;
	reg [0:0] andOp_347_in1;
	wire [0:0] andOp_347_out;
	andOp #(.WIDTH(1)) andOp_347(.in0(andOp_347_in0), .in1(andOp_347_in1), .out(andOp_347_out));

	reg [0:0] notOp_348_in0;
	wire [0:0] notOp_348_out;
	notOp #(.WIDTH(1)) notOp_348(.in(notOp_348_in0), .out(notOp_348_out));

	reg [0:0] andOp_349_in0;
	reg [0:0] andOp_349_in1;
	wire [0:0] andOp_349_out;
	andOp #(.WIDTH(1)) andOp_349(.in0(andOp_349_in0), .in1(andOp_349_in1), .out(andOp_349_out));

	reg [0:0] andOp_350_in0;
	reg [0:0] andOp_350_in1;
	wire [0:0] andOp_350_out;
	andOp #(.WIDTH(1)) andOp_350(.in0(andOp_350_in0), .in1(andOp_350_in1), .out(andOp_350_out));

	reg [31:0] eq_351_in0;
	reg [31:0] eq_351_in1;
	wire [0:0] eq_351_out;
	eq #(.WIDTH(32)) eq_351(.in0(eq_351_in0), .in1(eq_351_in1), .out(eq_351_out));

	reg [0:0] andOp_352_in0;
	reg [0:0] andOp_352_in1;
	wire [0:0] andOp_352_out;
	andOp #(.WIDTH(1)) andOp_352(.in0(andOp_352_in0), .in1(andOp_352_in1), .out(andOp_352_out));

	reg [0:0] notOp_353_in0;
	wire [0:0] notOp_353_out;
	notOp #(.WIDTH(1)) notOp_353(.in(notOp_353_in0), .out(notOp_353_out));

	reg [0:0] andOp_354_in0;
	reg [0:0] andOp_354_in1;
	wire [0:0] andOp_354_out;
	andOp #(.WIDTH(1)) andOp_354(.in0(andOp_354_in0), .in1(andOp_354_in1), .out(andOp_354_out));

	reg [31:0] eq_355_in0;
	reg [31:0] eq_355_in1;
	wire [0:0] eq_355_out;
	eq #(.WIDTH(32)) eq_355(.in0(eq_355_in0), .in1(eq_355_in1), .out(eq_355_out));

	reg [0:0] andOp_356_in0;
	reg [0:0] andOp_356_in1;
	wire [0:0] andOp_356_out;
	andOp #(.WIDTH(1)) andOp_356(.in0(andOp_356_in0), .in1(andOp_356_in1), .out(andOp_356_out));

	reg [0:0] notOp_357_in0;
	wire [0:0] notOp_357_out;
	notOp #(.WIDTH(1)) notOp_357(.in(notOp_357_in0), .out(notOp_357_out));

	reg [0:0] andOp_358_in0;
	reg [0:0] andOp_358_in1;
	wire [0:0] andOp_358_out;
	andOp #(.WIDTH(1)) andOp_358(.in0(andOp_358_in0), .in1(andOp_358_in1), .out(andOp_358_out));

	reg [0:0] andOp_359_in0;
	reg [0:0] andOp_359_in1;
	wire [0:0] andOp_359_out;
	andOp #(.WIDTH(1)) andOp_359(.in0(andOp_359_in0), .in1(andOp_359_in1), .out(andOp_359_out));

	reg [31:0] eq_360_in0;
	reg [31:0] eq_360_in1;
	wire [0:0] eq_360_out;
	eq #(.WIDTH(32)) eq_360(.in0(eq_360_in0), .in1(eq_360_in1), .out(eq_360_out));

	reg [0:0] andOp_361_in0;
	reg [0:0] andOp_361_in1;
	wire [0:0] andOp_361_out;
	andOp #(.WIDTH(1)) andOp_361(.in0(andOp_361_in0), .in1(andOp_361_in1), .out(andOp_361_out));

	reg [0:0] notOp_362_in0;
	wire [0:0] notOp_362_out;
	notOp #(.WIDTH(1)) notOp_362(.in(notOp_362_in0), .out(notOp_362_out));

	reg [0:0] andOp_363_in0;
	reg [0:0] andOp_363_in1;
	wire [0:0] andOp_363_out;
	andOp #(.WIDTH(1)) andOp_363(.in0(andOp_363_in0), .in1(andOp_363_in1), .out(andOp_363_out));

	reg [31:0] eq_364_in0;
	reg [31:0] eq_364_in1;
	wire [0:0] eq_364_out;
	eq #(.WIDTH(32)) eq_364(.in0(eq_364_in0), .in1(eq_364_in1), .out(eq_364_out));

	reg [0:0] andOp_365_in0;
	reg [0:0] andOp_365_in1;
	wire [0:0] andOp_365_out;
	andOp #(.WIDTH(1)) andOp_365(.in0(andOp_365_in0), .in1(andOp_365_in1), .out(andOp_365_out));

	reg [31:0] eq_366_in0;
	reg [31:0] eq_366_in1;
	wire [0:0] eq_366_out;
	eq #(.WIDTH(32)) eq_366(.in0(eq_366_in0), .in1(eq_366_in1), .out(eq_366_out));

	reg [0:0] andOp_367_in0;
	reg [0:0] andOp_367_in1;
	wire [0:0] andOp_367_out;
	andOp #(.WIDTH(1)) andOp_367(.in0(andOp_367_in0), .in1(andOp_367_in1), .out(andOp_367_out));

	reg [0:0] notOp_368_in0;
	wire [0:0] notOp_368_out;
	notOp #(.WIDTH(1)) notOp_368(.in(notOp_368_in0), .out(notOp_368_out));

	reg [0:0] andOp_369_in0;
	reg [0:0] andOp_369_in1;
	wire [0:0] andOp_369_out;
	andOp #(.WIDTH(1)) andOp_369(.in0(andOp_369_in0), .in1(andOp_369_in1), .out(andOp_369_out));

	reg [0:0] andOp_370_in0;
	reg [0:0] andOp_370_in1;
	wire [0:0] andOp_370_out;
	andOp #(.WIDTH(1)) andOp_370(.in0(andOp_370_in0), .in1(andOp_370_in1), .out(andOp_370_out));

	reg [31:0] eq_371_in0;
	reg [31:0] eq_371_in1;
	wire [0:0] eq_371_out;
	eq #(.WIDTH(32)) eq_371(.in0(eq_371_in0), .in1(eq_371_in1), .out(eq_371_out));

	reg [0:0] andOp_372_in0;
	reg [0:0] andOp_372_in1;
	wire [0:0] andOp_372_out;
	andOp #(.WIDTH(1)) andOp_372(.in0(andOp_372_in0), .in1(andOp_372_in1), .out(andOp_372_out));

	reg [0:0] notOp_373_in0;
	wire [0:0] notOp_373_out;
	notOp #(.WIDTH(1)) notOp_373(.in(notOp_373_in0), .out(notOp_373_out));

	reg [0:0] andOp_374_in0;
	reg [0:0] andOp_374_in1;
	wire [0:0] andOp_374_out;
	andOp #(.WIDTH(1)) andOp_374(.in0(andOp_374_in0), .in1(andOp_374_in1), .out(andOp_374_out));

	reg [31:0] eq_375_in0;
	reg [31:0] eq_375_in1;
	wire [0:0] eq_375_out;
	eq #(.WIDTH(32)) eq_375(.in0(eq_375_in0), .in1(eq_375_in1), .out(eq_375_out));

	reg [0:0] andOp_376_in0;
	reg [0:0] andOp_376_in1;
	wire [0:0] andOp_376_out;
	andOp #(.WIDTH(1)) andOp_376(.in0(andOp_376_in0), .in1(andOp_376_in1), .out(andOp_376_out));

	reg [31:0] eq_377_in0;
	reg [31:0] eq_377_in1;
	wire [0:0] eq_377_out;
	eq #(.WIDTH(32)) eq_377(.in0(eq_377_in0), .in1(eq_377_in1), .out(eq_377_out));

	reg [0:0] andOp_378_in0;
	reg [0:0] andOp_378_in1;
	wire [0:0] andOp_378_out;
	andOp #(.WIDTH(1)) andOp_378(.in0(andOp_378_in0), .in1(andOp_378_in1), .out(andOp_378_out));

	reg [0:0] notOp_379_in0;
	wire [0:0] notOp_379_out;
	notOp #(.WIDTH(1)) notOp_379(.in(notOp_379_in0), .out(notOp_379_out));

	reg [0:0] andOp_380_in0;
	reg [0:0] andOp_380_in1;
	wire [0:0] andOp_380_out;
	andOp #(.WIDTH(1)) andOp_380(.in0(andOp_380_in0), .in1(andOp_380_in1), .out(andOp_380_out));

	reg [0:0] andOp_381_in0;
	reg [0:0] andOp_381_in1;
	wire [0:0] andOp_381_out;
	andOp #(.WIDTH(1)) andOp_381(.in0(andOp_381_in0), .in1(andOp_381_in1), .out(andOp_381_out));

	reg [31:0] eq_382_in0;
	reg [31:0] eq_382_in1;
	wire [0:0] eq_382_out;
	eq #(.WIDTH(32)) eq_382(.in0(eq_382_in0), .in1(eq_382_in1), .out(eq_382_out));

	reg [0:0] andOp_383_in0;
	reg [0:0] andOp_383_in1;
	wire [0:0] andOp_383_out;
	andOp #(.WIDTH(1)) andOp_383(.in0(andOp_383_in0), .in1(andOp_383_in1), .out(andOp_383_out));

	reg [0:0] notOp_384_in0;
	wire [0:0] notOp_384_out;
	notOp #(.WIDTH(1)) notOp_384(.in(notOp_384_in0), .out(notOp_384_out));

	reg [0:0] andOp_385_in0;
	reg [0:0] andOp_385_in1;
	wire [0:0] andOp_385_out;
	andOp #(.WIDTH(1)) andOp_385(.in0(andOp_385_in0), .in1(andOp_385_in1), .out(andOp_385_out));

	reg [31:0] eq_386_in0;
	reg [31:0] eq_386_in1;
	wire [0:0] eq_386_out;
	eq #(.WIDTH(32)) eq_386(.in0(eq_386_in0), .in1(eq_386_in1), .out(eq_386_out));

	reg [0:0] andOp_387_in0;
	reg [0:0] andOp_387_in1;
	wire [0:0] andOp_387_out;
	andOp #(.WIDTH(1)) andOp_387(.in0(andOp_387_in0), .in1(andOp_387_in1), .out(andOp_387_out));

	reg [0:0] notOp_388_in0;
	wire [0:0] notOp_388_out;
	notOp #(.WIDTH(1)) notOp_388(.in(notOp_388_in0), .out(notOp_388_out));

	reg [0:0] andOp_389_in0;
	reg [0:0] andOp_389_in1;
	wire [0:0] andOp_389_out;
	andOp #(.WIDTH(1)) andOp_389(.in0(andOp_389_in0), .in1(andOp_389_in1), .out(andOp_389_out));

	reg [0:0] andOp_390_in0;
	reg [0:0] andOp_390_in1;
	wire [0:0] andOp_390_out;
	andOp #(.WIDTH(1)) andOp_390(.in0(andOp_390_in0), .in1(andOp_390_in1), .out(andOp_390_out));

	reg [31:0] eq_391_in0;
	reg [31:0] eq_391_in1;
	wire [0:0] eq_391_out;
	eq #(.WIDTH(32)) eq_391(.in0(eq_391_in0), .in1(eq_391_in1), .out(eq_391_out));

	reg [0:0] andOp_392_in0;
	reg [0:0] andOp_392_in1;
	wire [0:0] andOp_392_out;
	andOp #(.WIDTH(1)) andOp_392(.in0(andOp_392_in0), .in1(andOp_392_in1), .out(andOp_392_out));

	reg [0:0] notOp_393_in0;
	wire [0:0] notOp_393_out;
	notOp #(.WIDTH(1)) notOp_393(.in(notOp_393_in0), .out(notOp_393_out));

	reg [0:0] andOp_394_in0;
	reg [0:0] andOp_394_in1;
	wire [0:0] andOp_394_out;
	andOp #(.WIDTH(1)) andOp_394(.in0(andOp_394_in0), .in1(andOp_394_in1), .out(andOp_394_out));

	reg [31:0] eq_395_in0;
	reg [31:0] eq_395_in1;
	wire [0:0] eq_395_out;
	eq #(.WIDTH(32)) eq_395(.in0(eq_395_in0), .in1(eq_395_in1), .out(eq_395_out));

	reg [0:0] andOp_396_in0;
	reg [0:0] andOp_396_in1;
	wire [0:0] andOp_396_out;
	andOp #(.WIDTH(1)) andOp_396(.in0(andOp_396_in0), .in1(andOp_396_in1), .out(andOp_396_out));

	reg [31:0] eq_397_in0;
	reg [31:0] eq_397_in1;
	wire [0:0] eq_397_out;
	eq #(.WIDTH(32)) eq_397(.in0(eq_397_in0), .in1(eq_397_in1), .out(eq_397_out));

	reg [0:0] andOp_398_in0;
	reg [0:0] andOp_398_in1;
	wire [0:0] andOp_398_out;
	andOp #(.WIDTH(1)) andOp_398(.in0(andOp_398_in0), .in1(andOp_398_in1), .out(andOp_398_out));

	reg [0:0] notOp_399_in0;
	wire [0:0] notOp_399_out;
	notOp #(.WIDTH(1)) notOp_399(.in(notOp_399_in0), .out(notOp_399_out));

	reg [0:0] andOp_400_in0;
	reg [0:0] andOp_400_in1;
	wire [0:0] andOp_400_out;
	andOp #(.WIDTH(1)) andOp_400(.in0(andOp_400_in0), .in1(andOp_400_in1), .out(andOp_400_out));

	reg [0:0] andOp_401_in0;
	reg [0:0] andOp_401_in1;
	wire [0:0] andOp_401_out;
	andOp #(.WIDTH(1)) andOp_401(.in0(andOp_401_in0), .in1(andOp_401_in1), .out(andOp_401_out));

	reg [31:0] eq_402_in0;
	reg [31:0] eq_402_in1;
	wire [0:0] eq_402_out;
	eq #(.WIDTH(32)) eq_402(.in0(eq_402_in0), .in1(eq_402_in1), .out(eq_402_out));

	reg [0:0] andOp_403_in0;
	reg [0:0] andOp_403_in1;
	wire [0:0] andOp_403_out;
	andOp #(.WIDTH(1)) andOp_403(.in0(andOp_403_in0), .in1(andOp_403_in1), .out(andOp_403_out));

	reg [0:0] notOp_404_in0;
	wire [0:0] notOp_404_out;
	notOp #(.WIDTH(1)) notOp_404(.in(notOp_404_in0), .out(notOp_404_out));

	reg [0:0] andOp_405_in0;
	reg [0:0] andOp_405_in1;
	wire [0:0] andOp_405_out;
	andOp #(.WIDTH(1)) andOp_405(.in0(andOp_405_in0), .in1(andOp_405_in1), .out(andOp_405_out));

	reg [31:0] eq_406_in0;
	reg [31:0] eq_406_in1;
	wire [0:0] eq_406_out;
	eq #(.WIDTH(32)) eq_406(.in0(eq_406_in0), .in1(eq_406_in1), .out(eq_406_out));

	reg [0:0] andOp_407_in0;
	reg [0:0] andOp_407_in1;
	wire [0:0] andOp_407_out;
	andOp #(.WIDTH(1)) andOp_407(.in0(andOp_407_in0), .in1(andOp_407_in1), .out(andOp_407_out));

	reg [0:0] notOp_408_in0;
	wire [0:0] notOp_408_out;
	notOp #(.WIDTH(1)) notOp_408(.in(notOp_408_in0), .out(notOp_408_out));

	reg [0:0] andOp_409_in0;
	reg [0:0] andOp_409_in1;
	wire [0:0] andOp_409_out;
	andOp #(.WIDTH(1)) andOp_409(.in0(andOp_409_in0), .in1(andOp_409_in1), .out(andOp_409_out));

	reg [0:0] andOp_410_in0;
	reg [0:0] andOp_410_in1;
	wire [0:0] andOp_410_out;
	andOp #(.WIDTH(1)) andOp_410(.in0(andOp_410_in0), .in1(andOp_410_in1), .out(andOp_410_out));

	reg [31:0] eq_411_in0;
	reg [31:0] eq_411_in1;
	wire [0:0] eq_411_out;
	eq #(.WIDTH(32)) eq_411(.in0(eq_411_in0), .in1(eq_411_in1), .out(eq_411_out));

	reg [0:0] andOp_412_in0;
	reg [0:0] andOp_412_in1;
	wire [0:0] andOp_412_out;
	andOp #(.WIDTH(1)) andOp_412(.in0(andOp_412_in0), .in1(andOp_412_in1), .out(andOp_412_out));

	reg [0:0] notOp_413_in0;
	wire [0:0] notOp_413_out;
	notOp #(.WIDTH(1)) notOp_413(.in(notOp_413_in0), .out(notOp_413_out));

	reg [0:0] andOp_414_in0;
	reg [0:0] andOp_414_in1;
	wire [0:0] andOp_414_out;
	andOp #(.WIDTH(1)) andOp_414(.in0(andOp_414_in0), .in1(andOp_414_in1), .out(andOp_414_out));

	reg [31:0] eq_415_in0;
	reg [31:0] eq_415_in1;
	wire [0:0] eq_415_out;
	eq #(.WIDTH(32)) eq_415(.in0(eq_415_in0), .in1(eq_415_in1), .out(eq_415_out));

	reg [0:0] andOp_416_in0;
	reg [0:0] andOp_416_in1;
	wire [0:0] andOp_416_out;
	andOp #(.WIDTH(1)) andOp_416(.in0(andOp_416_in0), .in1(andOp_416_in1), .out(andOp_416_out));

	reg [0:0] notOp_417_in0;
	wire [0:0] notOp_417_out;
	notOp #(.WIDTH(1)) notOp_417(.in(notOp_417_in0), .out(notOp_417_out));

	reg [0:0] andOp_418_in0;
	reg [0:0] andOp_418_in1;
	wire [0:0] andOp_418_out;
	andOp #(.WIDTH(1)) andOp_418(.in0(andOp_418_in0), .in1(andOp_418_in1), .out(andOp_418_out));

	reg [0:0] andOp_419_in0;
	reg [0:0] andOp_419_in1;
	wire [0:0] andOp_419_out;
	andOp #(.WIDTH(1)) andOp_419(.in0(andOp_419_in0), .in1(andOp_419_in1), .out(andOp_419_out));

	reg [31:0] eq_420_in0;
	reg [31:0] eq_420_in1;
	wire [0:0] eq_420_out;
	eq #(.WIDTH(32)) eq_420(.in0(eq_420_in0), .in1(eq_420_in1), .out(eq_420_out));

	reg [0:0] andOp_421_in0;
	reg [0:0] andOp_421_in1;
	wire [0:0] andOp_421_out;
	andOp #(.WIDTH(1)) andOp_421(.in0(andOp_421_in0), .in1(andOp_421_in1), .out(andOp_421_out));

	reg [0:0] notOp_422_in0;
	wire [0:0] notOp_422_out;
	notOp #(.WIDTH(1)) notOp_422(.in(notOp_422_in0), .out(notOp_422_out));

	reg [0:0] andOp_423_in0;
	reg [0:0] andOp_423_in1;
	wire [0:0] andOp_423_out;
	andOp #(.WIDTH(1)) andOp_423(.in0(andOp_423_in0), .in1(andOp_423_in1), .out(andOp_423_out));

	reg [31:0] eq_424_in0;
	reg [31:0] eq_424_in1;
	wire [0:0] eq_424_out;
	eq #(.WIDTH(32)) eq_424(.in0(eq_424_in0), .in1(eq_424_in1), .out(eq_424_out));

	reg [0:0] andOp_425_in0;
	reg [0:0] andOp_425_in1;
	wire [0:0] andOp_425_out;
	andOp #(.WIDTH(1)) andOp_425(.in0(andOp_425_in0), .in1(andOp_425_in1), .out(andOp_425_out));

	reg [0:0] notOp_426_in0;
	wire [0:0] notOp_426_out;
	notOp #(.WIDTH(1)) notOp_426(.in(notOp_426_in0), .out(notOp_426_out));

	reg [0:0] andOp_427_in0;
	reg [0:0] andOp_427_in1;
	wire [0:0] andOp_427_out;
	andOp #(.WIDTH(1)) andOp_427(.in0(andOp_427_in0), .in1(andOp_427_in1), .out(andOp_427_out));

	reg [0:0] andOp_428_in0;
	reg [0:0] andOp_428_in1;
	wire [0:0] andOp_428_out;
	andOp #(.WIDTH(1)) andOp_428(.in0(andOp_428_in0), .in1(andOp_428_in1), .out(andOp_428_out));

	reg [31:0] eq_429_in0;
	reg [31:0] eq_429_in1;
	wire [0:0] eq_429_out;
	eq #(.WIDTH(32)) eq_429(.in0(eq_429_in0), .in1(eq_429_in1), .out(eq_429_out));

	reg [0:0] andOp_430_in0;
	reg [0:0] andOp_430_in1;
	wire [0:0] andOp_430_out;
	andOp #(.WIDTH(1)) andOp_430(.in0(andOp_430_in0), .in1(andOp_430_in1), .out(andOp_430_out));

	reg [0:0] notOp_431_in0;
	wire [0:0] notOp_431_out;
	notOp #(.WIDTH(1)) notOp_431(.in(notOp_431_in0), .out(notOp_431_out));

	reg [0:0] andOp_432_in0;
	reg [0:0] andOp_432_in1;
	wire [0:0] andOp_432_out;
	andOp #(.WIDTH(1)) andOp_432(.in0(andOp_432_in0), .in1(andOp_432_in1), .out(andOp_432_out));

	reg [31:0] eq_433_in0;
	reg [31:0] eq_433_in1;
	wire [0:0] eq_433_out;
	eq #(.WIDTH(32)) eq_433(.in0(eq_433_in0), .in1(eq_433_in1), .out(eq_433_out));

	reg [0:0] andOp_434_in0;
	reg [0:0] andOp_434_in1;
	wire [0:0] andOp_434_out;
	andOp #(.WIDTH(1)) andOp_434(.in0(andOp_434_in0), .in1(andOp_434_in1), .out(andOp_434_out));

	reg [0:0] notOp_435_in0;
	wire [0:0] notOp_435_out;
	notOp #(.WIDTH(1)) notOp_435(.in(notOp_435_in0), .out(notOp_435_out));

	reg [0:0] andOp_436_in0;
	reg [0:0] andOp_436_in1;
	wire [0:0] andOp_436_out;
	andOp #(.WIDTH(1)) andOp_436(.in0(andOp_436_in0), .in1(andOp_436_in1), .out(andOp_436_out));

	reg [0:0] andOp_437_in0;
	reg [0:0] andOp_437_in1;
	wire [0:0] andOp_437_out;
	andOp #(.WIDTH(1)) andOp_437(.in0(andOp_437_in0), .in1(andOp_437_in1), .out(andOp_437_out));

	reg [31:0] eq_438_in0;
	reg [31:0] eq_438_in1;
	wire [0:0] eq_438_out;
	eq #(.WIDTH(32)) eq_438(.in0(eq_438_in0), .in1(eq_438_in1), .out(eq_438_out));

	reg [0:0] andOp_439_in0;
	reg [0:0] andOp_439_in1;
	wire [0:0] andOp_439_out;
	andOp #(.WIDTH(1)) andOp_439(.in0(andOp_439_in0), .in1(andOp_439_in1), .out(andOp_439_out));

	reg [0:0] notOp_440_in0;
	wire [0:0] notOp_440_out;
	notOp #(.WIDTH(1)) notOp_440(.in(notOp_440_in0), .out(notOp_440_out));

	reg [0:0] andOp_441_in0;
	reg [0:0] andOp_441_in1;
	wire [0:0] andOp_441_out;
	andOp #(.WIDTH(1)) andOp_441(.in0(andOp_441_in0), .in1(andOp_441_in1), .out(andOp_441_out));

	reg [31:0] eq_442_in0;
	reg [31:0] eq_442_in1;
	wire [0:0] eq_442_out;
	eq #(.WIDTH(32)) eq_442(.in0(eq_442_in0), .in1(eq_442_in1), .out(eq_442_out));

	reg [0:0] andOp_443_in0;
	reg [0:0] andOp_443_in1;
	wire [0:0] andOp_443_out;
	andOp #(.WIDTH(1)) andOp_443(.in0(andOp_443_in0), .in1(andOp_443_in1), .out(andOp_443_out));

	reg [0:0] notOp_444_in0;
	wire [0:0] notOp_444_out;
	notOp #(.WIDTH(1)) notOp_444(.in(notOp_444_in0), .out(notOp_444_out));

	reg [0:0] andOp_445_in0;
	reg [0:0] andOp_445_in1;
	wire [0:0] andOp_445_out;
	andOp #(.WIDTH(1)) andOp_445(.in0(andOp_445_in0), .in1(andOp_445_in1), .out(andOp_445_out));

	reg [0:0] andOp_446_in0;
	reg [0:0] andOp_446_in1;
	wire [0:0] andOp_446_out;
	andOp #(.WIDTH(1)) andOp_446(.in0(andOp_446_in0), .in1(andOp_446_in1), .out(andOp_446_out));

	reg [31:0] eq_447_in0;
	reg [31:0] eq_447_in1;
	wire [0:0] eq_447_out;
	eq #(.WIDTH(32)) eq_447(.in0(eq_447_in0), .in1(eq_447_in1), .out(eq_447_out));

	reg [0:0] andOp_448_in0;
	reg [0:0] andOp_448_in1;
	wire [0:0] andOp_448_out;
	andOp #(.WIDTH(1)) andOp_448(.in0(andOp_448_in0), .in1(andOp_448_in1), .out(andOp_448_out));

	reg [0:0] notOp_449_in0;
	wire [0:0] notOp_449_out;
	notOp #(.WIDTH(1)) notOp_449(.in(notOp_449_in0), .out(notOp_449_out));

	reg [0:0] andOp_450_in0;
	reg [0:0] andOp_450_in1;
	wire [0:0] andOp_450_out;
	andOp #(.WIDTH(1)) andOp_450(.in0(andOp_450_in0), .in1(andOp_450_in1), .out(andOp_450_out));

	reg [31:0] eq_451_in0;
	reg [31:0] eq_451_in1;
	wire [0:0] eq_451_out;
	eq #(.WIDTH(32)) eq_451(.in0(eq_451_in0), .in1(eq_451_in1), .out(eq_451_out));

	reg [0:0] andOp_452_in0;
	reg [0:0] andOp_452_in1;
	wire [0:0] andOp_452_out;
	andOp #(.WIDTH(1)) andOp_452(.in0(andOp_452_in0), .in1(andOp_452_in1), .out(andOp_452_out));

	reg [31:0] eq_453_in0;
	reg [31:0] eq_453_in1;
	wire [0:0] eq_453_out;
	eq #(.WIDTH(32)) eq_453(.in0(eq_453_in0), .in1(eq_453_in1), .out(eq_453_out));

	reg [0:0] andOp_454_in0;
	reg [0:0] andOp_454_in1;
	wire [0:0] andOp_454_out;
	andOp #(.WIDTH(1)) andOp_454(.in0(andOp_454_in0), .in1(andOp_454_in1), .out(andOp_454_out));

	reg [0:0] notOp_455_in0;
	wire [0:0] notOp_455_out;
	notOp #(.WIDTH(1)) notOp_455(.in(notOp_455_in0), .out(notOp_455_out));

	reg [0:0] andOp_456_in0;
	reg [0:0] andOp_456_in1;
	wire [0:0] andOp_456_out;
	andOp #(.WIDTH(1)) andOp_456(.in0(andOp_456_in0), .in1(andOp_456_in1), .out(andOp_456_out));

	reg [0:0] andOp_457_in0;
	reg [0:0] andOp_457_in1;
	wire [0:0] andOp_457_out;
	andOp #(.WIDTH(1)) andOp_457(.in0(andOp_457_in0), .in1(andOp_457_in1), .out(andOp_457_out));

	reg [31:0] eq_458_in0;
	reg [31:0] eq_458_in1;
	wire [0:0] eq_458_out;
	eq #(.WIDTH(32)) eq_458(.in0(eq_458_in0), .in1(eq_458_in1), .out(eq_458_out));

	reg [0:0] andOp_459_in0;
	reg [0:0] andOp_459_in1;
	wire [0:0] andOp_459_out;
	andOp #(.WIDTH(1)) andOp_459(.in0(andOp_459_in0), .in1(andOp_459_in1), .out(andOp_459_out));

	reg [0:0] notOp_460_in0;
	wire [0:0] notOp_460_out;
	notOp #(.WIDTH(1)) notOp_460(.in(notOp_460_in0), .out(notOp_460_out));

	reg [0:0] andOp_461_in0;
	reg [0:0] andOp_461_in1;
	wire [0:0] andOp_461_out;
	andOp #(.WIDTH(1)) andOp_461(.in0(andOp_461_in0), .in1(andOp_461_in1), .out(andOp_461_out));

	reg [31:0] eq_462_in0;
	reg [31:0] eq_462_in1;
	wire [0:0] eq_462_out;
	eq #(.WIDTH(32)) eq_462(.in0(eq_462_in0), .in1(eq_462_in1), .out(eq_462_out));

	reg [0:0] andOp_463_in0;
	reg [0:0] andOp_463_in1;
	wire [0:0] andOp_463_out;
	andOp #(.WIDTH(1)) andOp_463(.in0(andOp_463_in0), .in1(andOp_463_in1), .out(andOp_463_out));

	reg [31:0] eq_464_in0;
	reg [31:0] eq_464_in1;
	wire [0:0] eq_464_out;
	eq #(.WIDTH(32)) eq_464(.in0(eq_464_in0), .in1(eq_464_in1), .out(eq_464_out));

	reg [0:0] andOp_465_in0;
	reg [0:0] andOp_465_in1;
	wire [0:0] andOp_465_out;
	andOp #(.WIDTH(1)) andOp_465(.in0(andOp_465_in0), .in1(andOp_465_in1), .out(andOp_465_out));

	reg [0:0] notOp_466_in0;
	wire [0:0] notOp_466_out;
	notOp #(.WIDTH(1)) notOp_466(.in(notOp_466_in0), .out(notOp_466_out));

	reg [0:0] andOp_467_in0;
	reg [0:0] andOp_467_in1;
	wire [0:0] andOp_467_out;
	andOp #(.WIDTH(1)) andOp_467(.in0(andOp_467_in0), .in1(andOp_467_in1), .out(andOp_467_out));

	reg [0:0] andOp_468_in0;
	reg [0:0] andOp_468_in1;
	wire [0:0] andOp_468_out;
	andOp #(.WIDTH(1)) andOp_468(.in0(andOp_468_in0), .in1(andOp_468_in1), .out(andOp_468_out));

	reg [31:0] eq_469_in0;
	reg [31:0] eq_469_in1;
	wire [0:0] eq_469_out;
	eq #(.WIDTH(32)) eq_469(.in0(eq_469_in0), .in1(eq_469_in1), .out(eq_469_out));

	reg [0:0] andOp_470_in0;
	reg [0:0] andOp_470_in1;
	wire [0:0] andOp_470_out;
	andOp #(.WIDTH(1)) andOp_470(.in0(andOp_470_in0), .in1(andOp_470_in1), .out(andOp_470_out));

	reg [0:0] notOp_471_in0;
	wire [0:0] notOp_471_out;
	notOp #(.WIDTH(1)) notOp_471(.in(notOp_471_in0), .out(notOp_471_out));

	reg [0:0] andOp_472_in0;
	reg [0:0] andOp_472_in1;
	wire [0:0] andOp_472_out;
	andOp #(.WIDTH(1)) andOp_472(.in0(andOp_472_in0), .in1(andOp_472_in1), .out(andOp_472_out));

	reg [31:0] eq_473_in0;
	reg [31:0] eq_473_in1;
	wire [0:0] eq_473_out;
	eq #(.WIDTH(32)) eq_473(.in0(eq_473_in0), .in1(eq_473_in1), .out(eq_473_out));

	reg [0:0] andOp_474_in0;
	reg [0:0] andOp_474_in1;
	wire [0:0] andOp_474_out;
	andOp #(.WIDTH(1)) andOp_474(.in0(andOp_474_in0), .in1(andOp_474_in1), .out(andOp_474_out));

	reg [0:0] notOp_475_in0;
	wire [0:0] notOp_475_out;
	notOp #(.WIDTH(1)) notOp_475(.in(notOp_475_in0), .out(notOp_475_out));

	reg [0:0] andOp_476_in0;
	reg [0:0] andOp_476_in1;
	wire [0:0] andOp_476_out;
	andOp #(.WIDTH(1)) andOp_476(.in0(andOp_476_in0), .in1(andOp_476_in1), .out(andOp_476_out));

	reg [0:0] andOp_477_in0;
	reg [0:0] andOp_477_in1;
	wire [0:0] andOp_477_out;
	andOp #(.WIDTH(1)) andOp_477(.in0(andOp_477_in0), .in1(andOp_477_in1), .out(andOp_477_out));

	reg [31:0] eq_478_in0;
	reg [31:0] eq_478_in1;
	wire [0:0] eq_478_out;
	eq #(.WIDTH(32)) eq_478(.in0(eq_478_in0), .in1(eq_478_in1), .out(eq_478_out));

	reg [0:0] andOp_479_in0;
	reg [0:0] andOp_479_in1;
	wire [0:0] andOp_479_out;
	andOp #(.WIDTH(1)) andOp_479(.in0(andOp_479_in0), .in1(andOp_479_in1), .out(andOp_479_out));

	reg [0:0] notOp_480_in0;
	wire [0:0] notOp_480_out;
	notOp #(.WIDTH(1)) notOp_480(.in(notOp_480_in0), .out(notOp_480_out));

	reg [0:0] andOp_481_in0;
	reg [0:0] andOp_481_in1;
	wire [0:0] andOp_481_out;
	andOp #(.WIDTH(1)) andOp_481(.in0(andOp_481_in0), .in1(andOp_481_in1), .out(andOp_481_out));

	reg [31:0] eq_482_in0;
	reg [31:0] eq_482_in1;
	wire [0:0] eq_482_out;
	eq #(.WIDTH(32)) eq_482(.in0(eq_482_in0), .in1(eq_482_in1), .out(eq_482_out));

	reg [0:0] andOp_483_in0;
	reg [0:0] andOp_483_in1;
	wire [0:0] andOp_483_out;
	andOp #(.WIDTH(1)) andOp_483(.in0(andOp_483_in0), .in1(andOp_483_in1), .out(andOp_483_out));

	reg [31:0] eq_484_in0;
	reg [31:0] eq_484_in1;
	wire [0:0] eq_484_out;
	eq #(.WIDTH(32)) eq_484(.in0(eq_484_in0), .in1(eq_484_in1), .out(eq_484_out));

	reg [0:0] andOp_485_in0;
	reg [0:0] andOp_485_in1;
	wire [0:0] andOp_485_out;
	andOp #(.WIDTH(1)) andOp_485(.in0(andOp_485_in0), .in1(andOp_485_in1), .out(andOp_485_out));

	reg [0:0] notOp_486_in0;
	wire [0:0] notOp_486_out;
	notOp #(.WIDTH(1)) notOp_486(.in(notOp_486_in0), .out(notOp_486_out));

	reg [0:0] andOp_487_in0;
	reg [0:0] andOp_487_in1;
	wire [0:0] andOp_487_out;
	andOp #(.WIDTH(1)) andOp_487(.in0(andOp_487_in0), .in1(andOp_487_in1), .out(andOp_487_out));

	reg [0:0] andOp_488_in0;
	reg [0:0] andOp_488_in1;
	wire [0:0] andOp_488_out;
	andOp #(.WIDTH(1)) andOp_488(.in0(andOp_488_in0), .in1(andOp_488_in1), .out(andOp_488_out));

	reg [31:0] eq_489_in0;
	reg [31:0] eq_489_in1;
	wire [0:0] eq_489_out;
	eq #(.WIDTH(32)) eq_489(.in0(eq_489_in0), .in1(eq_489_in1), .out(eq_489_out));

	reg [0:0] andOp_490_in0;
	reg [0:0] andOp_490_in1;
	wire [0:0] andOp_490_out;
	andOp #(.WIDTH(1)) andOp_490(.in0(andOp_490_in0), .in1(andOp_490_in1), .out(andOp_490_out));

	reg [0:0] notOp_491_in0;
	wire [0:0] notOp_491_out;
	notOp #(.WIDTH(1)) notOp_491(.in(notOp_491_in0), .out(notOp_491_out));

	reg [0:0] andOp_492_in0;
	reg [0:0] andOp_492_in1;
	wire [0:0] andOp_492_out;
	andOp #(.WIDTH(1)) andOp_492(.in0(andOp_492_in0), .in1(andOp_492_in1), .out(andOp_492_out));

	reg [0:0] notOp_493_in0;
	wire [0:0] notOp_493_out;
	notOp #(.WIDTH(1)) notOp_493(.in(notOp_493_in0), .out(notOp_493_out));

	reg [0:0] andOp_494_in0;
	reg [0:0] andOp_494_in1;
	wire [0:0] andOp_494_out;
	andOp #(.WIDTH(1)) andOp_494(.in0(andOp_494_in0), .in1(andOp_494_in1), .out(andOp_494_out));

	reg [0:0] andOp_495_in0;
	reg [0:0] andOp_495_in1;
	wire [0:0] andOp_495_out;
	andOp #(.WIDTH(1)) andOp_495(.in0(andOp_495_in0), .in1(andOp_495_in1), .out(andOp_495_out));

	reg [31:0] eq_496_in0;
	reg [31:0] eq_496_in1;
	wire [0:0] eq_496_out;
	eq #(.WIDTH(32)) eq_496(.in0(eq_496_in0), .in1(eq_496_in1), .out(eq_496_out));

	reg [0:0] andOp_497_in0;
	reg [0:0] andOp_497_in1;
	wire [0:0] andOp_497_out;
	andOp #(.WIDTH(1)) andOp_497(.in0(andOp_497_in0), .in1(andOp_497_in1), .out(andOp_497_out));

	reg [0:0] notOp_498_in0;
	wire [0:0] notOp_498_out;
	notOp #(.WIDTH(1)) notOp_498(.in(notOp_498_in0), .out(notOp_498_out));

	reg [0:0] andOp_499_in0;
	reg [0:0] andOp_499_in1;
	wire [0:0] andOp_499_out;
	andOp #(.WIDTH(1)) andOp_499(.in0(andOp_499_in0), .in1(andOp_499_in1), .out(andOp_499_out));

	reg [0:0] notOp_500_in0;
	wire [0:0] notOp_500_out;
	notOp #(.WIDTH(1)) notOp_500(.in(notOp_500_in0), .out(notOp_500_out));

	reg [0:0] andOp_501_in0;
	reg [0:0] andOp_501_in1;
	wire [0:0] andOp_501_out;
	andOp #(.WIDTH(1)) andOp_501(.in0(andOp_501_in0), .in1(andOp_501_in1), .out(andOp_501_out));

	reg [0:0] andOp_502_in0;
	reg [0:0] andOp_502_in1;
	wire [0:0] andOp_502_out;
	andOp #(.WIDTH(1)) andOp_502(.in0(andOp_502_in0), .in1(andOp_502_in1), .out(andOp_502_out));

	reg [31:0] eq_503_in0;
	reg [31:0] eq_503_in1;
	wire [0:0] eq_503_out;
	eq #(.WIDTH(32)) eq_503(.in0(eq_503_in0), .in1(eq_503_in1), .out(eq_503_out));

	reg [0:0] andOp_504_in0;
	reg [0:0] andOp_504_in1;
	wire [0:0] andOp_504_out;
	andOp #(.WIDTH(1)) andOp_504(.in0(andOp_504_in0), .in1(andOp_504_in1), .out(andOp_504_out));

	reg [0:0] notOp_505_in0;
	wire [0:0] notOp_505_out;
	notOp #(.WIDTH(1)) notOp_505(.in(notOp_505_in0), .out(notOp_505_out));

	reg [0:0] andOp_506_in0;
	reg [0:0] andOp_506_in1;
	wire [0:0] andOp_506_out;
	andOp #(.WIDTH(1)) andOp_506(.in0(andOp_506_in0), .in1(andOp_506_in1), .out(andOp_506_out));

	reg [0:0] notOp_507_in0;
	wire [0:0] notOp_507_out;
	notOp #(.WIDTH(1)) notOp_507(.in(notOp_507_in0), .out(notOp_507_out));

	reg [0:0] andOp_508_in0;
	reg [0:0] andOp_508_in1;
	wire [0:0] andOp_508_out;
	andOp #(.WIDTH(1)) andOp_508(.in0(andOp_508_in0), .in1(andOp_508_in1), .out(andOp_508_out));

	reg [0:0] andOp_509_in0;
	reg [0:0] andOp_509_in1;
	wire [0:0] andOp_509_out;
	andOp #(.WIDTH(1)) andOp_509(.in0(andOp_509_in0), .in1(andOp_509_in1), .out(andOp_509_out));

	reg [31:0] eq_510_in0;
	reg [31:0] eq_510_in1;
	wire [0:0] eq_510_out;
	eq #(.WIDTH(32)) eq_510(.in0(eq_510_in0), .in1(eq_510_in1), .out(eq_510_out));

	reg [0:0] andOp_511_in0;
	reg [0:0] andOp_511_in1;
	wire [0:0] andOp_511_out;
	andOp #(.WIDTH(1)) andOp_511(.in0(andOp_511_in0), .in1(andOp_511_in1), .out(andOp_511_out));

	reg [0:0] notOp_512_in0;
	wire [0:0] notOp_512_out;
	notOp #(.WIDTH(1)) notOp_512(.in(notOp_512_in0), .out(notOp_512_out));

	reg [0:0] andOp_513_in0;
	reg [0:0] andOp_513_in1;
	wire [0:0] andOp_513_out;
	andOp #(.WIDTH(1)) andOp_513(.in0(andOp_513_in0), .in1(andOp_513_in1), .out(andOp_513_out));

	reg [0:0] notOp_514_in0;
	wire [0:0] notOp_514_out;
	notOp #(.WIDTH(1)) notOp_514(.in(notOp_514_in0), .out(notOp_514_out));

	reg [0:0] andOp_515_in0;
	reg [0:0] andOp_515_in1;
	wire [0:0] andOp_515_out;
	andOp #(.WIDTH(1)) andOp_515(.in0(andOp_515_in0), .in1(andOp_515_in1), .out(andOp_515_out));

	reg [0:0] andOp_516_in0;
	reg [0:0] andOp_516_in1;
	wire [0:0] andOp_516_out;
	andOp #(.WIDTH(1)) andOp_516(.in0(andOp_516_in0), .in1(andOp_516_in1), .out(andOp_516_out));

	reg [31:0] eq_517_in0;
	reg [31:0] eq_517_in1;
	wire [0:0] eq_517_out;
	eq #(.WIDTH(32)) eq_517(.in0(eq_517_in0), .in1(eq_517_in1), .out(eq_517_out));

	reg [0:0] andOp_518_in0;
	reg [0:0] andOp_518_in1;
	wire [0:0] andOp_518_out;
	andOp #(.WIDTH(1)) andOp_518(.in0(andOp_518_in0), .in1(andOp_518_in1), .out(andOp_518_out));

	reg [0:0] notOp_519_in0;
	wire [0:0] notOp_519_out;
	notOp #(.WIDTH(1)) notOp_519(.in(notOp_519_in0), .out(notOp_519_out));

	reg [0:0] andOp_520_in0;
	reg [0:0] andOp_520_in1;
	wire [0:0] andOp_520_out;
	andOp #(.WIDTH(1)) andOp_520(.in0(andOp_520_in0), .in1(andOp_520_in1), .out(andOp_520_out));

	reg [31:0] eq_521_in0;
	reg [31:0] eq_521_in1;
	wire [0:0] eq_521_out;
	eq #(.WIDTH(32)) eq_521(.in0(eq_521_in0), .in1(eq_521_in1), .out(eq_521_out));

	reg [0:0] andOp_522_in0;
	reg [0:0] andOp_522_in1;
	wire [0:0] andOp_522_out;
	andOp #(.WIDTH(1)) andOp_522(.in0(andOp_522_in0), .in1(andOp_522_in1), .out(andOp_522_out));

	reg [0:0] notOp_523_in0;
	wire [0:0] notOp_523_out;
	notOp #(.WIDTH(1)) notOp_523(.in(notOp_523_in0), .out(notOp_523_out));

	reg [0:0] andOp_524_in0;
	reg [0:0] andOp_524_in1;
	wire [0:0] andOp_524_out;
	andOp #(.WIDTH(1)) andOp_524(.in0(andOp_524_in0), .in1(andOp_524_in1), .out(andOp_524_out));

	reg [0:0] andOp_525_in0;
	reg [0:0] andOp_525_in1;
	wire [0:0] andOp_525_out;
	andOp #(.WIDTH(1)) andOp_525(.in0(andOp_525_in0), .in1(andOp_525_in1), .out(andOp_525_out));

	reg [31:0] eq_526_in0;
	reg [31:0] eq_526_in1;
	wire [0:0] eq_526_out;
	eq #(.WIDTH(32)) eq_526(.in0(eq_526_in0), .in1(eq_526_in1), .out(eq_526_out));

	reg [0:0] andOp_527_in0;
	reg [0:0] andOp_527_in1;
	wire [0:0] andOp_527_out;
	andOp #(.WIDTH(1)) andOp_527(.in0(andOp_527_in0), .in1(andOp_527_in1), .out(andOp_527_out));

	reg [0:0] notOp_528_in0;
	wire [0:0] notOp_528_out;
	notOp #(.WIDTH(1)) notOp_528(.in(notOp_528_in0), .out(notOp_528_out));

	reg [0:0] andOp_529_in0;
	reg [0:0] andOp_529_in1;
	wire [0:0] andOp_529_out;
	andOp #(.WIDTH(1)) andOp_529(.in0(andOp_529_in0), .in1(andOp_529_in1), .out(andOp_529_out));

	reg [31:0] eq_530_in0;
	reg [31:0] eq_530_in1;
	wire [0:0] eq_530_out;
	eq #(.WIDTH(32)) eq_530(.in0(eq_530_in0), .in1(eq_530_in1), .out(eq_530_out));

	reg [0:0] andOp_531_in0;
	reg [0:0] andOp_531_in1;
	wire [0:0] andOp_531_out;
	andOp #(.WIDTH(1)) andOp_531(.in0(andOp_531_in0), .in1(andOp_531_in1), .out(andOp_531_out));

	reg [31:0] eq_532_in0;
	reg [31:0] eq_532_in1;
	wire [0:0] eq_532_out;
	eq #(.WIDTH(32)) eq_532(.in0(eq_532_in0), .in1(eq_532_in1), .out(eq_532_out));

	reg [0:0] andOp_533_in0;
	reg [0:0] andOp_533_in1;
	wire [0:0] andOp_533_out;
	andOp #(.WIDTH(1)) andOp_533(.in0(andOp_533_in0), .in1(andOp_533_in1), .out(andOp_533_out));

	reg [0:0] notOp_534_in0;
	wire [0:0] notOp_534_out;
	notOp #(.WIDTH(1)) notOp_534(.in(notOp_534_in0), .out(notOp_534_out));

	reg [0:0] andOp_535_in0;
	reg [0:0] andOp_535_in1;
	wire [0:0] andOp_535_out;
	andOp #(.WIDTH(1)) andOp_535(.in0(andOp_535_in0), .in1(andOp_535_in1), .out(andOp_535_out));

	reg [0:0] andOp_536_in0;
	reg [0:0] andOp_536_in1;
	wire [0:0] andOp_536_out;
	andOp #(.WIDTH(1)) andOp_536(.in0(andOp_536_in0), .in1(andOp_536_in1), .out(andOp_536_out));

	reg [31:0] eq_537_in0;
	reg [31:0] eq_537_in1;
	wire [0:0] eq_537_out;
	eq #(.WIDTH(32)) eq_537(.in0(eq_537_in0), .in1(eq_537_in1), .out(eq_537_out));

	reg [0:0] andOp_538_in0;
	reg [0:0] andOp_538_in1;
	wire [0:0] andOp_538_out;
	andOp #(.WIDTH(1)) andOp_538(.in0(andOp_538_in0), .in1(andOp_538_in1), .out(andOp_538_out));

	reg [0:0] notOp_539_in0;
	wire [0:0] notOp_539_out;
	notOp #(.WIDTH(1)) notOp_539(.in(notOp_539_in0), .out(notOp_539_out));

	reg [0:0] andOp_540_in0;
	reg [0:0] andOp_540_in1;
	wire [0:0] andOp_540_out;
	andOp #(.WIDTH(1)) andOp_540(.in0(andOp_540_in0), .in1(andOp_540_in1), .out(andOp_540_out));

	reg [31:0] eq_541_in0;
	reg [31:0] eq_541_in1;
	wire [0:0] eq_541_out;
	eq #(.WIDTH(32)) eq_541(.in0(eq_541_in0), .in1(eq_541_in1), .out(eq_541_out));

	reg [0:0] andOp_542_in0;
	reg [0:0] andOp_542_in1;
	wire [0:0] andOp_542_out;
	andOp #(.WIDTH(1)) andOp_542(.in0(andOp_542_in0), .in1(andOp_542_in1), .out(andOp_542_out));

	reg [31:0] eq_543_in0;
	reg [31:0] eq_543_in1;
	wire [0:0] eq_543_out;
	eq #(.WIDTH(32)) eq_543(.in0(eq_543_in0), .in1(eq_543_in1), .out(eq_543_out));

	reg [0:0] andOp_544_in0;
	reg [0:0] andOp_544_in1;
	wire [0:0] andOp_544_out;
	andOp #(.WIDTH(1)) andOp_544(.in0(andOp_544_in0), .in1(andOp_544_in1), .out(andOp_544_out));

	reg [0:0] notOp_545_in0;
	wire [0:0] notOp_545_out;
	notOp #(.WIDTH(1)) notOp_545(.in(notOp_545_in0), .out(notOp_545_out));

	reg [0:0] andOp_546_in0;
	reg [0:0] andOp_546_in1;
	wire [0:0] andOp_546_out;
	andOp #(.WIDTH(1)) andOp_546(.in0(andOp_546_in0), .in1(andOp_546_in1), .out(andOp_546_out));

	reg [0:0] andOp_547_in0;
	reg [0:0] andOp_547_in1;
	wire [0:0] andOp_547_out;
	andOp #(.WIDTH(1)) andOp_547(.in0(andOp_547_in0), .in1(andOp_547_in1), .out(andOp_547_out));

	reg [31:0] eq_548_in0;
	reg [31:0] eq_548_in1;
	wire [0:0] eq_548_out;
	eq #(.WIDTH(32)) eq_548(.in0(eq_548_in0), .in1(eq_548_in1), .out(eq_548_out));

	reg [0:0] andOp_549_in0;
	reg [0:0] andOp_549_in1;
	wire [0:0] andOp_549_out;
	andOp #(.WIDTH(1)) andOp_549(.in0(andOp_549_in0), .in1(andOp_549_in1), .out(andOp_549_out));

	reg [0:0] notOp_550_in0;
	wire [0:0] notOp_550_out;
	notOp #(.WIDTH(1)) notOp_550(.in(notOp_550_in0), .out(notOp_550_out));

	reg [0:0] andOp_551_in0;
	reg [0:0] andOp_551_in1;
	wire [0:0] andOp_551_out;
	andOp #(.WIDTH(1)) andOp_551(.in0(andOp_551_in0), .in1(andOp_551_in1), .out(andOp_551_out));

	reg [31:0] eq_552_in0;
	reg [31:0] eq_552_in1;
	wire [0:0] eq_552_out;
	eq #(.WIDTH(32)) eq_552(.in0(eq_552_in0), .in1(eq_552_in1), .out(eq_552_out));

	reg [0:0] andOp_553_in0;
	reg [0:0] andOp_553_in1;
	wire [0:0] andOp_553_out;
	andOp #(.WIDTH(1)) andOp_553(.in0(andOp_553_in0), .in1(andOp_553_in1), .out(andOp_553_out));

	reg [0:0] notOp_554_in0;
	wire [0:0] notOp_554_out;
	notOp #(.WIDTH(1)) notOp_554(.in(notOp_554_in0), .out(notOp_554_out));

	reg [0:0] andOp_555_in0;
	reg [0:0] andOp_555_in1;
	wire [0:0] andOp_555_out;
	andOp #(.WIDTH(1)) andOp_555(.in0(andOp_555_in0), .in1(andOp_555_in1), .out(andOp_555_out));

	reg [0:0] andOp_556_in0;
	reg [0:0] andOp_556_in1;
	wire [0:0] andOp_556_out;
	andOp #(.WIDTH(1)) andOp_556(.in0(andOp_556_in0), .in1(andOp_556_in1), .out(andOp_556_out));

	reg [31:0] eq_557_in0;
	reg [31:0] eq_557_in1;
	wire [0:0] eq_557_out;
	eq #(.WIDTH(32)) eq_557(.in0(eq_557_in0), .in1(eq_557_in1), .out(eq_557_out));

	reg [0:0] andOp_558_in0;
	reg [0:0] andOp_558_in1;
	wire [0:0] andOp_558_out;
	andOp #(.WIDTH(1)) andOp_558(.in0(andOp_558_in0), .in1(andOp_558_in1), .out(andOp_558_out));

	reg [0:0] notOp_559_in0;
	wire [0:0] notOp_559_out;
	notOp #(.WIDTH(1)) notOp_559(.in(notOp_559_in0), .out(notOp_559_out));

	reg [0:0] andOp_560_in0;
	reg [0:0] andOp_560_in1;
	wire [0:0] andOp_560_out;
	andOp #(.WIDTH(1)) andOp_560(.in0(andOp_560_in0), .in1(andOp_560_in1), .out(andOp_560_out));

	reg [31:0] eq_561_in0;
	reg [31:0] eq_561_in1;
	wire [0:0] eq_561_out;
	eq #(.WIDTH(32)) eq_561(.in0(eq_561_in0), .in1(eq_561_in1), .out(eq_561_out));

	reg [0:0] andOp_562_in0;
	reg [0:0] andOp_562_in1;
	wire [0:0] andOp_562_out;
	andOp #(.WIDTH(1)) andOp_562(.in0(andOp_562_in0), .in1(andOp_562_in1), .out(andOp_562_out));

	reg [31:0] eq_563_in0;
	reg [31:0] eq_563_in1;
	wire [0:0] eq_563_out;
	eq #(.WIDTH(32)) eq_563(.in0(eq_563_in0), .in1(eq_563_in1), .out(eq_563_out));

	reg [0:0] andOp_564_in0;
	reg [0:0] andOp_564_in1;
	wire [0:0] andOp_564_out;
	andOp #(.WIDTH(1)) andOp_564(.in0(andOp_564_in0), .in1(andOp_564_in1), .out(andOp_564_out));

	reg [0:0] notOp_565_in0;
	wire [0:0] notOp_565_out;
	notOp #(.WIDTH(1)) notOp_565(.in(notOp_565_in0), .out(notOp_565_out));

	reg [0:0] andOp_566_in0;
	reg [0:0] andOp_566_in1;
	wire [0:0] andOp_566_out;
	andOp #(.WIDTH(1)) andOp_566(.in0(andOp_566_in0), .in1(andOp_566_in1), .out(andOp_566_out));

	reg [0:0] andOp_567_in0;
	reg [0:0] andOp_567_in1;
	wire [0:0] andOp_567_out;
	andOp #(.WIDTH(1)) andOp_567(.in0(andOp_567_in0), .in1(andOp_567_in1), .out(andOp_567_out));

	reg [31:0] eq_568_in0;
	reg [31:0] eq_568_in1;
	wire [0:0] eq_568_out;
	eq #(.WIDTH(32)) eq_568(.in0(eq_568_in0), .in1(eq_568_in1), .out(eq_568_out));

	reg [0:0] andOp_569_in0;
	reg [0:0] andOp_569_in1;
	wire [0:0] andOp_569_out;
	andOp #(.WIDTH(1)) andOp_569(.in0(andOp_569_in0), .in1(andOp_569_in1), .out(andOp_569_out));

	reg [0:0] notOp_570_in0;
	wire [0:0] notOp_570_out;
	notOp #(.WIDTH(1)) notOp_570(.in(notOp_570_in0), .out(notOp_570_out));

	reg [0:0] andOp_571_in0;
	reg [0:0] andOp_571_in1;
	wire [0:0] andOp_571_out;
	andOp #(.WIDTH(1)) andOp_571(.in0(andOp_571_in0), .in1(andOp_571_in1), .out(andOp_571_out));

	reg [31:0] eq_572_in0;
	reg [31:0] eq_572_in1;
	wire [0:0] eq_572_out;
	eq #(.WIDTH(32)) eq_572(.in0(eq_572_in0), .in1(eq_572_in1), .out(eq_572_out));

	reg [0:0] andOp_573_in0;
	reg [0:0] andOp_573_in1;
	wire [0:0] andOp_573_out;
	andOp #(.WIDTH(1)) andOp_573(.in0(andOp_573_in0), .in1(andOp_573_in1), .out(andOp_573_out));

	reg [0:0] notOp_574_in0;
	wire [0:0] notOp_574_out;
	notOp #(.WIDTH(1)) notOp_574(.in(notOp_574_in0), .out(notOp_574_out));

	reg [0:0] andOp_575_in0;
	reg [0:0] andOp_575_in1;
	wire [0:0] andOp_575_out;
	andOp #(.WIDTH(1)) andOp_575(.in0(andOp_575_in0), .in1(andOp_575_in1), .out(andOp_575_out));

	reg [0:0] andOp_576_in0;
	reg [0:0] andOp_576_in1;
	wire [0:0] andOp_576_out;
	andOp #(.WIDTH(1)) andOp_576(.in0(andOp_576_in0), .in1(andOp_576_in1), .out(andOp_576_out));

	reg [31:0] eq_577_in0;
	reg [31:0] eq_577_in1;
	wire [0:0] eq_577_out;
	eq #(.WIDTH(32)) eq_577(.in0(eq_577_in0), .in1(eq_577_in1), .out(eq_577_out));

	reg [0:0] andOp_578_in0;
	reg [0:0] andOp_578_in1;
	wire [0:0] andOp_578_out;
	andOp #(.WIDTH(1)) andOp_578(.in0(andOp_578_in0), .in1(andOp_578_in1), .out(andOp_578_out));

	reg [0:0] notOp_579_in0;
	wire [0:0] notOp_579_out;
	notOp #(.WIDTH(1)) notOp_579(.in(notOp_579_in0), .out(notOp_579_out));

	reg [0:0] andOp_580_in0;
	reg [0:0] andOp_580_in1;
	wire [0:0] andOp_580_out;
	andOp #(.WIDTH(1)) andOp_580(.in0(andOp_580_in0), .in1(andOp_580_in1), .out(andOp_580_out));

	reg [31:0] eq_581_in0;
	reg [31:0] eq_581_in1;
	wire [0:0] eq_581_out;
	eq #(.WIDTH(32)) eq_581(.in0(eq_581_in0), .in1(eq_581_in1), .out(eq_581_out));

	reg [0:0] andOp_582_in0;
	reg [0:0] andOp_582_in1;
	wire [0:0] andOp_582_out;
	andOp #(.WIDTH(1)) andOp_582(.in0(andOp_582_in0), .in1(andOp_582_in1), .out(andOp_582_out));

	reg [0:0] notOp_583_in0;
	wire [0:0] notOp_583_out;
	notOp #(.WIDTH(1)) notOp_583(.in(notOp_583_in0), .out(notOp_583_out));

	reg [0:0] andOp_584_in0;
	reg [0:0] andOp_584_in1;
	wire [0:0] andOp_584_out;
	andOp #(.WIDTH(1)) andOp_584(.in0(andOp_584_in0), .in1(andOp_584_in1), .out(andOp_584_out));

	reg [0:0] andOp_585_in0;
	reg [0:0] andOp_585_in1;
	wire [0:0] andOp_585_out;
	andOp #(.WIDTH(1)) andOp_585(.in0(andOp_585_in0), .in1(andOp_585_in1), .out(andOp_585_out));

	reg [31:0] eq_586_in0;
	reg [31:0] eq_586_in1;
	wire [0:0] eq_586_out;
	eq #(.WIDTH(32)) eq_586(.in0(eq_586_in0), .in1(eq_586_in1), .out(eq_586_out));

	reg [0:0] andOp_587_in0;
	reg [0:0] andOp_587_in1;
	wire [0:0] andOp_587_out;
	andOp #(.WIDTH(1)) andOp_587(.in0(andOp_587_in0), .in1(andOp_587_in1), .out(andOp_587_out));

	reg [0:0] notOp_588_in0;
	wire [0:0] notOp_588_out;
	notOp #(.WIDTH(1)) notOp_588(.in(notOp_588_in0), .out(notOp_588_out));

	reg [0:0] andOp_589_in0;
	reg [0:0] andOp_589_in1;
	wire [0:0] andOp_589_out;
	andOp #(.WIDTH(1)) andOp_589(.in0(andOp_589_in0), .in1(andOp_589_in1), .out(andOp_589_out));

	reg [31:0] eq_590_in0;
	reg [31:0] eq_590_in1;
	wire [0:0] eq_590_out;
	eq #(.WIDTH(32)) eq_590(.in0(eq_590_in0), .in1(eq_590_in1), .out(eq_590_out));

	reg [0:0] andOp_591_in0;
	reg [0:0] andOp_591_in1;
	wire [0:0] andOp_591_out;
	andOp #(.WIDTH(1)) andOp_591(.in0(andOp_591_in0), .in1(andOp_591_in1), .out(andOp_591_out));

	reg [0:0] notOp_592_in0;
	wire [0:0] notOp_592_out;
	notOp #(.WIDTH(1)) notOp_592(.in(notOp_592_in0), .out(notOp_592_out));

	reg [0:0] andOp_593_in0;
	reg [0:0] andOp_593_in1;
	wire [0:0] andOp_593_out;
	andOp #(.WIDTH(1)) andOp_593(.in0(andOp_593_in0), .in1(andOp_593_in1), .out(andOp_593_out));

	reg [0:0] andOp_594_in0;
	reg [0:0] andOp_594_in1;
	wire [0:0] andOp_594_out;
	andOp #(.WIDTH(1)) andOp_594(.in0(andOp_594_in0), .in1(andOp_594_in1), .out(andOp_594_out));

	reg [31:0] eq_595_in0;
	reg [31:0] eq_595_in1;
	wire [0:0] eq_595_out;
	eq #(.WIDTH(32)) eq_595(.in0(eq_595_in0), .in1(eq_595_in1), .out(eq_595_out));

	reg [0:0] andOp_596_in0;
	reg [0:0] andOp_596_in1;
	wire [0:0] andOp_596_out;
	andOp #(.WIDTH(1)) andOp_596(.in0(andOp_596_in0), .in1(andOp_596_in1), .out(andOp_596_out));

	reg [0:0] notOp_597_in0;
	wire [0:0] notOp_597_out;
	notOp #(.WIDTH(1)) notOp_597(.in(notOp_597_in0), .out(notOp_597_out));

	reg [0:0] andOp_598_in0;
	reg [0:0] andOp_598_in1;
	wire [0:0] andOp_598_out;
	andOp #(.WIDTH(1)) andOp_598(.in0(andOp_598_in0), .in1(andOp_598_in1), .out(andOp_598_out));

	reg [31:0] eq_599_in0;
	reg [31:0] eq_599_in1;
	wire [0:0] eq_599_out;
	eq #(.WIDTH(32)) eq_599(.in0(eq_599_in0), .in1(eq_599_in1), .out(eq_599_out));

	reg [0:0] andOp_600_in0;
	reg [0:0] andOp_600_in1;
	wire [0:0] andOp_600_out;
	andOp #(.WIDTH(1)) andOp_600(.in0(andOp_600_in0), .in1(andOp_600_in1), .out(andOp_600_out));

	reg [0:0] notOp_601_in0;
	wire [0:0] notOp_601_out;
	notOp #(.WIDTH(1)) notOp_601(.in(notOp_601_in0), .out(notOp_601_out));

	reg [0:0] andOp_602_in0;
	reg [0:0] andOp_602_in1;
	wire [0:0] andOp_602_out;
	andOp #(.WIDTH(1)) andOp_602(.in0(andOp_602_in0), .in1(andOp_602_in1), .out(andOp_602_out));

	reg [0:0] andOp_603_in0;
	reg [0:0] andOp_603_in1;
	wire [0:0] andOp_603_out;
	andOp #(.WIDTH(1)) andOp_603(.in0(andOp_603_in0), .in1(andOp_603_in1), .out(andOp_603_out));

	reg [31:0] eq_604_in0;
	reg [31:0] eq_604_in1;
	wire [0:0] eq_604_out;
	eq #(.WIDTH(32)) eq_604(.in0(eq_604_in0), .in1(eq_604_in1), .out(eq_604_out));

	reg [0:0] andOp_605_in0;
	reg [0:0] andOp_605_in1;
	wire [0:0] andOp_605_out;
	andOp #(.WIDTH(1)) andOp_605(.in0(andOp_605_in0), .in1(andOp_605_in1), .out(andOp_605_out));

	reg [0:0] notOp_606_in0;
	wire [0:0] notOp_606_out;
	notOp #(.WIDTH(1)) notOp_606(.in(notOp_606_in0), .out(notOp_606_out));

	reg [0:0] andOp_607_in0;
	reg [0:0] andOp_607_in1;
	wire [0:0] andOp_607_out;
	andOp #(.WIDTH(1)) andOp_607(.in0(andOp_607_in0), .in1(andOp_607_in1), .out(andOp_607_out));

	reg [0:0] notOp_608_in0;
	wire [0:0] notOp_608_out;
	notOp #(.WIDTH(1)) notOp_608(.in(notOp_608_in0), .out(notOp_608_out));

	reg [0:0] andOp_609_in0;
	reg [0:0] andOp_609_in1;
	wire [0:0] andOp_609_out;
	andOp #(.WIDTH(1)) andOp_609(.in0(andOp_609_in0), .in1(andOp_609_in1), .out(andOp_609_out));

	reg [0:0] andOp_610_in0;
	reg [0:0] andOp_610_in1;
	wire [0:0] andOp_610_out;
	andOp #(.WIDTH(1)) andOp_610(.in0(andOp_610_in0), .in1(andOp_610_in1), .out(andOp_610_out));

	reg [31:0] eq_611_in0;
	reg [31:0] eq_611_in1;
	wire [0:0] eq_611_out;
	eq #(.WIDTH(32)) eq_611(.in0(eq_611_in0), .in1(eq_611_in1), .out(eq_611_out));

	reg [0:0] andOp_612_in0;
	reg [0:0] andOp_612_in1;
	wire [0:0] andOp_612_out;
	andOp #(.WIDTH(1)) andOp_612(.in0(andOp_612_in0), .in1(andOp_612_in1), .out(andOp_612_out));

	reg [0:0] notOp_613_in0;
	wire [0:0] notOp_613_out;
	notOp #(.WIDTH(1)) notOp_613(.in(notOp_613_in0), .out(notOp_613_out));

	reg [0:0] andOp_614_in0;
	reg [0:0] andOp_614_in1;
	wire [0:0] andOp_614_out;
	andOp #(.WIDTH(1)) andOp_614(.in0(andOp_614_in0), .in1(andOp_614_in1), .out(andOp_614_out));

	reg [31:0] eq_615_in0;
	reg [31:0] eq_615_in1;
	wire [0:0] eq_615_out;
	eq #(.WIDTH(32)) eq_615(.in0(eq_615_in0), .in1(eq_615_in1), .out(eq_615_out));

	reg [0:0] andOp_616_in0;
	reg [0:0] andOp_616_in1;
	wire [0:0] andOp_616_out;
	andOp #(.WIDTH(1)) andOp_616(.in0(andOp_616_in0), .in1(andOp_616_in1), .out(andOp_616_out));

	// End Functional Units

	reg [31:0] add_tmp_5;
	reg [31:0] call_tmp_2;
	reg [0:0] data_store_0_0;
	reg [31:0] data_store_0_1;
	reg [31:0] data_store_0_2;
	reg [31:0] data_store_0_3;
	reg [31:0] data_store_0_4;
	reg [31:0] data_store_0_5;
	reg [0:0] data_store_0_6;
	reg [31:0] data_store_0_7;
	reg [0:0] data_store_0_8;
	reg [31:0] data_store_1_10;
	reg [31:0] data_store_1_11;
	reg [31:0] data_store_1_12;
	reg [31:0] data_store_1_13;
	reg [31:0] data_store_1_14;
	reg [0:0] data_store_1_15;
	reg [31:0] data_store_1_16;
	reg [0:0] data_store_1_17;
	reg [0:0] data_store_1_9;
	reg [0:0] data_store_2_18;
	reg [31:0] data_store_2_19;
	reg [31:0] data_store_2_20;
	reg [31:0] data_store_2_21;
	reg [31:0] data_store_2_22;
	reg [31:0] data_store_2_23;
	reg [0:0] data_store_2_24;
	reg [31:0] data_store_2_25;
	reg [0:0] data_store_2_26;
	reg [0:0] data_store_3_27;
	reg [31:0] data_store_3_28;
	reg [31:0] data_store_3_29;
	reg [31:0] data_store_3_30;
	reg [31:0] data_store_3_31;
	reg [31:0] data_store_3_32;
	reg [0:0] data_store_3_33;
	reg [31:0] data_store_3_34;
	reg [0:0] data_store_3_35;
	reg [0:0] data_store_4_36;
	reg [31:0] data_store_4_37;
	reg [31:0] data_store_4_38;
	reg [31:0] data_store_4_39;
	reg [31:0] data_store_4_40;
	reg [31:0] data_store_4_41;
	reg [0:0] data_store_4_42;
	reg [31:0] data_store_4_43;
	reg [0:0] data_store_4_44;
	reg [31:0] global_state;
	reg [0:0] icmp_tmp_6;
	reg [31:0] phi_tmp_1;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;

	// controller for add_add_13.add_in0_add_13
	// controller for add_add_13.add_in1_add_13
	// Insensitive connections
	always @(*) begin
		add_in0_add_13 = valid ? rdata_ram_0 : rdata_ram_0;
		add_in1_add_13 = valid ? tmp_output_165_out_data : tmp_output_165_out_data;
	end
	// controller for add_add_15.add_in0_add_15
	// controller for add_add_15.add_in1_add_15
	// Insensitive connections
	always @(*) begin
		add_in0_add_15 = valid ? phi_tmp_1 : phi_tmp_1;
		add_in1_add_15 = valid ? 32'd1 : 32'd1;
	end
	// controller for andOp_122.andOp_122_in0
	// controller for andOp_122.andOp_122_in1
	// Insensitive connections
	always @(*) begin
		andOp_122_in0 = valid ? notOp_121_out : notOp_121_out;
		andOp_122_in1 = valid ? andOp_55_out : andOp_55_out;
	end
	// controller for andOp_126.andOp_126_in0
	// controller for andOp_126.andOp_126_in1
	// Insensitive connections
	always @(*) begin
		andOp_126_in0 = valid ? notOp_125_out : notOp_125_out;
		andOp_126_in1 = valid ? andOp_46_out : andOp_46_out;
	end
	// controller for andOp_129.andOp_129_in0
	// controller for andOp_129.andOp_129_in1
	// Insensitive connections
	always @(*) begin
		andOp_129_in0 = valid ? notOp_128_out : notOp_128_out;
		andOp_129_in1 = valid ? andOp_49_out : andOp_49_out;
	end
	// controller for andOp_133.andOp_133_in0
	// controller for andOp_133.andOp_133_in1
	// Insensitive connections
	always @(*) begin
		andOp_133_in0 = valid ? notOp_132_out : notOp_132_out;
		andOp_133_in1 = valid ? andOp_64_out : andOp_64_out;
	end
	// controller for andOp_137.andOp_137_in0
	// controller for andOp_137.andOp_137_in1
	// Insensitive connections
	always @(*) begin
		andOp_137_in0 = valid ? notOp_136_out : notOp_136_out;
		andOp_137_in1 = valid ? andOp_94_out : andOp_94_out;
	end
	// controller for andOp_140.andOp_140_in0
	// controller for andOp_140.andOp_140_in1
	// Insensitive connections
	always @(*) begin
		andOp_140_in0 = valid ? notOp_139_out : notOp_139_out;
		andOp_140_in1 = valid ? andOp_76_out : andOp_76_out;
	end
	// controller for andOp_143.andOp_143_in0
	// controller for andOp_143.andOp_143_in1
	// Insensitive connections
	always @(*) begin
		andOp_143_in0 = valid ? notOp_142_out : notOp_142_out;
		andOp_143_in1 = valid ? andOp_81_out : andOp_81_out;
	end
	// controller for andOp_147.andOp_147_in0
	// controller for andOp_147.andOp_147_in1
	// Insensitive connections
	always @(*) begin
		andOp_147_in0 = valid ? notOp_146_out : notOp_146_out;
		andOp_147_in1 = valid ? andOp_85_out : andOp_85_out;
	end
	// controller for andOp_150.andOp_150_in0
	// controller for andOp_150.andOp_150_in1
	// Insensitive connections
	always @(*) begin
		andOp_150_in0 = valid ? notOp_149_out : notOp_149_out;
		andOp_150_in1 = valid ? andOp_69_out : andOp_69_out;
	end
	// controller for andOp_151.andOp_151_in0
	// controller for andOp_151.andOp_151_in1
	// Insensitive connections
	always @(*) begin
		andOp_151_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_151_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_152.andOp_152_in0
	// controller for andOp_152.andOp_152_in1
	// Insensitive connections
	always @(*) begin
		andOp_152_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_152_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_153.andOp_153_in0
	// controller for andOp_153.andOp_153_in1
	// Insensitive connections
	always @(*) begin
		andOp_153_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_153_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_154.andOp_154_in0
	// controller for andOp_154.andOp_154_in1
	// Insensitive connections
	always @(*) begin
		andOp_154_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_154_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_155.andOp_155_in0
	// controller for andOp_155.andOp_155_in1
	// Insensitive connections
	always @(*) begin
		andOp_155_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_155_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_156.andOp_156_in0
	// controller for andOp_156.andOp_156_in1
	// Insensitive connections
	always @(*) begin
		andOp_156_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_156_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_157.andOp_157_in0
	// controller for andOp_157.andOp_157_in1
	// Insensitive connections
	always @(*) begin
		andOp_157_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_157_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_158.andOp_158_in0
	// controller for andOp_158.andOp_158_in1
	// Insensitive connections
	always @(*) begin
		andOp_158_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
		andOp_158_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_159.andOp_159_in0
	// controller for andOp_159.andOp_159_in1
	// Insensitive connections
	always @(*) begin
		andOp_159_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_159_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_160.andOp_160_in0
	// controller for andOp_160.andOp_160_in1
	// Insensitive connections
	always @(*) begin
		andOp_160_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_160_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_161.andOp_161_in0
	// controller for andOp_161.andOp_161_in1
	// Insensitive connections
	always @(*) begin
		andOp_161_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_161_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_164.andOp_164_in0
	// controller for andOp_164.andOp_164_in1
	// Insensitive connections
	always @(*) begin
		andOp_164_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_164_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_167.andOp_167_in0
	// controller for andOp_167.andOp_167_in1
	// Insensitive connections
	always @(*) begin
		andOp_167_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_167_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_168.andOp_168_in0
	// controller for andOp_168.andOp_168_in1
	// Insensitive connections
	always @(*) begin
		andOp_168_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_168_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_169.andOp_169_in0
	// controller for andOp_169.andOp_169_in1
	// Insensitive connections
	always @(*) begin
		andOp_169_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_169_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_170.andOp_170_in0
	// controller for andOp_170.andOp_170_in1
	// Insensitive connections
	always @(*) begin
		andOp_170_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_170_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_171.andOp_171_in0
	// controller for andOp_171.andOp_171_in1
	// Insensitive connections
	always @(*) begin
		andOp_171_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_171_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_172.andOp_172_in0
	// controller for andOp_172.andOp_172_in1
	// Insensitive connections
	always @(*) begin
		andOp_172_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_172_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_173.andOp_173_in0
	// controller for andOp_173.andOp_173_in1
	// Insensitive connections
	always @(*) begin
		andOp_173_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
		andOp_173_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_174.andOp_174_in0
	// controller for andOp_174.andOp_174_in1
	// Insensitive connections
	always @(*) begin
		andOp_174_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_174_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_175.andOp_175_in0
	// controller for andOp_175.andOp_175_in1
	// Insensitive connections
	always @(*) begin
		andOp_175_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_175_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_176.andOp_176_in0
	// controller for andOp_176.andOp_176_in1
	// Insensitive connections
	always @(*) begin
		andOp_176_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_176_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_177.andOp_177_in0
	// controller for andOp_177.andOp_177_in1
	// Insensitive connections
	always @(*) begin
		andOp_177_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_177_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_179.andOp_179_in0
	// controller for andOp_179.andOp_179_in1
	// Insensitive connections
	always @(*) begin
		andOp_179_in0 = valid ? notOp_178_out : notOp_178_out;
		andOp_179_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_181.andOp_181_in0
	// controller for andOp_181.andOp_181_in1
	// Insensitive connections
	always @(*) begin
		andOp_181_in0 = valid ? notOp_180_out : notOp_180_out;
		andOp_181_in1 = valid ? andOp_179_out : andOp_179_out;
	end
	// controller for andOp_183.andOp_183_in0
	// controller for andOp_183.andOp_183_in1
	// Insensitive connections
	always @(*) begin
		andOp_183_in0 = valid ? notOp_182_out : notOp_182_out;
		andOp_183_in1 = valid ? andOp_181_out : andOp_181_out;
	end
	// controller for andOp_185.andOp_185_in0
	// controller for andOp_185.andOp_185_in1
	// Insensitive connections
	always @(*) begin
		andOp_185_in0 = valid ? notOp_184_out : notOp_184_out;
		andOp_185_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_187.andOp_187_in0
	// controller for andOp_187.andOp_187_in1
	// Insensitive connections
	always @(*) begin
		andOp_187_in0 = valid ? notOp_186_out : notOp_186_out;
		andOp_187_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_189.andOp_189_in0
	// controller for andOp_189.andOp_189_in1
	// Insensitive connections
	always @(*) begin
		andOp_189_in0 = valid ? notOp_188_out : notOp_188_out;
		andOp_189_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_191.andOp_191_in0
	// controller for andOp_191.andOp_191_in1
	// Insensitive connections
	always @(*) begin
		andOp_191_in0 = valid ? notOp_190_out : notOp_190_out;
		andOp_191_in1 = valid ? andOp_189_out : andOp_189_out;
	end
	// controller for andOp_193.andOp_193_in0
	// controller for andOp_193.andOp_193_in1
	// Insensitive connections
	always @(*) begin
		andOp_193_in0 = valid ? notOp_192_out : notOp_192_out;
		andOp_193_in1 = valid ? andOp_191_out : andOp_191_out;
	end
	// controller for andOp_194.andOp_194_in0
	// controller for andOp_194.andOp_194_in1
	// Insensitive connections
	always @(*) begin
		andOp_194_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_194_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_195.andOp_195_in0
	// controller for andOp_195.andOp_195_in1
	// Insensitive connections
	always @(*) begin
		andOp_195_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_195_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_196.andOp_196_in0
	// controller for andOp_196.andOp_196_in1
	// Insensitive connections
	always @(*) begin
		andOp_196_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_196_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_197.andOp_197_in0
	// controller for andOp_197.andOp_197_in1
	// Insensitive connections
	always @(*) begin
		andOp_197_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_197_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_199.andOp_199_in0
	// controller for andOp_199.andOp_199_in1
	// Insensitive connections
	always @(*) begin
		andOp_199_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_199_in1 = valid ? notOp_198_out : notOp_198_out;
	end
	// controller for andOp_200.andOp_200_in0
	// controller for andOp_200.andOp_200_in1
	// Insensitive connections
	always @(*) begin
		andOp_200_in0 = valid ? 1'd0 : 1'd0;
		andOp_200_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_202.andOp_202_in0
	// controller for andOp_202.andOp_202_in1
	// Insensitive connections
	always @(*) begin
		andOp_202_in0 = valid ? andOp_199_out : andOp_199_out;
		andOp_202_in1 = valid ? eq_201_out : eq_201_out;
	end
	// controller for andOp_204.andOp_204_in0
	// controller for andOp_204.andOp_204_in1
	// Insensitive connections
	always @(*) begin
		andOp_204_in0 = valid ? andOp_199_out : andOp_199_out;
		andOp_204_in1 = valid ? notOp_203_out : notOp_203_out;
	end
	// controller for andOp_206.andOp_206_in0
	// controller for andOp_206.andOp_206_in1
	// Insensitive connections
	always @(*) begin
		andOp_206_in0 = valid ? andOp_204_out : andOp_204_out;
		andOp_206_in1 = valid ? eq_205_out : eq_205_out;
	end
	// controller for andOp_208.andOp_208_in0
	// controller for andOp_208.andOp_208_in1
	// Insensitive connections
	always @(*) begin
		andOp_208_in0 = valid ? andOp_204_out : andOp_204_out;
		andOp_208_in1 = valid ? eq_207_out : eq_207_out;
	end
	// controller for andOp_210.andOp_210_in0
	// controller for andOp_210.andOp_210_in1
	// Insensitive connections
	always @(*) begin
		andOp_210_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_210_in1 = valid ? notOp_209_out : notOp_209_out;
	end
	// controller for andOp_211.andOp_211_in0
	// controller for andOp_211.andOp_211_in1
	// Insensitive connections
	always @(*) begin
		andOp_211_in0 = valid ? 1'd0 : 1'd0;
		andOp_211_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_213.andOp_213_in0
	// controller for andOp_213.andOp_213_in1
	// Insensitive connections
	always @(*) begin
		andOp_213_in0 = valid ? andOp_210_out : andOp_210_out;
		andOp_213_in1 = valid ? eq_212_out : eq_212_out;
	end
	// controller for andOp_215.andOp_215_in0
	// controller for andOp_215.andOp_215_in1
	// Insensitive connections
	always @(*) begin
		andOp_215_in0 = valid ? andOp_210_out : andOp_210_out;
		andOp_215_in1 = valid ? notOp_214_out : notOp_214_out;
	end
	// controller for andOp_217.andOp_217_in0
	// controller for andOp_217.andOp_217_in1
	// Insensitive connections
	always @(*) begin
		andOp_217_in0 = valid ? andOp_215_out : andOp_215_out;
		andOp_217_in1 = valid ? eq_216_out : eq_216_out;
	end
	// controller for andOp_219.andOp_219_in0
	// controller for andOp_219.andOp_219_in1
	// Insensitive connections
	always @(*) begin
		andOp_219_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_219_in1 = valid ? notOp_218_out : notOp_218_out;
	end
	// controller for andOp_220.andOp_220_in0
	// controller for andOp_220.andOp_220_in1
	// Insensitive connections
	always @(*) begin
		andOp_220_in0 = valid ? 1'd0 : 1'd0;
		andOp_220_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_222.andOp_222_in0
	// controller for andOp_222.andOp_222_in1
	// Insensitive connections
	always @(*) begin
		andOp_222_in0 = valid ? andOp_219_out : andOp_219_out;
		andOp_222_in1 = valid ? eq_221_out : eq_221_out;
	end
	// controller for andOp_224.andOp_224_in0
	// controller for andOp_224.andOp_224_in1
	// Insensitive connections
	always @(*) begin
		andOp_224_in0 = valid ? andOp_219_out : andOp_219_out;
		andOp_224_in1 = valid ? notOp_223_out : notOp_223_out;
	end
	// controller for andOp_226.andOp_226_in0
	// controller for andOp_226.andOp_226_in1
	// Insensitive connections
	always @(*) begin
		andOp_226_in0 = valid ? andOp_224_out : andOp_224_out;
		andOp_226_in1 = valid ? eq_225_out : eq_225_out;
	end
	// controller for andOp_228.andOp_228_in0
	// controller for andOp_228.andOp_228_in1
	// Insensitive connections
	always @(*) begin
		andOp_228_in0 = valid ? andOp_224_out : andOp_224_out;
		andOp_228_in1 = valid ? eq_227_out : eq_227_out;
	end
	// controller for andOp_230.andOp_230_in0
	// controller for andOp_230.andOp_230_in1
	// Insensitive connections
	always @(*) begin
		andOp_230_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_230_in1 = valid ? notOp_229_out : notOp_229_out;
	end
	// controller for andOp_231.andOp_231_in0
	// controller for andOp_231.andOp_231_in1
	// Insensitive connections
	always @(*) begin
		andOp_231_in0 = valid ? 1'd0 : 1'd0;
		andOp_231_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_233.andOp_233_in0
	// controller for andOp_233.andOp_233_in1
	// Insensitive connections
	always @(*) begin
		andOp_233_in0 = valid ? andOp_230_out : andOp_230_out;
		andOp_233_in1 = valid ? eq_232_out : eq_232_out;
	end
	// controller for andOp_235.andOp_235_in0
	// controller for andOp_235.andOp_235_in1
	// Insensitive connections
	always @(*) begin
		andOp_235_in0 = valid ? andOp_230_out : andOp_230_out;
		andOp_235_in1 = valid ? notOp_234_out : notOp_234_out;
	end
	// controller for andOp_237.andOp_237_in0
	// controller for andOp_237.andOp_237_in1
	// Insensitive connections
	always @(*) begin
		andOp_237_in0 = valid ? andOp_235_out : andOp_235_out;
		andOp_237_in1 = valid ? eq_236_out : eq_236_out;
	end
	// controller for andOp_239.andOp_239_in0
	// controller for andOp_239.andOp_239_in1
	// Insensitive connections
	always @(*) begin
		andOp_239_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_239_in1 = valid ? notOp_238_out : notOp_238_out;
	end
	// controller for andOp_240.andOp_240_in0
	// controller for andOp_240.andOp_240_in1
	// Insensitive connections
	always @(*) begin
		andOp_240_in0 = valid ? 1'd0 : 1'd0;
		andOp_240_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_242.andOp_242_in0
	// controller for andOp_242.andOp_242_in1
	// Insensitive connections
	always @(*) begin
		andOp_242_in0 = valid ? andOp_239_out : andOp_239_out;
		andOp_242_in1 = valid ? eq_241_out : eq_241_out;
	end
	// controller for andOp_244.andOp_244_in0
	// controller for andOp_244.andOp_244_in1
	// Insensitive connections
	always @(*) begin
		andOp_244_in0 = valid ? andOp_239_out : andOp_239_out;
		andOp_244_in1 = valid ? notOp_243_out : notOp_243_out;
	end
	// controller for andOp_246.andOp_246_in0
	// controller for andOp_246.andOp_246_in1
	// Insensitive connections
	always @(*) begin
		andOp_246_in0 = valid ? andOp_244_out : andOp_244_out;
		andOp_246_in1 = valid ? eq_245_out : eq_245_out;
	end
	// controller for andOp_248.andOp_248_in0
	// controller for andOp_248.andOp_248_in1
	// Insensitive connections
	always @(*) begin
		andOp_248_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_248_in1 = valid ? notOp_247_out : notOp_247_out;
	end
	// controller for andOp_249.andOp_249_in0
	// controller for andOp_249.andOp_249_in1
	// Insensitive connections
	always @(*) begin
		andOp_249_in0 = valid ? 1'd0 : 1'd0;
		andOp_249_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_251.andOp_251_in0
	// controller for andOp_251.andOp_251_in1
	// Insensitive connections
	always @(*) begin
		andOp_251_in0 = valid ? andOp_248_out : andOp_248_out;
		andOp_251_in1 = valid ? eq_250_out : eq_250_out;
	end
	// controller for andOp_253.andOp_253_in0
	// controller for andOp_253.andOp_253_in1
	// Insensitive connections
	always @(*) begin
		andOp_253_in0 = valid ? andOp_248_out : andOp_248_out;
		andOp_253_in1 = valid ? notOp_252_out : notOp_252_out;
	end
	// controller for andOp_255.andOp_255_in0
	// controller for andOp_255.andOp_255_in1
	// Insensitive connections
	always @(*) begin
		andOp_255_in0 = valid ? andOp_253_out : andOp_253_out;
		andOp_255_in1 = valid ? eq_254_out : eq_254_out;
	end
	// controller for andOp_257.andOp_257_in0
	// controller for andOp_257.andOp_257_in1
	// Insensitive connections
	always @(*) begin
		andOp_257_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_257_in1 = valid ? notOp_256_out : notOp_256_out;
	end
	// controller for andOp_258.andOp_258_in0
	// controller for andOp_258.andOp_258_in1
	// Insensitive connections
	always @(*) begin
		andOp_258_in0 = valid ? 1'd0 : 1'd0;
		andOp_258_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_260.andOp_260_in0
	// controller for andOp_260.andOp_260_in1
	// Insensitive connections
	always @(*) begin
		andOp_260_in0 = valid ? andOp_257_out : andOp_257_out;
		andOp_260_in1 = valid ? eq_259_out : eq_259_out;
	end
	// controller for andOp_262.andOp_262_in0
	// controller for andOp_262.andOp_262_in1
	// Insensitive connections
	always @(*) begin
		andOp_262_in0 = valid ? andOp_257_out : andOp_257_out;
		andOp_262_in1 = valid ? notOp_261_out : notOp_261_out;
	end
	// controller for andOp_264.andOp_264_in0
	// controller for andOp_264.andOp_264_in1
	// Insensitive connections
	always @(*) begin
		andOp_264_in0 = valid ? andOp_262_out : andOp_262_out;
		andOp_264_in1 = valid ? eq_263_out : eq_263_out;
	end
	// controller for andOp_266.andOp_266_in0
	// controller for andOp_266.andOp_266_in1
	// Insensitive connections
	always @(*) begin
		andOp_266_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_266_in1 = valid ? notOp_265_out : notOp_265_out;
	end
	// controller for andOp_267.andOp_267_in0
	// controller for andOp_267.andOp_267_in1
	// Insensitive connections
	always @(*) begin
		andOp_267_in0 = valid ? 1'd0 : 1'd0;
		andOp_267_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_269.andOp_269_in0
	// controller for andOp_269.andOp_269_in1
	// Insensitive connections
	always @(*) begin
		andOp_269_in0 = valid ? andOp_266_out : andOp_266_out;
		andOp_269_in1 = valid ? eq_268_out : eq_268_out;
	end
	// controller for andOp_271.andOp_271_in0
	// controller for andOp_271.andOp_271_in1
	// Insensitive connections
	always @(*) begin
		andOp_271_in0 = valid ? andOp_266_out : andOp_266_out;
		andOp_271_in1 = valid ? notOp_270_out : notOp_270_out;
	end
	// controller for andOp_273.andOp_273_in0
	// controller for andOp_273.andOp_273_in1
	// Insensitive connections
	always @(*) begin
		andOp_273_in0 = valid ? andOp_271_out : andOp_271_out;
		andOp_273_in1 = valid ? eq_272_out : eq_272_out;
	end
	// controller for andOp_275.andOp_275_in0
	// controller for andOp_275.andOp_275_in1
	// Insensitive connections
	always @(*) begin
		andOp_275_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_275_in1 = valid ? notOp_274_out : notOp_274_out;
	end
	// controller for andOp_276.andOp_276_in0
	// controller for andOp_276.andOp_276_in1
	// Insensitive connections
	always @(*) begin
		andOp_276_in0 = valid ? 1'd0 : 1'd0;
		andOp_276_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_278.andOp_278_in0
	// controller for andOp_278.andOp_278_in1
	// Insensitive connections
	always @(*) begin
		andOp_278_in0 = valid ? andOp_275_out : andOp_275_out;
		andOp_278_in1 = valid ? eq_277_out : eq_277_out;
	end
	// controller for andOp_280.andOp_280_in0
	// controller for andOp_280.andOp_280_in1
	// Insensitive connections
	always @(*) begin
		andOp_280_in0 = valid ? andOp_275_out : andOp_275_out;
		andOp_280_in1 = valid ? notOp_279_out : notOp_279_out;
	end
	// controller for andOp_282.andOp_282_in0
	// controller for andOp_282.andOp_282_in1
	// Insensitive connections
	always @(*) begin
		andOp_282_in0 = valid ? andOp_280_out : andOp_280_out;
		andOp_282_in1 = valid ? eq_281_out : eq_281_out;
	end
	// controller for andOp_284.andOp_284_in0
	// controller for andOp_284.andOp_284_in1
	// Insensitive connections
	always @(*) begin
		andOp_284_in0 = valid ? andOp_280_out : andOp_280_out;
		andOp_284_in1 = valid ? eq_283_out : eq_283_out;
	end
	// controller for andOp_286.andOp_286_in0
	// controller for andOp_286.andOp_286_in1
	// Insensitive connections
	always @(*) begin
		andOp_286_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_286_in1 = valid ? notOp_285_out : notOp_285_out;
	end
	// controller for andOp_287.andOp_287_in0
	// controller for andOp_287.andOp_287_in1
	// Insensitive connections
	always @(*) begin
		andOp_287_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
		andOp_287_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_289.andOp_289_in0
	// controller for andOp_289.andOp_289_in1
	// Insensitive connections
	always @(*) begin
		andOp_289_in0 = valid ? andOp_286_out : andOp_286_out;
		andOp_289_in1 = valid ? eq_288_out : eq_288_out;
	end
	// controller for andOp_291.andOp_291_in0
	// controller for andOp_291.andOp_291_in1
	// Insensitive connections
	always @(*) begin
		andOp_291_in0 = valid ? andOp_286_out : andOp_286_out;
		andOp_291_in1 = valid ? notOp_290_out : notOp_290_out;
	end
	// controller for andOp_293.andOp_293_in0
	// controller for andOp_293.andOp_293_in1
	// Insensitive connections
	always @(*) begin
		andOp_293_in0 = valid ? andOp_291_out : andOp_291_out;
		andOp_293_in1 = valid ? eq_292_out : eq_292_out;
	end
	// controller for andOp_295.andOp_295_in0
	// controller for andOp_295.andOp_295_in1
	// Insensitive connections
	always @(*) begin
		andOp_295_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_295_in1 = valid ? notOp_294_out : notOp_294_out;
	end
	// controller for andOp_296.andOp_296_in0
	// controller for andOp_296.andOp_296_in1
	// Insensitive connections
	always @(*) begin
		andOp_296_in0 = valid ? 1'd0 : 1'd0;
		andOp_296_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_298.andOp_298_in0
	// controller for andOp_298.andOp_298_in1
	// Insensitive connections
	always @(*) begin
		andOp_298_in0 = valid ? andOp_295_out : andOp_295_out;
		andOp_298_in1 = valid ? eq_297_out : eq_297_out;
	end
	// controller for andOp_300.andOp_300_in0
	// controller for andOp_300.andOp_300_in1
	// Insensitive connections
	always @(*) begin
		andOp_300_in0 = valid ? andOp_295_out : andOp_295_out;
		andOp_300_in1 = valid ? notOp_299_out : notOp_299_out;
	end
	// controller for andOp_302.andOp_302_in0
	// controller for andOp_302.andOp_302_in1
	// Insensitive connections
	always @(*) begin
		andOp_302_in0 = valid ? andOp_300_out : andOp_300_out;
		andOp_302_in1 = valid ? eq_301_out : eq_301_out;
	end
	// controller for andOp_304.andOp_304_in0
	// controller for andOp_304.andOp_304_in1
	// Insensitive connections
	always @(*) begin
		andOp_304_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_304_in1 = valid ? notOp_303_out : notOp_303_out;
	end
	// controller for andOp_305.andOp_305_in0
	// controller for andOp_305.andOp_305_in1
	// Insensitive connections
	always @(*) begin
		andOp_305_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_305_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_307.andOp_307_in0
	// controller for andOp_307.andOp_307_in1
	// Insensitive connections
	always @(*) begin
		andOp_307_in0 = valid ? andOp_304_out : andOp_304_out;
		andOp_307_in1 = valid ? eq_306_out : eq_306_out;
	end
	// controller for andOp_309.andOp_309_in0
	// controller for andOp_309.andOp_309_in1
	// Insensitive connections
	always @(*) begin
		andOp_309_in0 = valid ? andOp_304_out : andOp_304_out;
		andOp_309_in1 = valid ? notOp_308_out : notOp_308_out;
	end
	// controller for andOp_311.andOp_311_in0
	// controller for andOp_311.andOp_311_in1
	// Insensitive connections
	always @(*) begin
		andOp_311_in0 = valid ? andOp_309_out : andOp_309_out;
		andOp_311_in1 = valid ? eq_310_out : eq_310_out;
	end
	// controller for andOp_313.andOp_313_in0
	// controller for andOp_313.andOp_313_in1
	// Insensitive connections
	always @(*) begin
		andOp_313_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_313_in1 = valid ? notOp_312_out : notOp_312_out;
	end
	// controller for andOp_314.andOp_314_in0
	// controller for andOp_314.andOp_314_in1
	// Insensitive connections
	always @(*) begin
		andOp_314_in0 = valid ? 1'd0 : 1'd0;
		andOp_314_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_316.andOp_316_in0
	// controller for andOp_316.andOp_316_in1
	// Insensitive connections
	always @(*) begin
		andOp_316_in0 = valid ? andOp_313_out : andOp_313_out;
		andOp_316_in1 = valid ? eq_315_out : eq_315_out;
	end
	// controller for andOp_318.andOp_318_in0
	// controller for andOp_318.andOp_318_in1
	// Insensitive connections
	always @(*) begin
		andOp_318_in0 = valid ? andOp_313_out : andOp_313_out;
		andOp_318_in1 = valid ? notOp_317_out : notOp_317_out;
	end
	// controller for andOp_320.andOp_320_in0
	// controller for andOp_320.andOp_320_in1
	// Insensitive connections
	always @(*) begin
		andOp_320_in0 = valid ? andOp_318_out : andOp_318_out;
		andOp_320_in1 = valid ? eq_319_out : eq_319_out;
	end
	// controller for andOp_322.andOp_322_in0
	// controller for andOp_322.andOp_322_in1
	// Insensitive connections
	always @(*) begin
		andOp_322_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_322_in1 = valid ? notOp_321_out : notOp_321_out;
	end
	// controller for andOp_323.andOp_323_in0
	// controller for andOp_323.andOp_323_in1
	// Insensitive connections
	always @(*) begin
		andOp_323_in0 = valid ? 1'd0 : 1'd0;
		andOp_323_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_325.andOp_325_in0
	// controller for andOp_325.andOp_325_in1
	// Insensitive connections
	always @(*) begin
		andOp_325_in0 = valid ? andOp_322_out : andOp_322_out;
		andOp_325_in1 = valid ? eq_324_out : eq_324_out;
	end
	// controller for andOp_327.andOp_327_in0
	// controller for andOp_327.andOp_327_in1
	// Insensitive connections
	always @(*) begin
		andOp_327_in0 = valid ? andOp_322_out : andOp_322_out;
		andOp_327_in1 = valid ? notOp_326_out : notOp_326_out;
	end
	// controller for andOp_329.andOp_329_in0
	// controller for andOp_329.andOp_329_in1
	// Insensitive connections
	always @(*) begin
		andOp_329_in0 = valid ? andOp_327_out : andOp_327_out;
		andOp_329_in1 = valid ? eq_328_out : eq_328_out;
	end
	// controller for andOp_331.andOp_331_in0
	// controller for andOp_331.andOp_331_in1
	// Insensitive connections
	always @(*) begin
		andOp_331_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_331_in1 = valid ? notOp_330_out : notOp_330_out;
	end
	// controller for andOp_332.andOp_332_in0
	// controller for andOp_332.andOp_332_in1
	// Insensitive connections
	always @(*) begin
		andOp_332_in0 = valid ? 1'd0 : 1'd0;
		andOp_332_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_334.andOp_334_in0
	// controller for andOp_334.andOp_334_in1
	// Insensitive connections
	always @(*) begin
		andOp_334_in0 = valid ? andOp_331_out : andOp_331_out;
		andOp_334_in1 = valid ? eq_333_out : eq_333_out;
	end
	// controller for andOp_336.andOp_336_in0
	// controller for andOp_336.andOp_336_in1
	// Insensitive connections
	always @(*) begin
		andOp_336_in0 = valid ? andOp_331_out : andOp_331_out;
		andOp_336_in1 = valid ? notOp_335_out : notOp_335_out;
	end
	// controller for andOp_338.andOp_338_in0
	// controller for andOp_338.andOp_338_in1
	// Insensitive connections
	always @(*) begin
		andOp_338_in0 = valid ? andOp_336_out : andOp_336_out;
		andOp_338_in1 = valid ? eq_337_out : eq_337_out;
	end
	// controller for andOp_340.andOp_340_in0
	// controller for andOp_340.andOp_340_in1
	// Insensitive connections
	always @(*) begin
		andOp_340_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_340_in1 = valid ? notOp_339_out : notOp_339_out;
	end
	// controller for andOp_341.andOp_341_in0
	// controller for andOp_341.andOp_341_in1
	// Insensitive connections
	always @(*) begin
		andOp_341_in0 = valid ? 1'd0 : 1'd0;
		andOp_341_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_343.andOp_343_in0
	// controller for andOp_343.andOp_343_in1
	// Insensitive connections
	always @(*) begin
		andOp_343_in0 = valid ? andOp_340_out : andOp_340_out;
		andOp_343_in1 = valid ? eq_342_out : eq_342_out;
	end
	// controller for andOp_345.andOp_345_in0
	// controller for andOp_345.andOp_345_in1
	// Insensitive connections
	always @(*) begin
		andOp_345_in0 = valid ? andOp_340_out : andOp_340_out;
		andOp_345_in1 = valid ? notOp_344_out : notOp_344_out;
	end
	// controller for andOp_347.andOp_347_in0
	// controller for andOp_347.andOp_347_in1
	// Insensitive connections
	always @(*) begin
		andOp_347_in0 = valid ? andOp_345_out : andOp_345_out;
		andOp_347_in1 = valid ? eq_346_out : eq_346_out;
	end
	// controller for andOp_349.andOp_349_in0
	// controller for andOp_349.andOp_349_in1
	// Insensitive connections
	always @(*) begin
		andOp_349_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_349_in1 = valid ? notOp_348_out : notOp_348_out;
	end
	// controller for andOp_350.andOp_350_in0
	// controller for andOp_350.andOp_350_in1
	// Insensitive connections
	always @(*) begin
		andOp_350_in0 = valid ? 1'd0 : 1'd0;
		andOp_350_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_352.andOp_352_in0
	// controller for andOp_352.andOp_352_in1
	// Insensitive connections
	always @(*) begin
		andOp_352_in0 = valid ? andOp_349_out : andOp_349_out;
		andOp_352_in1 = valid ? eq_351_out : eq_351_out;
	end
	// controller for andOp_354.andOp_354_in0
	// controller for andOp_354.andOp_354_in1
	// Insensitive connections
	always @(*) begin
		andOp_354_in0 = valid ? andOp_349_out : andOp_349_out;
		andOp_354_in1 = valid ? notOp_353_out : notOp_353_out;
	end
	// controller for andOp_356.andOp_356_in0
	// controller for andOp_356.andOp_356_in1
	// Insensitive connections
	always @(*) begin
		andOp_356_in0 = valid ? andOp_354_out : andOp_354_out;
		andOp_356_in1 = valid ? eq_355_out : eq_355_out;
	end
	// controller for andOp_358.andOp_358_in0
	// controller for andOp_358.andOp_358_in1
	// Insensitive connections
	always @(*) begin
		andOp_358_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_358_in1 = valid ? notOp_357_out : notOp_357_out;
	end
	// controller for andOp_359.andOp_359_in0
	// controller for andOp_359.andOp_359_in1
	// Insensitive connections
	always @(*) begin
		andOp_359_in0 = valid ? 1'd0 : 1'd0;
		andOp_359_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_361.andOp_361_in0
	// controller for andOp_361.andOp_361_in1
	// Insensitive connections
	always @(*) begin
		andOp_361_in0 = valid ? andOp_358_out : andOp_358_out;
		andOp_361_in1 = valid ? eq_360_out : eq_360_out;
	end
	// controller for andOp_363.andOp_363_in0
	// controller for andOp_363.andOp_363_in1
	// Insensitive connections
	always @(*) begin
		andOp_363_in0 = valid ? andOp_358_out : andOp_358_out;
		andOp_363_in1 = valid ? notOp_362_out : notOp_362_out;
	end
	// controller for andOp_365.andOp_365_in0
	// controller for andOp_365.andOp_365_in1
	// Insensitive connections
	always @(*) begin
		andOp_365_in0 = valid ? andOp_363_out : andOp_363_out;
		andOp_365_in1 = valid ? eq_364_out : eq_364_out;
	end
	// controller for andOp_367.andOp_367_in0
	// controller for andOp_367.andOp_367_in1
	// Insensitive connections
	always @(*) begin
		andOp_367_in0 = valid ? andOp_363_out : andOp_363_out;
		andOp_367_in1 = valid ? eq_366_out : eq_366_out;
	end
	// controller for andOp_369.andOp_369_in0
	// controller for andOp_369.andOp_369_in1
	// Insensitive connections
	always @(*) begin
		andOp_369_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_369_in1 = valid ? notOp_368_out : notOp_368_out;
	end
	// controller for andOp_370.andOp_370_in0
	// controller for andOp_370.andOp_370_in1
	// Insensitive connections
	always @(*) begin
		andOp_370_in0 = valid ? 1'd0 : 1'd0;
		andOp_370_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_372.andOp_372_in0
	// controller for andOp_372.andOp_372_in1
	// Insensitive connections
	always @(*) begin
		andOp_372_in0 = valid ? andOp_369_out : andOp_369_out;
		andOp_372_in1 = valid ? eq_371_out : eq_371_out;
	end
	// controller for andOp_374.andOp_374_in0
	// controller for andOp_374.andOp_374_in1
	// Insensitive connections
	always @(*) begin
		andOp_374_in0 = valid ? andOp_369_out : andOp_369_out;
		andOp_374_in1 = valid ? notOp_373_out : notOp_373_out;
	end
	// controller for andOp_376.andOp_376_in0
	// controller for andOp_376.andOp_376_in1
	// Insensitive connections
	always @(*) begin
		andOp_376_in0 = valid ? andOp_374_out : andOp_374_out;
		andOp_376_in1 = valid ? eq_375_out : eq_375_out;
	end
	// controller for andOp_378.andOp_378_in0
	// controller for andOp_378.andOp_378_in1
	// Insensitive connections
	always @(*) begin
		andOp_378_in0 = valid ? andOp_374_out : andOp_374_out;
		andOp_378_in1 = valid ? eq_377_out : eq_377_out;
	end
	// controller for andOp_380.andOp_380_in0
	// controller for andOp_380.andOp_380_in1
	// Insensitive connections
	always @(*) begin
		andOp_380_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_380_in1 = valid ? notOp_379_out : notOp_379_out;
	end
	// controller for andOp_381.andOp_381_in0
	// controller for andOp_381.andOp_381_in1
	// Insensitive connections
	always @(*) begin
		andOp_381_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_381_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_383.andOp_383_in0
	// controller for andOp_383.andOp_383_in1
	// Insensitive connections
	always @(*) begin
		andOp_383_in0 = valid ? andOp_380_out : andOp_380_out;
		andOp_383_in1 = valid ? eq_382_out : eq_382_out;
	end
	// controller for andOp_385.andOp_385_in0
	// controller for andOp_385.andOp_385_in1
	// Insensitive connections
	always @(*) begin
		andOp_385_in0 = valid ? andOp_380_out : andOp_380_out;
		andOp_385_in1 = valid ? notOp_384_out : notOp_384_out;
	end
	// controller for andOp_387.andOp_387_in0
	// controller for andOp_387.andOp_387_in1
	// Insensitive connections
	always @(*) begin
		andOp_387_in0 = valid ? andOp_385_out : andOp_385_out;
		andOp_387_in1 = valid ? eq_386_out : eq_386_out;
	end
	// controller for andOp_389.andOp_389_in0
	// controller for andOp_389.andOp_389_in1
	// Insensitive connections
	always @(*) begin
		andOp_389_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_389_in1 = valid ? notOp_388_out : notOp_388_out;
	end
	// controller for andOp_390.andOp_390_in0
	// controller for andOp_390.andOp_390_in1
	// Insensitive connections
	always @(*) begin
		andOp_390_in0 = valid ? 1'd0 : 1'd0;
		andOp_390_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_392.andOp_392_in0
	// controller for andOp_392.andOp_392_in1
	// Insensitive connections
	always @(*) begin
		andOp_392_in0 = valid ? andOp_389_out : andOp_389_out;
		andOp_392_in1 = valid ? eq_391_out : eq_391_out;
	end
	// controller for andOp_394.andOp_394_in0
	// controller for andOp_394.andOp_394_in1
	// Insensitive connections
	always @(*) begin
		andOp_394_in0 = valid ? andOp_389_out : andOp_389_out;
		andOp_394_in1 = valid ? notOp_393_out : notOp_393_out;
	end
	// controller for andOp_396.andOp_396_in0
	// controller for andOp_396.andOp_396_in1
	// Insensitive connections
	always @(*) begin
		andOp_396_in0 = valid ? andOp_394_out : andOp_394_out;
		andOp_396_in1 = valid ? eq_395_out : eq_395_out;
	end
	// controller for andOp_398.andOp_398_in0
	// controller for andOp_398.andOp_398_in1
	// Insensitive connections
	always @(*) begin
		andOp_398_in0 = valid ? andOp_394_out : andOp_394_out;
		andOp_398_in1 = valid ? eq_397_out : eq_397_out;
	end
	// controller for andOp_400.andOp_400_in0
	// controller for andOp_400.andOp_400_in1
	// Insensitive connections
	always @(*) begin
		andOp_400_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_400_in1 = valid ? notOp_399_out : notOp_399_out;
	end
	// controller for andOp_401.andOp_401_in0
	// controller for andOp_401.andOp_401_in1
	// Insensitive connections
	always @(*) begin
		andOp_401_in0 = valid ? 1'd0 : 1'd0;
		andOp_401_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_403.andOp_403_in0
	// controller for andOp_403.andOp_403_in1
	// Insensitive connections
	always @(*) begin
		andOp_403_in0 = valid ? andOp_400_out : andOp_400_out;
		andOp_403_in1 = valid ? eq_402_out : eq_402_out;
	end
	// controller for andOp_405.andOp_405_in0
	// controller for andOp_405.andOp_405_in1
	// Insensitive connections
	always @(*) begin
		andOp_405_in0 = valid ? andOp_400_out : andOp_400_out;
		andOp_405_in1 = valid ? notOp_404_out : notOp_404_out;
	end
	// controller for andOp_407.andOp_407_in0
	// controller for andOp_407.andOp_407_in1
	// Insensitive connections
	always @(*) begin
		andOp_407_in0 = valid ? andOp_405_out : andOp_405_out;
		andOp_407_in1 = valid ? eq_406_out : eq_406_out;
	end
	// controller for andOp_409.andOp_409_in0
	// controller for andOp_409.andOp_409_in1
	// Insensitive connections
	always @(*) begin
		andOp_409_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_409_in1 = valid ? notOp_408_out : notOp_408_out;
	end
	// controller for andOp_410.andOp_410_in0
	// controller for andOp_410.andOp_410_in1
	// Insensitive connections
	always @(*) begin
		andOp_410_in0 = valid ? 1'd0 : 1'd0;
		andOp_410_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_412.andOp_412_in0
	// controller for andOp_412.andOp_412_in1
	// Insensitive connections
	always @(*) begin
		andOp_412_in0 = valid ? andOp_409_out : andOp_409_out;
		andOp_412_in1 = valid ? eq_411_out : eq_411_out;
	end
	// controller for andOp_414.andOp_414_in0
	// controller for andOp_414.andOp_414_in1
	// Insensitive connections
	always @(*) begin
		andOp_414_in0 = valid ? andOp_409_out : andOp_409_out;
		andOp_414_in1 = valid ? notOp_413_out : notOp_413_out;
	end
	// controller for andOp_416.andOp_416_in0
	// controller for andOp_416.andOp_416_in1
	// Insensitive connections
	always @(*) begin
		andOp_416_in0 = valid ? andOp_414_out : andOp_414_out;
		andOp_416_in1 = valid ? eq_415_out : eq_415_out;
	end
	// controller for andOp_418.andOp_418_in0
	// controller for andOp_418.andOp_418_in1
	// Insensitive connections
	always @(*) begin
		andOp_418_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_418_in1 = valid ? notOp_417_out : notOp_417_out;
	end
	// controller for andOp_419.andOp_419_in0
	// controller for andOp_419.andOp_419_in1
	// Insensitive connections
	always @(*) begin
		andOp_419_in0 = valid ? 1'd0 : 1'd0;
		andOp_419_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_421.andOp_421_in0
	// controller for andOp_421.andOp_421_in1
	// Insensitive connections
	always @(*) begin
		andOp_421_in0 = valid ? andOp_418_out : andOp_418_out;
		andOp_421_in1 = valid ? eq_420_out : eq_420_out;
	end
	// controller for andOp_423.andOp_423_in0
	// controller for andOp_423.andOp_423_in1
	// Insensitive connections
	always @(*) begin
		andOp_423_in0 = valid ? andOp_418_out : andOp_418_out;
		andOp_423_in1 = valid ? notOp_422_out : notOp_422_out;
	end
	// controller for andOp_425.andOp_425_in0
	// controller for andOp_425.andOp_425_in1
	// Insensitive connections
	always @(*) begin
		andOp_425_in0 = valid ? andOp_423_out : andOp_423_out;
		andOp_425_in1 = valid ? eq_424_out : eq_424_out;
	end
	// controller for andOp_427.andOp_427_in0
	// controller for andOp_427.andOp_427_in1
	// Insensitive connections
	always @(*) begin
		andOp_427_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_427_in1 = valid ? notOp_426_out : notOp_426_out;
	end
	// controller for andOp_428.andOp_428_in0
	// controller for andOp_428.andOp_428_in1
	// Insensitive connections
	always @(*) begin
		andOp_428_in0 = valid ? 1'd0 : 1'd0;
		andOp_428_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_430.andOp_430_in0
	// controller for andOp_430.andOp_430_in1
	// Insensitive connections
	always @(*) begin
		andOp_430_in0 = valid ? andOp_427_out : andOp_427_out;
		andOp_430_in1 = valid ? eq_429_out : eq_429_out;
	end
	// controller for andOp_432.andOp_432_in0
	// controller for andOp_432.andOp_432_in1
	// Insensitive connections
	always @(*) begin
		andOp_432_in0 = valid ? andOp_427_out : andOp_427_out;
		andOp_432_in1 = valid ? notOp_431_out : notOp_431_out;
	end
	// controller for andOp_434.andOp_434_in0
	// controller for andOp_434.andOp_434_in1
	// Insensitive connections
	always @(*) begin
		andOp_434_in0 = valid ? andOp_432_out : andOp_432_out;
		andOp_434_in1 = valid ? eq_433_out : eq_433_out;
	end
	// controller for andOp_436.andOp_436_in0
	// controller for andOp_436.andOp_436_in1
	// Insensitive connections
	always @(*) begin
		andOp_436_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_436_in1 = valid ? notOp_435_out : notOp_435_out;
	end
	// controller for andOp_437.andOp_437_in0
	// controller for andOp_437.andOp_437_in1
	// Insensitive connections
	always @(*) begin
		andOp_437_in0 = valid ? 1'd0 : 1'd0;
		andOp_437_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_439.andOp_439_in0
	// controller for andOp_439.andOp_439_in1
	// Insensitive connections
	always @(*) begin
		andOp_439_in0 = valid ? andOp_436_out : andOp_436_out;
		andOp_439_in1 = valid ? eq_438_out : eq_438_out;
	end
	// controller for andOp_441.andOp_441_in0
	// controller for andOp_441.andOp_441_in1
	// Insensitive connections
	always @(*) begin
		andOp_441_in0 = valid ? andOp_436_out : andOp_436_out;
		andOp_441_in1 = valid ? notOp_440_out : notOp_440_out;
	end
	// controller for andOp_443.andOp_443_in0
	// controller for andOp_443.andOp_443_in1
	// Insensitive connections
	always @(*) begin
		andOp_443_in0 = valid ? andOp_441_out : andOp_441_out;
		andOp_443_in1 = valid ? eq_442_out : eq_442_out;
	end
	// controller for andOp_445.andOp_445_in0
	// controller for andOp_445.andOp_445_in1
	// Insensitive connections
	always @(*) begin
		andOp_445_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_445_in1 = valid ? notOp_444_out : notOp_444_out;
	end
	// controller for andOp_446.andOp_446_in0
	// controller for andOp_446.andOp_446_in1
	// Insensitive connections
	always @(*) begin
		andOp_446_in0 = valid ? 1'd0 : 1'd0;
		andOp_446_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_448.andOp_448_in0
	// controller for andOp_448.andOp_448_in1
	// Insensitive connections
	always @(*) begin
		andOp_448_in0 = valid ? andOp_445_out : andOp_445_out;
		andOp_448_in1 = valid ? eq_447_out : eq_447_out;
	end
	// controller for andOp_45.andOp_45_in0
	// controller for andOp_45.andOp_45_in1
	// Insensitive connections
	always @(*) begin
		andOp_45_in0 = valid ? bb_0_active_in_state_1_out_data : bb_0_active_in_state_1_out_data;
		andOp_45_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_450.andOp_450_in0
	// controller for andOp_450.andOp_450_in1
	// Insensitive connections
	always @(*) begin
		andOp_450_in0 = valid ? andOp_445_out : andOp_445_out;
		andOp_450_in1 = valid ? notOp_449_out : notOp_449_out;
	end
	// controller for andOp_452.andOp_452_in0
	// controller for andOp_452.andOp_452_in1
	// Insensitive connections
	always @(*) begin
		andOp_452_in0 = valid ? andOp_450_out : andOp_450_out;
		andOp_452_in1 = valid ? eq_451_out : eq_451_out;
	end
	// controller for andOp_454.andOp_454_in0
	// controller for andOp_454.andOp_454_in1
	// Insensitive connections
	always @(*) begin
		andOp_454_in0 = valid ? andOp_450_out : andOp_450_out;
		andOp_454_in1 = valid ? eq_453_out : eq_453_out;
	end
	// controller for andOp_456.andOp_456_in0
	// controller for andOp_456.andOp_456_in1
	// Insensitive connections
	always @(*) begin
		andOp_456_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_456_in1 = valid ? notOp_455_out : notOp_455_out;
	end
	// controller for andOp_457.andOp_457_in0
	// controller for andOp_457.andOp_457_in1
	// Insensitive connections
	always @(*) begin
		andOp_457_in0 = valid ? 1'd0 : 1'd0;
		andOp_457_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_459.andOp_459_in0
	// controller for andOp_459.andOp_459_in1
	// Insensitive connections
	always @(*) begin
		andOp_459_in0 = valid ? andOp_456_out : andOp_456_out;
		andOp_459_in1 = valid ? eq_458_out : eq_458_out;
	end
	// controller for andOp_46.andOp_46_in0
	// controller for andOp_46.andOp_46_in1
	// Insensitive connections
	always @(*) begin
		andOp_46_in0 = valid ? andOp_45_out : andOp_45_out;
		andOp_46_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_461.andOp_461_in0
	// controller for andOp_461.andOp_461_in1
	// Insensitive connections
	always @(*) begin
		andOp_461_in0 = valid ? andOp_456_out : andOp_456_out;
		andOp_461_in1 = valid ? notOp_460_out : notOp_460_out;
	end
	// controller for andOp_463.andOp_463_in0
	// controller for andOp_463.andOp_463_in1
	// Insensitive connections
	always @(*) begin
		andOp_463_in0 = valid ? andOp_461_out : andOp_461_out;
		andOp_463_in1 = valid ? eq_462_out : eq_462_out;
	end
	// controller for andOp_465.andOp_465_in0
	// controller for andOp_465.andOp_465_in1
	// Insensitive connections
	always @(*) begin
		andOp_465_in0 = valid ? andOp_461_out : andOp_461_out;
		andOp_465_in1 = valid ? eq_464_out : eq_464_out;
	end
	// controller for andOp_467.andOp_467_in0
	// controller for andOp_467.andOp_467_in1
	// Insensitive connections
	always @(*) begin
		andOp_467_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_467_in1 = valid ? notOp_466_out : notOp_466_out;
	end
	// controller for andOp_468.andOp_468_in0
	// controller for andOp_468.andOp_468_in1
	// Insensitive connections
	always @(*) begin
		andOp_468_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_468_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_470.andOp_470_in0
	// controller for andOp_470.andOp_470_in1
	// Insensitive connections
	always @(*) begin
		andOp_470_in0 = valid ? andOp_467_out : andOp_467_out;
		andOp_470_in1 = valid ? eq_469_out : eq_469_out;
	end
	// controller for andOp_472.andOp_472_in0
	// controller for andOp_472.andOp_472_in1
	// Insensitive connections
	always @(*) begin
		andOp_472_in0 = valid ? andOp_467_out : andOp_467_out;
		andOp_472_in1 = valid ? notOp_471_out : notOp_471_out;
	end
	// controller for andOp_474.andOp_474_in0
	// controller for andOp_474.andOp_474_in1
	// Insensitive connections
	always @(*) begin
		andOp_474_in0 = valid ? andOp_472_out : andOp_472_out;
		andOp_474_in1 = valid ? eq_473_out : eq_473_out;
	end
	// controller for andOp_476.andOp_476_in0
	// controller for andOp_476.andOp_476_in1
	// Insensitive connections
	always @(*) begin
		andOp_476_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_476_in1 = valid ? notOp_475_out : notOp_475_out;
	end
	// controller for andOp_477.andOp_477_in0
	// controller for andOp_477.andOp_477_in1
	// Insensitive connections
	always @(*) begin
		andOp_477_in0 = valid ? 1'd0 : 1'd0;
		andOp_477_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_479.andOp_479_in0
	// controller for andOp_479.andOp_479_in1
	// Insensitive connections
	always @(*) begin
		andOp_479_in0 = valid ? andOp_476_out : andOp_476_out;
		andOp_479_in1 = valid ? eq_478_out : eq_478_out;
	end
	// controller for andOp_48.andOp_48_in0
	// controller for andOp_48.andOp_48_in1
	// Insensitive connections
	always @(*) begin
		andOp_48_in0 = valid ? bb_8_active_in_state_1_out_data : bb_8_active_in_state_1_out_data;
		andOp_48_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_481.andOp_481_in0
	// controller for andOp_481.andOp_481_in1
	// Insensitive connections
	always @(*) begin
		andOp_481_in0 = valid ? andOp_476_out : andOp_476_out;
		andOp_481_in1 = valid ? notOp_480_out : notOp_480_out;
	end
	// controller for andOp_483.andOp_483_in0
	// controller for andOp_483.andOp_483_in1
	// Insensitive connections
	always @(*) begin
		andOp_483_in0 = valid ? andOp_481_out : andOp_481_out;
		andOp_483_in1 = valid ? eq_482_out : eq_482_out;
	end
	// controller for andOp_485.andOp_485_in0
	// controller for andOp_485.andOp_485_in1
	// Insensitive connections
	always @(*) begin
		andOp_485_in0 = valid ? andOp_481_out : andOp_481_out;
		andOp_485_in1 = valid ? eq_484_out : eq_484_out;
	end
	// controller for andOp_487.andOp_487_in0
	// controller for andOp_487.andOp_487_in1
	// Insensitive connections
	always @(*) begin
		andOp_487_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_487_in1 = valid ? notOp_486_out : notOp_486_out;
	end
	// controller for andOp_488.andOp_488_in0
	// controller for andOp_488.andOp_488_in1
	// Insensitive connections
	always @(*) begin
		andOp_488_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_488_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_49.andOp_49_in0
	// controller for andOp_49.andOp_49_in1
	// Insensitive connections
	always @(*) begin
		andOp_49_in0 = valid ? andOp_48_out : andOp_48_out;
		andOp_49_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_490.andOp_490_in0
	// controller for andOp_490.andOp_490_in1
	// Insensitive connections
	always @(*) begin
		andOp_490_in0 = valid ? andOp_487_out : andOp_487_out;
		andOp_490_in1 = valid ? eq_489_out : eq_489_out;
	end
	// controller for andOp_492.andOp_492_in0
	// controller for andOp_492.andOp_492_in1
	// Insensitive connections
	always @(*) begin
		andOp_492_in0 = valid ? andOp_487_out : andOp_487_out;
		andOp_492_in1 = valid ? notOp_491_out : notOp_491_out;
	end
	// controller for andOp_494.andOp_494_in0
	// controller for andOp_494.andOp_494_in1
	// Insensitive connections
	always @(*) begin
		andOp_494_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_494_in1 = valid ? notOp_493_out : notOp_493_out;
	end
	// controller for andOp_495.andOp_495_in0
	// controller for andOp_495.andOp_495_in1
	// Insensitive connections
	always @(*) begin
		andOp_495_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_495_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_497.andOp_497_in0
	// controller for andOp_497.andOp_497_in1
	// Insensitive connections
	always @(*) begin
		andOp_497_in0 = valid ? andOp_494_out : andOp_494_out;
		andOp_497_in1 = valid ? eq_496_out : eq_496_out;
	end
	// controller for andOp_499.andOp_499_in0
	// controller for andOp_499.andOp_499_in1
	// Insensitive connections
	always @(*) begin
		andOp_499_in0 = valid ? andOp_494_out : andOp_494_out;
		andOp_499_in1 = valid ? notOp_498_out : notOp_498_out;
	end
	// controller for andOp_501.andOp_501_in0
	// controller for andOp_501.andOp_501_in1
	// Insensitive connections
	always @(*) begin
		andOp_501_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_501_in1 = valid ? notOp_500_out : notOp_500_out;
	end
	// controller for andOp_502.andOp_502_in0
	// controller for andOp_502.andOp_502_in1
	// Insensitive connections
	always @(*) begin
		andOp_502_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_502_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_504.andOp_504_in0
	// controller for andOp_504.andOp_504_in1
	// Insensitive connections
	always @(*) begin
		andOp_504_in0 = valid ? andOp_501_out : andOp_501_out;
		andOp_504_in1 = valid ? eq_503_out : eq_503_out;
	end
	// controller for andOp_506.andOp_506_in0
	// controller for andOp_506.andOp_506_in1
	// Insensitive connections
	always @(*) begin
		andOp_506_in0 = valid ? andOp_501_out : andOp_501_out;
		andOp_506_in1 = valid ? notOp_505_out : notOp_505_out;
	end
	// controller for andOp_508.andOp_508_in0
	// controller for andOp_508.andOp_508_in1
	// Insensitive connections
	always @(*) begin
		andOp_508_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_508_in1 = valid ? notOp_507_out : notOp_507_out;
	end
	// controller for andOp_509.andOp_509_in0
	// controller for andOp_509.andOp_509_in1
	// Insensitive connections
	always @(*) begin
		andOp_509_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_509_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_51.andOp_51_in0
	// controller for andOp_51.andOp_51_in1
	// Insensitive connections
	always @(*) begin
		andOp_51_in0 = valid ? bb_0_active_in_state_1_out_data : bb_0_active_in_state_1_out_data;
		andOp_51_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_511.andOp_511_in0
	// controller for andOp_511.andOp_511_in1
	// Insensitive connections
	always @(*) begin
		andOp_511_in0 = valid ? andOp_508_out : andOp_508_out;
		andOp_511_in1 = valid ? eq_510_out : eq_510_out;
	end
	// controller for andOp_513.andOp_513_in0
	// controller for andOp_513.andOp_513_in1
	// Insensitive connections
	always @(*) begin
		andOp_513_in0 = valid ? andOp_508_out : andOp_508_out;
		andOp_513_in1 = valid ? notOp_512_out : notOp_512_out;
	end
	// controller for andOp_515.andOp_515_in0
	// controller for andOp_515.andOp_515_in1
	// Insensitive connections
	always @(*) begin
		andOp_515_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_515_in1 = valid ? notOp_514_out : notOp_514_out;
	end
	// controller for andOp_516.andOp_516_in0
	// controller for andOp_516.andOp_516_in1
	// Insensitive connections
	always @(*) begin
		andOp_516_in0 = valid ? 1'd0 : 1'd0;
		andOp_516_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_518.andOp_518_in0
	// controller for andOp_518.andOp_518_in1
	// Insensitive connections
	always @(*) begin
		andOp_518_in0 = valid ? andOp_515_out : andOp_515_out;
		andOp_518_in1 = valid ? eq_517_out : eq_517_out;
	end
	// controller for andOp_52.andOp_52_in0
	// controller for andOp_52.andOp_52_in1
	// Insensitive connections
	always @(*) begin
		andOp_52_in0 = valid ? andOp_51_out : andOp_51_out;
		andOp_52_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_520.andOp_520_in0
	// controller for andOp_520.andOp_520_in1
	// Insensitive connections
	always @(*) begin
		andOp_520_in0 = valid ? andOp_515_out : andOp_515_out;
		andOp_520_in1 = valid ? notOp_519_out : notOp_519_out;
	end
	// controller for andOp_522.andOp_522_in0
	// controller for andOp_522.andOp_522_in1
	// Insensitive connections
	always @(*) begin
		andOp_522_in0 = valid ? andOp_520_out : andOp_520_out;
		andOp_522_in1 = valid ? eq_521_out : eq_521_out;
	end
	// controller for andOp_524.andOp_524_in0
	// controller for andOp_524.andOp_524_in1
	// Insensitive connections
	always @(*) begin
		andOp_524_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_524_in1 = valid ? notOp_523_out : notOp_523_out;
	end
	// controller for andOp_525.andOp_525_in0
	// controller for andOp_525.andOp_525_in1
	// Insensitive connections
	always @(*) begin
		andOp_525_in0 = valid ? 1'd0 : 1'd0;
		andOp_525_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_527.andOp_527_in0
	// controller for andOp_527.andOp_527_in1
	// Insensitive connections
	always @(*) begin
		andOp_527_in0 = valid ? andOp_524_out : andOp_524_out;
		andOp_527_in1 = valid ? eq_526_out : eq_526_out;
	end
	// controller for andOp_529.andOp_529_in0
	// controller for andOp_529.andOp_529_in1
	// Insensitive connections
	always @(*) begin
		andOp_529_in0 = valid ? andOp_524_out : andOp_524_out;
		andOp_529_in1 = valid ? notOp_528_out : notOp_528_out;
	end
	// controller for andOp_531.andOp_531_in0
	// controller for andOp_531.andOp_531_in1
	// Insensitive connections
	always @(*) begin
		andOp_531_in0 = valid ? andOp_529_out : andOp_529_out;
		andOp_531_in1 = valid ? eq_530_out : eq_530_out;
	end
	// controller for andOp_533.andOp_533_in0
	// controller for andOp_533.andOp_533_in1
	// Insensitive connections
	always @(*) begin
		andOp_533_in0 = valid ? andOp_529_out : andOp_529_out;
		andOp_533_in1 = valid ? eq_532_out : eq_532_out;
	end
	// controller for andOp_535.andOp_535_in0
	// controller for andOp_535.andOp_535_in1
	// Insensitive connections
	always @(*) begin
		andOp_535_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_535_in1 = valid ? notOp_534_out : notOp_534_out;
	end
	// controller for andOp_536.andOp_536_in0
	// controller for andOp_536.andOp_536_in1
	// Insensitive connections
	always @(*) begin
		andOp_536_in0 = valid ? 1'd0 : 1'd0;
		andOp_536_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_538.andOp_538_in0
	// controller for andOp_538.andOp_538_in1
	// Insensitive connections
	always @(*) begin
		andOp_538_in0 = valid ? andOp_535_out : andOp_535_out;
		andOp_538_in1 = valid ? eq_537_out : eq_537_out;
	end
	// controller for andOp_54.andOp_54_in0
	// controller for andOp_54.andOp_54_in1
	// Insensitive connections
	always @(*) begin
		andOp_54_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_54_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_540.andOp_540_in0
	// controller for andOp_540.andOp_540_in1
	// Insensitive connections
	always @(*) begin
		andOp_540_in0 = valid ? andOp_535_out : andOp_535_out;
		andOp_540_in1 = valid ? notOp_539_out : notOp_539_out;
	end
	// controller for andOp_542.andOp_542_in0
	// controller for andOp_542.andOp_542_in1
	// Insensitive connections
	always @(*) begin
		andOp_542_in0 = valid ? andOp_540_out : andOp_540_out;
		andOp_542_in1 = valid ? eq_541_out : eq_541_out;
	end
	// controller for andOp_544.andOp_544_in0
	// controller for andOp_544.andOp_544_in1
	// Insensitive connections
	always @(*) begin
		andOp_544_in0 = valid ? andOp_540_out : andOp_540_out;
		andOp_544_in1 = valid ? eq_543_out : eq_543_out;
	end
	// controller for andOp_546.andOp_546_in0
	// controller for andOp_546.andOp_546_in1
	// Insensitive connections
	always @(*) begin
		andOp_546_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_546_in1 = valid ? notOp_545_out : notOp_545_out;
	end
	// controller for andOp_547.andOp_547_in0
	// controller for andOp_547.andOp_547_in1
	// Insensitive connections
	always @(*) begin
		andOp_547_in0 = valid ? 1'd0 : 1'd0;
		andOp_547_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_549.andOp_549_in0
	// controller for andOp_549.andOp_549_in1
	// Insensitive connections
	always @(*) begin
		andOp_549_in0 = valid ? andOp_546_out : andOp_546_out;
		andOp_549_in1 = valid ? eq_548_out : eq_548_out;
	end
	// controller for andOp_55.andOp_55_in0
	// controller for andOp_55.andOp_55_in1
	// Insensitive connections
	always @(*) begin
		andOp_55_in0 = valid ? andOp_54_out : andOp_54_out;
		andOp_55_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_551.andOp_551_in0
	// controller for andOp_551.andOp_551_in1
	// Insensitive connections
	always @(*) begin
		andOp_551_in0 = valid ? andOp_546_out : andOp_546_out;
		andOp_551_in1 = valid ? notOp_550_out : notOp_550_out;
	end
	// controller for andOp_553.andOp_553_in0
	// controller for andOp_553.andOp_553_in1
	// Insensitive connections
	always @(*) begin
		andOp_553_in0 = valid ? andOp_551_out : andOp_551_out;
		andOp_553_in1 = valid ? eq_552_out : eq_552_out;
	end
	// controller for andOp_555.andOp_555_in0
	// controller for andOp_555.andOp_555_in1
	// Insensitive connections
	always @(*) begin
		andOp_555_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_555_in1 = valid ? notOp_554_out : notOp_554_out;
	end
	// controller for andOp_556.andOp_556_in0
	// controller for andOp_556.andOp_556_in1
	// Insensitive connections
	always @(*) begin
		andOp_556_in0 = valid ? 1'd0 : 1'd0;
		andOp_556_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_558.andOp_558_in0
	// controller for andOp_558.andOp_558_in1
	// Insensitive connections
	always @(*) begin
		andOp_558_in0 = valid ? andOp_555_out : andOp_555_out;
		andOp_558_in1 = valid ? eq_557_out : eq_557_out;
	end
	// controller for andOp_560.andOp_560_in0
	// controller for andOp_560.andOp_560_in1
	// Insensitive connections
	always @(*) begin
		andOp_560_in0 = valid ? andOp_555_out : andOp_555_out;
		andOp_560_in1 = valid ? notOp_559_out : notOp_559_out;
	end
	// controller for andOp_562.andOp_562_in0
	// controller for andOp_562.andOp_562_in1
	// Insensitive connections
	always @(*) begin
		andOp_562_in0 = valid ? andOp_560_out : andOp_560_out;
		andOp_562_in1 = valid ? eq_561_out : eq_561_out;
	end
	// controller for andOp_564.andOp_564_in0
	// controller for andOp_564.andOp_564_in1
	// Insensitive connections
	always @(*) begin
		andOp_564_in0 = valid ? andOp_560_out : andOp_560_out;
		andOp_564_in1 = valid ? eq_563_out : eq_563_out;
	end
	// controller for andOp_566.andOp_566_in0
	// controller for andOp_566.andOp_566_in1
	// Insensitive connections
	always @(*) begin
		andOp_566_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_566_in1 = valid ? notOp_565_out : notOp_565_out;
	end
	// controller for andOp_567.andOp_567_in0
	// controller for andOp_567.andOp_567_in1
	// Insensitive connections
	always @(*) begin
		andOp_567_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_567_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_569.andOp_569_in0
	// controller for andOp_569.andOp_569_in1
	// Insensitive connections
	always @(*) begin
		andOp_569_in0 = valid ? andOp_566_out : andOp_566_out;
		andOp_569_in1 = valid ? eq_568_out : eq_568_out;
	end
	// controller for andOp_57.andOp_57_in0
	// controller for andOp_57.andOp_57_in1
	// Insensitive connections
	always @(*) begin
		andOp_57_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
		andOp_57_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_571.andOp_571_in0
	// controller for andOp_571.andOp_571_in1
	// Insensitive connections
	always @(*) begin
		andOp_571_in0 = valid ? andOp_566_out : andOp_566_out;
		andOp_571_in1 = valid ? notOp_570_out : notOp_570_out;
	end
	// controller for andOp_573.andOp_573_in0
	// controller for andOp_573.andOp_573_in1
	// Insensitive connections
	always @(*) begin
		andOp_573_in0 = valid ? andOp_571_out : andOp_571_out;
		andOp_573_in1 = valid ? eq_572_out : eq_572_out;
	end
	// controller for andOp_575.andOp_575_in0
	// controller for andOp_575.andOp_575_in1
	// Insensitive connections
	always @(*) begin
		andOp_575_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_575_in1 = valid ? notOp_574_out : notOp_574_out;
	end
	// controller for andOp_576.andOp_576_in0
	// controller for andOp_576.andOp_576_in1
	// Insensitive connections
	always @(*) begin
		andOp_576_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_576_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_578.andOp_578_in0
	// controller for andOp_578.andOp_578_in1
	// Insensitive connections
	always @(*) begin
		andOp_578_in0 = valid ? andOp_575_out : andOp_575_out;
		andOp_578_in1 = valid ? eq_577_out : eq_577_out;
	end
	// controller for andOp_58.andOp_58_in0
	// controller for andOp_58.andOp_58_in1
	// Insensitive connections
	always @(*) begin
		andOp_58_in0 = valid ? andOp_57_out : andOp_57_out;
		andOp_58_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_580.andOp_580_in0
	// controller for andOp_580.andOp_580_in1
	// Insensitive connections
	always @(*) begin
		andOp_580_in0 = valid ? andOp_575_out : andOp_575_out;
		andOp_580_in1 = valid ? notOp_579_out : notOp_579_out;
	end
	// controller for andOp_582.andOp_582_in0
	// controller for andOp_582.andOp_582_in1
	// Insensitive connections
	always @(*) begin
		andOp_582_in0 = valid ? andOp_580_out : andOp_580_out;
		andOp_582_in1 = valid ? eq_581_out : eq_581_out;
	end
	// controller for andOp_584.andOp_584_in0
	// controller for andOp_584.andOp_584_in1
	// Insensitive connections
	always @(*) begin
		andOp_584_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_584_in1 = valid ? notOp_583_out : notOp_583_out;
	end
	// controller for andOp_585.andOp_585_in0
	// controller for andOp_585.andOp_585_in1
	// Insensitive connections
	always @(*) begin
		andOp_585_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_585_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_587.andOp_587_in0
	// controller for andOp_587.andOp_587_in1
	// Insensitive connections
	always @(*) begin
		andOp_587_in0 = valid ? andOp_584_out : andOp_584_out;
		andOp_587_in1 = valid ? eq_586_out : eq_586_out;
	end
	// controller for andOp_589.andOp_589_in0
	// controller for andOp_589.andOp_589_in1
	// Insensitive connections
	always @(*) begin
		andOp_589_in0 = valid ? andOp_584_out : andOp_584_out;
		andOp_589_in1 = valid ? notOp_588_out : notOp_588_out;
	end
	// controller for andOp_591.andOp_591_in0
	// controller for andOp_591.andOp_591_in1
	// Insensitive connections
	always @(*) begin
		andOp_591_in0 = valid ? andOp_589_out : andOp_589_out;
		andOp_591_in1 = valid ? eq_590_out : eq_590_out;
	end
	// controller for andOp_593.andOp_593_in0
	// controller for andOp_593.andOp_593_in1
	// Insensitive connections
	always @(*) begin
		andOp_593_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_593_in1 = valid ? notOp_592_out : notOp_592_out;
	end
	// controller for andOp_594.andOp_594_in0
	// controller for andOp_594.andOp_594_in1
	// Insensitive connections
	always @(*) begin
		andOp_594_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_594_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_596.andOp_596_in0
	// controller for andOp_596.andOp_596_in1
	// Insensitive connections
	always @(*) begin
		andOp_596_in0 = valid ? andOp_593_out : andOp_593_out;
		andOp_596_in1 = valid ? eq_595_out : eq_595_out;
	end
	// controller for andOp_598.andOp_598_in0
	// controller for andOp_598.andOp_598_in1
	// Insensitive connections
	always @(*) begin
		andOp_598_in0 = valid ? andOp_593_out : andOp_593_out;
		andOp_598_in1 = valid ? notOp_597_out : notOp_597_out;
	end
	// controller for andOp_60.andOp_60_in0
	// controller for andOp_60.andOp_60_in1
	// Insensitive connections
	always @(*) begin
		andOp_60_in0 = valid ? andOp_58_out : andOp_58_out;
		andOp_60_in1 = valid ? in_read_ready : in_read_ready;
	end
	// controller for andOp_600.andOp_600_in0
	// controller for andOp_600.andOp_600_in1
	// Insensitive connections
	always @(*) begin
		andOp_600_in0 = valid ? andOp_598_out : andOp_598_out;
		andOp_600_in1 = valid ? eq_599_out : eq_599_out;
	end
	// controller for andOp_602.andOp_602_in0
	// controller for andOp_602.andOp_602_in1
	// Insensitive connections
	always @(*) begin
		andOp_602_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_602_in1 = valid ? notOp_601_out : notOp_601_out;
	end
	// controller for andOp_603.andOp_603_in0
	// controller for andOp_603.andOp_603_in1
	// Insensitive connections
	always @(*) begin
		andOp_603_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_603_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_605.andOp_605_in0
	// controller for andOp_605.andOp_605_in1
	// Insensitive connections
	always @(*) begin
		andOp_605_in0 = valid ? andOp_602_out : andOp_602_out;
		andOp_605_in1 = valid ? eq_604_out : eq_604_out;
	end
	// controller for andOp_607.andOp_607_in0
	// controller for andOp_607.andOp_607_in1
	// Insensitive connections
	always @(*) begin
		andOp_607_in0 = valid ? andOp_602_out : andOp_602_out;
		andOp_607_in1 = valid ? notOp_606_out : notOp_606_out;
	end
	// controller for andOp_609.andOp_609_in0
	// controller for andOp_609.andOp_609_in1
	// Insensitive connections
	always @(*) begin
		andOp_609_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_609_in1 = valid ? notOp_608_out : notOp_608_out;
	end
	// controller for andOp_610.andOp_610_in0
	// controller for andOp_610.andOp_610_in1
	// Insensitive connections
	always @(*) begin
		andOp_610_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
		andOp_610_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_612.andOp_612_in0
	// controller for andOp_612.andOp_612_in1
	// Insensitive connections
	always @(*) begin
		andOp_612_in0 = valid ? andOp_609_out : andOp_609_out;
		andOp_612_in1 = valid ? eq_611_out : eq_611_out;
	end
	// controller for andOp_614.andOp_614_in0
	// controller for andOp_614.andOp_614_in1
	// Insensitive connections
	always @(*) begin
		andOp_614_in0 = valid ? andOp_609_out : andOp_609_out;
		andOp_614_in1 = valid ? notOp_613_out : notOp_613_out;
	end
	// controller for andOp_616.andOp_616_in0
	// controller for andOp_616.andOp_616_in1
	// Insensitive connections
	always @(*) begin
		andOp_616_in0 = valid ? andOp_614_out : andOp_614_out;
		andOp_616_in1 = valid ? eq_615_out : eq_615_out;
	end
	// controller for andOp_62.andOp_62_in0
	// controller for andOp_62.andOp_62_in1
	// Insensitive connections
	always @(*) begin
		andOp_62_in0 = valid ? andOp_58_out : andOp_58_out;
		andOp_62_in1 = valid ? notOp_61_out : notOp_61_out;
	end
	// controller for andOp_63.andOp_63_in0
	// controller for andOp_63.andOp_63_in1
	// Insensitive connections
	always @(*) begin
		andOp_63_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_63_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_64.andOp_64_in0
	// controller for andOp_64.andOp_64_in1
	// Insensitive connections
	always @(*) begin
		andOp_64_in0 = valid ? andOp_63_out : andOp_63_out;
		andOp_64_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_66.andOp_66_in0
	// controller for andOp_66.andOp_66_in1
	// Insensitive connections
	always @(*) begin
		andOp_66_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_66_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_67.andOp_67_in0
	// controller for andOp_67.andOp_67_in1
	// Insensitive connections
	always @(*) begin
		andOp_67_in0 = valid ? andOp_66_out : andOp_66_out;
		andOp_67_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_69.andOp_69_in0
	// controller for andOp_69.andOp_69_in1
	// Insensitive connections
	always @(*) begin
		andOp_69_in0 = valid ? andOp_67_out : andOp_67_out;
		andOp_69_in1 = valid ? icmp_tmp_6 : icmp_tmp_6;
	end
	// controller for andOp_71.andOp_71_in0
	// controller for andOp_71.andOp_71_in1
	// Insensitive connections
	always @(*) begin
		andOp_71_in0 = valid ? andOp_67_out : andOp_67_out;
		andOp_71_in1 = valid ? notOp_70_out : notOp_70_out;
	end
	// controller for andOp_72.andOp_72_in0
	// controller for andOp_72.andOp_72_in1
	// Insensitive connections
	always @(*) begin
		andOp_72_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_72_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_73.andOp_73_in0
	// controller for andOp_73.andOp_73_in1
	// Insensitive connections
	always @(*) begin
		andOp_73_in0 = valid ? andOp_72_out : andOp_72_out;
		andOp_73_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_75.andOp_75_in0
	// controller for andOp_75.andOp_75_in1
	// Insensitive connections
	always @(*) begin
		andOp_75_in0 = valid ? bb_5_active_in_state_4_out_data : bb_5_active_in_state_4_out_data;
		andOp_75_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_76.andOp_76_in0
	// controller for andOp_76.andOp_76_in1
	// Insensitive connections
	always @(*) begin
		andOp_76_in0 = valid ? andOp_75_out : andOp_75_out;
		andOp_76_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_78.andOp_78_in0
	// controller for andOp_78.andOp_78_in1
	// Insensitive connections
	always @(*) begin
		andOp_78_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
		andOp_78_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_79.andOp_79_in0
	// controller for andOp_79.andOp_79_in1
	// Insensitive connections
	always @(*) begin
		andOp_79_in0 = valid ? andOp_78_out : andOp_78_out;
		andOp_79_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_81.andOp_81_in0
	// controller for andOp_81.andOp_81_in1
	// Insensitive connections
	always @(*) begin
		andOp_81_in0 = valid ? andOp_79_out : andOp_79_out;
		andOp_81_in1 = valid ? out_write_ready : out_write_ready;
	end
	// controller for andOp_83.andOp_83_in0
	// controller for andOp_83.andOp_83_in1
	// Insensitive connections
	always @(*) begin
		andOp_83_in0 = valid ? andOp_79_out : andOp_79_out;
		andOp_83_in1 = valid ? notOp_82_out : notOp_82_out;
	end
	// controller for andOp_84.andOp_84_in0
	// controller for andOp_84.andOp_84_in1
	// Insensitive connections
	always @(*) begin
		andOp_84_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_84_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_85.andOp_85_in0
	// controller for andOp_85.andOp_85_in1
	// Insensitive connections
	always @(*) begin
		andOp_85_in0 = valid ? andOp_84_out : andOp_84_out;
		andOp_85_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_87.andOp_87_in0
	// controller for andOp_87.andOp_87_in1
	// Insensitive connections
	always @(*) begin
		andOp_87_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_87_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_88.andOp_88_in0
	// controller for andOp_88.andOp_88_in1
	// Insensitive connections
	always @(*) begin
		andOp_88_in0 = valid ? andOp_87_out : andOp_87_out;
		andOp_88_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_90.andOp_90_in0
	// controller for andOp_90.andOp_90_in1
	// Insensitive connections
	always @(*) begin
		andOp_90_in0 = valid ? andOp_88_out : andOp_88_out;
		andOp_90_in1 = valid ? icmp_tmp_6 : icmp_tmp_6;
	end
	// controller for andOp_92.andOp_92_in0
	// controller for andOp_92.andOp_92_in1
	// Insensitive connections
	always @(*) begin
		andOp_92_in0 = valid ? andOp_88_out : andOp_88_out;
		andOp_92_in1 = valid ? notOp_91_out : notOp_91_out;
	end
	// controller for andOp_93.andOp_93_in0
	// controller for andOp_93.andOp_93_in1
	// Insensitive connections
	always @(*) begin
		andOp_93_in0 = valid ? bb_1_active_in_state_4_out_data : bb_1_active_in_state_4_out_data;
		andOp_93_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_94.andOp_94_in0
	// controller for andOp_94.andOp_94_in1
	// Insensitive connections
	always @(*) begin
		andOp_94_in0 = valid ? andOp_93_out : andOp_93_out;
		andOp_94_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_96_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_active_in_state_1.bb_0_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_1_in_data = eq_99_out;
		end else begin
			bb_0_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_119_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_1.bb_0_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_123_out) begin 
			bb_0_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_2.bb_10_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_2_in_data = eq_104_out;
		end else begin
			bb_10_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_3.bb_10_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_3_in_data = eq_107_out;
		end else begin
			bb_10_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_2.bb_10_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_130_out) begin 
			bb_10_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_3.bb_10_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_134_out) begin 
			bb_10_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_4.bb_1_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_4_in_data = orOp_118_out;
		end else begin
			bb_1_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_4.bb_1_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_150_out) begin 
			bb_1_predecessor_in_state_4_in_data = 32'd4;
		end else if (eq_148_out) begin 
			bb_1_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_4.bb_2_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_4_in_data = orOp_116_out;
		end else begin
			bb_2_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_4.bb_2_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_147_out) begin 
			bb_2_predecessor_in_state_4_in_data = 32'd7;
		end else if (eq_145_out) begin 
			bb_2_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_1.bb_3_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_1_in_data = orOp_101_out;
		end else begin
			bb_3_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_1.bb_3_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_126_out) begin 
			bb_3_predecessor_in_state_1_in_data = 32'd0;
		end else if (eq_124_out) begin 
			bb_3_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_3.bb_4_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_3_in_data = orOp_106_out;
		end else begin
			bb_4_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_4.bb_4_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_4_in_data = eq_114_out;
		end else begin
			bb_4_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_3.bb_4_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_133_out) begin 
			bb_4_predecessor_in_state_3_in_data = 32'd10;
		end else if (eq_131_out) begin 
			bb_4_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_4.bb_4_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_144_out) begin 
			bb_4_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_5_active_in_state_4.bb_5_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_5_active_in_state_4_in_data = orOp_109_out;
		end else begin
			bb_5_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_5_predecessor_in_state_4.bb_5_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_137_out) begin 
			bb_5_predecessor_in_state_4_in_data = 32'd1;
		end else if (eq_135_out) begin 
			bb_5_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_5_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_6_active_in_state_4.bb_6_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_6_active_in_state_4_in_data = orOp_111_out;
		end else begin
			bb_6_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_6_predecessor_in_state_4.bb_6_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_140_out) begin 
			bb_6_predecessor_in_state_4_in_data = 32'd5;
		end else if (eq_138_out) begin 
			bb_6_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_6_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_7_active_in_state_4.bb_7_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_7_active_in_state_4_in_data = orOp_113_out;
		end else begin
			bb_7_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_7_predecessor_in_state_4.bb_7_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_143_out) begin 
			bb_7_predecessor_in_state_4_in_data = 32'd6;
		end else if (eq_141_out) begin 
			bb_7_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_7_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_8_active_in_state_1.bb_8_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_state_1_in_data = orOp_98_out;
		end else begin
			bb_8_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_8_predecessor_in_state_1.bb_8_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_122_out) begin 
			bb_8_predecessor_in_state_1_in_data = 32'd3;
		end else if (eq_120_out) begin 
			bb_8_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_8_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_9_active_in_state_1.bb_9_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_9_active_in_state_1_in_data = orOp_103_out;
		end else begin
			bb_9_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_9_predecessor_in_state_1.bb_9_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_129_out) begin 
			bb_9_predecessor_in_state_1_in_data = 32'd8;
		end else if (eq_127_out) begin 
			bb_9_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_9_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_46_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_47_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_1.br_0_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_52_out) begin 
			br_0_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_53_out) begin 
			br_0_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_2.br_10_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_64_out) begin 
			br_10_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_65_out) begin 
			br_10_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_3.br_10_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_73_out) begin 
			br_10_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_74_out) begin 
			br_10_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_1_happened_in_state_4.br_1_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_94_out) begin 
			br_1_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_95_out) begin 
			br_1_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_1_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_1.br_3_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_55_out) begin 
			br_3_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_56_out) begin 
			br_3_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_3.br_4_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_67_out) begin 
			br_4_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_68_out) begin 
			br_4_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_4.br_4_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_88_out) begin 
			br_4_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_89_out) begin 
			br_4_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_5_happened_in_state_4.br_5_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_76_out) begin 
			br_5_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_77_out) begin 
			br_5_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_5_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_6_happened_in_state_4.br_6_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_79_out) begin 
			br_6_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_80_out) begin 
			br_6_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_6_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_7_happened_in_state_4.br_7_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_85_out) begin 
			br_7_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_86_out) begin 
			br_7_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_7_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_8_happened_in_state_1.br_8_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_49_out) begin 
			br_8_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_50_out) begin 
			br_8_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_8_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_9_happened_in_state_1.br_9_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_58_out) begin 
			br_9_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_59_out) begin 
			br_9_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_9_happened_in_state_1_in_data = 0;
		end
	end
	// controller for concat_162.concat_162_in0
	// controller for concat_162.concat_162_in1
	// Insensitive connections
	always @(*) begin
		concat_162_in0 = valid ? add_tmp_5 : add_tmp_5;
		concat_162_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for concat_163.concat_163_in0
	// controller for concat_163.concat_163_in1
	// Insensitive connections
	always @(*) begin
		concat_163_in0 = valid ? 32'd4 : 32'd4;
		concat_163_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_100.eq_100_in0
	// controller for eq_100.eq_100_in1
	// Insensitive connections
	always @(*) begin
		eq_100_in0 = valid ? 32'd3 : 32'd3;
		eq_100_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_102.eq_102_in0
	// controller for eq_102.eq_102_in1
	// Insensitive connections
	always @(*) begin
		eq_102_in0 = valid ? 32'd9 : 32'd9;
		eq_102_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_104.eq_104_in0
	// controller for eq_104.eq_104_in1
	// Insensitive connections
	always @(*) begin
		eq_104_in0 = valid ? 32'd10 : 32'd10;
		eq_104_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_105.eq_105_in0
	// controller for eq_105.eq_105_in1
	// Insensitive connections
	always @(*) begin
		eq_105_in0 = valid ? 32'd4 : 32'd4;
		eq_105_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_107.eq_107_in0
	// controller for eq_107.eq_107_in1
	// Insensitive connections
	always @(*) begin
		eq_107_in0 = valid ? 32'd10 : 32'd10;
		eq_107_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_108.eq_108_in0
	// controller for eq_108.eq_108_in1
	// Insensitive connections
	always @(*) begin
		eq_108_in0 = valid ? 32'd5 : 32'd5;
		eq_108_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_110.eq_110_in0
	// controller for eq_110.eq_110_in1
	// Insensitive connections
	always @(*) begin
		eq_110_in0 = valid ? 32'd6 : 32'd6;
		eq_110_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_112.eq_112_in0
	// controller for eq_112.eq_112_in1
	// Insensitive connections
	always @(*) begin
		eq_112_in0 = valid ? 32'd7 : 32'd7;
		eq_112_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_114.eq_114_in0
	// controller for eq_114.eq_114_in1
	// Insensitive connections
	always @(*) begin
		eq_114_in0 = valid ? 32'd4 : 32'd4;
		eq_114_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_115.eq_115_in0
	// controller for eq_115.eq_115_in1
	// Insensitive connections
	always @(*) begin
		eq_115_in0 = valid ? 32'd2 : 32'd2;
		eq_115_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_117.eq_117_in0
	// controller for eq_117.eq_117_in1
	// Insensitive connections
	always @(*) begin
		eq_117_in0 = valid ? 32'd1 : 32'd1;
		eq_117_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_119.eq_119_in0
	// controller for eq_119.eq_119_in1
	// Insensitive connections
	always @(*) begin
		eq_119_in0 = valid ? 32'd0 : 32'd0;
		eq_119_in1 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
	end
	// controller for eq_120.eq_120_in0
	// controller for eq_120.eq_120_in1
	// Insensitive connections
	always @(*) begin
		eq_120_in0 = valid ? 32'd8 : 32'd8;
		eq_120_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_123.eq_123_in0
	// controller for eq_123.eq_123_in1
	// Insensitive connections
	always @(*) begin
		eq_123_in0 = valid ? 32'd0 : 32'd0;
		eq_123_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_124.eq_124_in0
	// controller for eq_124.eq_124_in1
	// Insensitive connections
	always @(*) begin
		eq_124_in0 = valid ? 32'd3 : 32'd3;
		eq_124_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_127.eq_127_in0
	// controller for eq_127.eq_127_in1
	// Insensitive connections
	always @(*) begin
		eq_127_in0 = valid ? 32'd9 : 32'd9;
		eq_127_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_130.eq_130_in0
	// controller for eq_130.eq_130_in1
	// Insensitive connections
	always @(*) begin
		eq_130_in0 = valid ? 32'd10 : 32'd10;
		eq_130_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_131.eq_131_in0
	// controller for eq_131.eq_131_in1
	// Insensitive connections
	always @(*) begin
		eq_131_in0 = valid ? 32'd4 : 32'd4;
		eq_131_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_134.eq_134_in0
	// controller for eq_134.eq_134_in1
	// Insensitive connections
	always @(*) begin
		eq_134_in0 = valid ? 32'd10 : 32'd10;
		eq_134_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_135.eq_135_in0
	// controller for eq_135.eq_135_in1
	// Insensitive connections
	always @(*) begin
		eq_135_in0 = valid ? 32'd5 : 32'd5;
		eq_135_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_138.eq_138_in0
	// controller for eq_138.eq_138_in1
	// Insensitive connections
	always @(*) begin
		eq_138_in0 = valid ? 32'd6 : 32'd6;
		eq_138_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_141.eq_141_in0
	// controller for eq_141.eq_141_in1
	// Insensitive connections
	always @(*) begin
		eq_141_in0 = valid ? 32'd7 : 32'd7;
		eq_141_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_144.eq_144_in0
	// controller for eq_144.eq_144_in1
	// Insensitive connections
	always @(*) begin
		eq_144_in0 = valid ? 32'd4 : 32'd4;
		eq_144_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_145.eq_145_in0
	// controller for eq_145.eq_145_in1
	// Insensitive connections
	always @(*) begin
		eq_145_in0 = valid ? 32'd2 : 32'd2;
		eq_145_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_148.eq_148_in0
	// controller for eq_148.eq_148_in1
	// Insensitive connections
	always @(*) begin
		eq_148_in0 = valid ? 32'd1 : 32'd1;
		eq_148_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_166.eq_166_in0
	// controller for eq_166.eq_166_in1
	// Insensitive connections
	always @(*) begin
		eq_166_in0 = valid ? 32'd10 : 32'd10;
		eq_166_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_201.eq_201_in0
	// controller for eq_201.eq_201_in1
	// Insensitive connections
	always @(*) begin
		eq_201_in0 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
		eq_201_in1 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
	end
	// controller for eq_205.eq_205_in0
	// controller for eq_205.eq_205_in1
	// Insensitive connections
	always @(*) begin
		eq_205_in0 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
		eq_205_in1 = valid ? 32'd8 : 32'd8;
	end
	// controller for eq_207.eq_207_in0
	// controller for eq_207.eq_207_in1
	// Insensitive connections
	always @(*) begin
		eq_207_in0 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
		eq_207_in1 = valid ? 32'd9 : 32'd9;
	end
	// controller for eq_212.eq_212_in0
	// controller for eq_212.eq_212_in1
	// Insensitive connections
	always @(*) begin
		eq_212_in0 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
		eq_212_in1 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
	end
	// controller for eq_216.eq_216_in0
	// controller for eq_216.eq_216_in1
	// Insensitive connections
	always @(*) begin
		eq_216_in0 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
		eq_216_in1 = valid ? 32'd9 : 32'd9;
	end
	// controller for eq_221.eq_221_in0
	// controller for eq_221.eq_221_in1
	// Insensitive connections
	always @(*) begin
		eq_221_in0 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
		eq_221_in1 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
	end
	// controller for eq_225.eq_225_in0
	// controller for eq_225.eq_225_in1
	// Insensitive connections
	always @(*) begin
		eq_225_in0 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
		eq_225_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_227.eq_227_in0
	// controller for eq_227.eq_227_in1
	// Insensitive connections
	always @(*) begin
		eq_227_in0 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
		eq_227_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_232.eq_232_in0
	// controller for eq_232.eq_232_in1
	// Insensitive connections
	always @(*) begin
		eq_232_in0 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
		eq_232_in1 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
	end
	// controller for eq_236.eq_236_in0
	// controller for eq_236.eq_236_in1
	// Insensitive connections
	always @(*) begin
		eq_236_in0 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
		eq_236_in1 = valid ? 32'd10 : 32'd10;
	end
	// controller for eq_241.eq_241_in0
	// controller for eq_241.eq_241_in1
	// Insensitive connections
	always @(*) begin
		eq_241_in0 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
		eq_241_in1 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
	end
	// controller for eq_245.eq_245_in0
	// controller for eq_245.eq_245_in1
	// Insensitive connections
	always @(*) begin
		eq_245_in0 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
		eq_245_in1 = valid ? 32'd10 : 32'd10;
	end
	// controller for eq_250.eq_250_in0
	// controller for eq_250.eq_250_in1
	// Insensitive connections
	always @(*) begin
		eq_250_in0 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
		eq_250_in1 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
	end
	// controller for eq_254.eq_254_in0
	// controller for eq_254.eq_254_in1
	// Insensitive connections
	always @(*) begin
		eq_254_in0 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
		eq_254_in1 = valid ? 32'd10 : 32'd10;
	end
	// controller for eq_259.eq_259_in0
	// controller for eq_259.eq_259_in1
	// Insensitive connections
	always @(*) begin
		eq_259_in0 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
		eq_259_in1 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
	end
	// controller for eq_263.eq_263_in0
	// controller for eq_263.eq_263_in1
	// Insensitive connections
	always @(*) begin
		eq_263_in0 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
		eq_263_in1 = valid ? 32'd10 : 32'd10;
	end
	// controller for eq_268.eq_268_in0
	// controller for eq_268.eq_268_in1
	// Insensitive connections
	always @(*) begin
		eq_268_in0 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
		eq_268_in1 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
	end
	// controller for eq_272.eq_272_in0
	// controller for eq_272.eq_272_in1
	// Insensitive connections
	always @(*) begin
		eq_272_in0 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
		eq_272_in1 = valid ? 32'd6 : 32'd6;
	end
	// controller for eq_277.eq_277_in0
	// controller for eq_277.eq_277_in1
	// Insensitive connections
	always @(*) begin
		eq_277_in0 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
		eq_277_in1 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
	end
	// controller for eq_281.eq_281_in0
	// controller for eq_281.eq_281_in1
	// Insensitive connections
	always @(*) begin
		eq_281_in0 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
		eq_281_in1 = valid ? 32'd5 : 32'd5;
	end
	// controller for eq_283.eq_283_in0
	// controller for eq_283.eq_283_in1
	// Insensitive connections
	always @(*) begin
		eq_283_in0 = valid ? state_0_last_BB_reg : state_0_last_BB_reg;
		eq_283_in1 = valid ? 32'd6 : 32'd6;
	end
	// controller for eq_288.eq_288_in0
	// controller for eq_288.eq_288_in1
	// Insensitive connections
	always @(*) begin
		eq_288_in0 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
		eq_288_in1 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
	end
	// controller for eq_292.eq_292_in0
	// controller for eq_292.eq_292_in1
	// Insensitive connections
	always @(*) begin
		eq_292_in0 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
		eq_292_in1 = valid ? 32'd9 : 32'd9;
	end
	// controller for eq_297.eq_297_in0
	// controller for eq_297.eq_297_in1
	// Insensitive connections
	always @(*) begin
		eq_297_in0 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
		eq_297_in1 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
	end
	// controller for eq_301.eq_301_in0
	// controller for eq_301.eq_301_in1
	// Insensitive connections
	always @(*) begin
		eq_301_in0 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
		eq_301_in1 = valid ? 32'd9 : 32'd9;
	end
	// controller for eq_306.eq_306_in0
	// controller for eq_306.eq_306_in1
	// Insensitive connections
	always @(*) begin
		eq_306_in0 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
		eq_306_in1 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
	end
	// controller for eq_310.eq_310_in0
	// controller for eq_310.eq_310_in1
	// Insensitive connections
	always @(*) begin
		eq_310_in0 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
		eq_310_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_315.eq_315_in0
	// controller for eq_315.eq_315_in1
	// Insensitive connections
	always @(*) begin
		eq_315_in0 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
		eq_315_in1 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
	end
	// controller for eq_319.eq_319_in0
	// controller for eq_319.eq_319_in1
	// Insensitive connections
	always @(*) begin
		eq_319_in0 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
		eq_319_in1 = valid ? 32'd10 : 32'd10;
	end
	// controller for eq_324.eq_324_in0
	// controller for eq_324.eq_324_in1
	// Insensitive connections
	always @(*) begin
		eq_324_in0 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
		eq_324_in1 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
	end
	// controller for eq_328.eq_328_in0
	// controller for eq_328.eq_328_in1
	// Insensitive connections
	always @(*) begin
		eq_328_in0 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
		eq_328_in1 = valid ? 32'd10 : 32'd10;
	end
	// controller for eq_333.eq_333_in0
	// controller for eq_333.eq_333_in1
	// Insensitive connections
	always @(*) begin
		eq_333_in0 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
		eq_333_in1 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
	end
	// controller for eq_337.eq_337_in0
	// controller for eq_337.eq_337_in1
	// Insensitive connections
	always @(*) begin
		eq_337_in0 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
		eq_337_in1 = valid ? 32'd10 : 32'd10;
	end
	// controller for eq_342.eq_342_in0
	// controller for eq_342.eq_342_in1
	// Insensitive connections
	always @(*) begin
		eq_342_in0 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
		eq_342_in1 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
	end
	// controller for eq_346.eq_346_in0
	// controller for eq_346.eq_346_in1
	// Insensitive connections
	always @(*) begin
		eq_346_in0 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
		eq_346_in1 = valid ? 32'd10 : 32'd10;
	end
	// controller for eq_351.eq_351_in0
	// controller for eq_351.eq_351_in1
	// Insensitive connections
	always @(*) begin
		eq_351_in0 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
		eq_351_in1 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
	end
	// controller for eq_355.eq_355_in0
	// controller for eq_355.eq_355_in1
	// Insensitive connections
	always @(*) begin
		eq_355_in0 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
		eq_355_in1 = valid ? 32'd6 : 32'd6;
	end
	// controller for eq_360.eq_360_in0
	// controller for eq_360.eq_360_in1
	// Insensitive connections
	always @(*) begin
		eq_360_in0 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
		eq_360_in1 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
	end
	// controller for eq_364.eq_364_in0
	// controller for eq_364.eq_364_in1
	// Insensitive connections
	always @(*) begin
		eq_364_in0 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
		eq_364_in1 = valid ? 32'd5 : 32'd5;
	end
	// controller for eq_366.eq_366_in0
	// controller for eq_366.eq_366_in1
	// Insensitive connections
	always @(*) begin
		eq_366_in0 = valid ? state_1_last_BB_reg : state_1_last_BB_reg;
		eq_366_in1 = valid ? 32'd6 : 32'd6;
	end
	// controller for eq_371.eq_371_in0
	// controller for eq_371.eq_371_in1
	// Insensitive connections
	always @(*) begin
		eq_371_in0 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
		eq_371_in1 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
	end
	// controller for eq_375.eq_375_in0
	// controller for eq_375.eq_375_in1
	// Insensitive connections
	always @(*) begin
		eq_375_in0 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
		eq_375_in1 = valid ? 32'd8 : 32'd8;
	end
	// controller for eq_377.eq_377_in0
	// controller for eq_377.eq_377_in1
	// Insensitive connections
	always @(*) begin
		eq_377_in0 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
		eq_377_in1 = valid ? 32'd9 : 32'd9;
	end
	// controller for eq_382.eq_382_in0
	// controller for eq_382.eq_382_in1
	// Insensitive connections
	always @(*) begin
		eq_382_in0 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
		eq_382_in1 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
	end
	// controller for eq_386.eq_386_in0
	// controller for eq_386.eq_386_in1
	// Insensitive connections
	always @(*) begin
		eq_386_in0 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
		eq_386_in1 = valid ? 32'd9 : 32'd9;
	end
	// controller for eq_391.eq_391_in0
	// controller for eq_391.eq_391_in1
	// Insensitive connections
	always @(*) begin
		eq_391_in0 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
		eq_391_in1 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
	end
	// controller for eq_395.eq_395_in0
	// controller for eq_395.eq_395_in1
	// Insensitive connections
	always @(*) begin
		eq_395_in0 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
		eq_395_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_397.eq_397_in0
	// controller for eq_397.eq_397_in1
	// Insensitive connections
	always @(*) begin
		eq_397_in0 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
		eq_397_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_402.eq_402_in0
	// controller for eq_402.eq_402_in1
	// Insensitive connections
	always @(*) begin
		eq_402_in0 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
		eq_402_in1 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
	end
	// controller for eq_406.eq_406_in0
	// controller for eq_406.eq_406_in1
	// Insensitive connections
	always @(*) begin
		eq_406_in0 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
		eq_406_in1 = valid ? 32'd10 : 32'd10;
	end
	// controller for eq_411.eq_411_in0
	// controller for eq_411.eq_411_in1
	// Insensitive connections
	always @(*) begin
		eq_411_in0 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
		eq_411_in1 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
	end
	// controller for eq_415.eq_415_in0
	// controller for eq_415.eq_415_in1
	// Insensitive connections
	always @(*) begin
		eq_415_in0 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
		eq_415_in1 = valid ? 32'd10 : 32'd10;
	end
	// controller for eq_420.eq_420_in0
	// controller for eq_420.eq_420_in1
	// Insensitive connections
	always @(*) begin
		eq_420_in0 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
		eq_420_in1 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
	end
	// controller for eq_424.eq_424_in0
	// controller for eq_424.eq_424_in1
	// Insensitive connections
	always @(*) begin
		eq_424_in0 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
		eq_424_in1 = valid ? 32'd10 : 32'd10;
	end
	// controller for eq_429.eq_429_in0
	// controller for eq_429.eq_429_in1
	// Insensitive connections
	always @(*) begin
		eq_429_in0 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
		eq_429_in1 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
	end
	// controller for eq_433.eq_433_in0
	// controller for eq_433.eq_433_in1
	// Insensitive connections
	always @(*) begin
		eq_433_in0 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
		eq_433_in1 = valid ? 32'd10 : 32'd10;
	end
	// controller for eq_438.eq_438_in0
	// controller for eq_438.eq_438_in1
	// Insensitive connections
	always @(*) begin
		eq_438_in0 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
		eq_438_in1 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
	end
	// controller for eq_442.eq_442_in0
	// controller for eq_442.eq_442_in1
	// Insensitive connections
	always @(*) begin
		eq_442_in0 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
		eq_442_in1 = valid ? 32'd6 : 32'd6;
	end
	// controller for eq_447.eq_447_in0
	// controller for eq_447.eq_447_in1
	// Insensitive connections
	always @(*) begin
		eq_447_in0 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
		eq_447_in1 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
	end
	// controller for eq_451.eq_451_in0
	// controller for eq_451.eq_451_in1
	// Insensitive connections
	always @(*) begin
		eq_451_in0 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
		eq_451_in1 = valid ? 32'd5 : 32'd5;
	end
	// controller for eq_453.eq_453_in0
	// controller for eq_453.eq_453_in1
	// Insensitive connections
	always @(*) begin
		eq_453_in0 = valid ? state_2_last_BB_reg : state_2_last_BB_reg;
		eq_453_in1 = valid ? 32'd6 : 32'd6;
	end
	// controller for eq_458.eq_458_in0
	// controller for eq_458.eq_458_in1
	// Insensitive connections
	always @(*) begin
		eq_458_in0 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
		eq_458_in1 = valid ? state_3_last_BB_reg : state_3_last_BB_reg;
	end
	// controller for eq_462.eq_462_in0
	// controller for eq_462.eq_462_in1
	// Insensitive connections
	always @(*) begin
		eq_462_in0 = valid ? state_3_last_BB_reg : state_3_last_BB_reg;
		eq_462_in1 = valid ? 32'd8 : 32'd8;
	end
	// controller for eq_464.eq_464_in0
	// controller for eq_464.eq_464_in1
	// Insensitive connections
	always @(*) begin
		eq_464_in0 = valid ? state_3_last_BB_reg : state_3_last_BB_reg;
		eq_464_in1 = valid ? 32'd9 : 32'd9;
	end
	// controller for eq_469.eq_469_in0
	// controller for eq_469.eq_469_in1
	// Insensitive connections
	always @(*) begin
		eq_469_in0 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
		eq_469_in1 = valid ? state_3_last_BB_reg : state_3_last_BB_reg;
	end
	// controller for eq_473.eq_473_in0
	// controller for eq_473.eq_473_in1
	// Insensitive connections
	always @(*) begin
		eq_473_in0 = valid ? state_3_last_BB_reg : state_3_last_BB_reg;
		eq_473_in1 = valid ? 32'd9 : 32'd9;
	end
	// controller for eq_478.eq_478_in0
	// controller for eq_478.eq_478_in1
	// Insensitive connections
	always @(*) begin
		eq_478_in0 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
		eq_478_in1 = valid ? state_3_last_BB_reg : state_3_last_BB_reg;
	end
	// controller for eq_482.eq_482_in0
	// controller for eq_482.eq_482_in1
	// Insensitive connections
	always @(*) begin
		eq_482_in0 = valid ? state_3_last_BB_reg : state_3_last_BB_reg;
		eq_482_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_484.eq_484_in0
	// controller for eq_484.eq_484_in1
	// Insensitive connections
	always @(*) begin
		eq_484_in0 = valid ? state_3_last_BB_reg : state_3_last_BB_reg;
		eq_484_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_489.eq_489_in0
	// controller for eq_489.eq_489_in1
	// Insensitive connections
	always @(*) begin
		eq_489_in0 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
		eq_489_in1 = valid ? state_3_last_BB_reg : state_3_last_BB_reg;
	end
	// controller for eq_496.eq_496_in0
	// controller for eq_496.eq_496_in1
	// Insensitive connections
	always @(*) begin
		eq_496_in0 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
		eq_496_in1 = valid ? state_3_last_BB_reg : state_3_last_BB_reg;
	end
	// controller for eq_503.eq_503_in0
	// controller for eq_503.eq_503_in1
	// Insensitive connections
	always @(*) begin
		eq_503_in0 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
		eq_503_in1 = valid ? state_3_last_BB_reg : state_3_last_BB_reg;
	end
	// controller for eq_510.eq_510_in0
	// controller for eq_510.eq_510_in1
	// Insensitive connections
	always @(*) begin
		eq_510_in0 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
		eq_510_in1 = valid ? state_3_last_BB_reg : state_3_last_BB_reg;
	end
	// controller for eq_517.eq_517_in0
	// controller for eq_517.eq_517_in1
	// Insensitive connections
	always @(*) begin
		eq_517_in0 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
		eq_517_in1 = valid ? state_3_last_BB_reg : state_3_last_BB_reg;
	end
	// controller for eq_521.eq_521_in0
	// controller for eq_521.eq_521_in1
	// Insensitive connections
	always @(*) begin
		eq_521_in0 = valid ? state_3_last_BB_reg : state_3_last_BB_reg;
		eq_521_in1 = valid ? 32'd6 : 32'd6;
	end
	// controller for eq_526.eq_526_in0
	// controller for eq_526.eq_526_in1
	// Insensitive connections
	always @(*) begin
		eq_526_in0 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
		eq_526_in1 = valid ? state_3_last_BB_reg : state_3_last_BB_reg;
	end
	// controller for eq_530.eq_530_in0
	// controller for eq_530.eq_530_in1
	// Insensitive connections
	always @(*) begin
		eq_530_in0 = valid ? state_3_last_BB_reg : state_3_last_BB_reg;
		eq_530_in1 = valid ? 32'd5 : 32'd5;
	end
	// controller for eq_532.eq_532_in0
	// controller for eq_532.eq_532_in1
	// Insensitive connections
	always @(*) begin
		eq_532_in0 = valid ? state_3_last_BB_reg : state_3_last_BB_reg;
		eq_532_in1 = valid ? 32'd6 : 32'd6;
	end
	// controller for eq_537.eq_537_in0
	// controller for eq_537.eq_537_in1
	// Insensitive connections
	always @(*) begin
		eq_537_in0 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
		eq_537_in1 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
	end
	// controller for eq_541.eq_541_in0
	// controller for eq_541.eq_541_in1
	// Insensitive connections
	always @(*) begin
		eq_541_in0 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
		eq_541_in1 = valid ? 32'd8 : 32'd8;
	end
	// controller for eq_543.eq_543_in0
	// controller for eq_543.eq_543_in1
	// Insensitive connections
	always @(*) begin
		eq_543_in0 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
		eq_543_in1 = valid ? 32'd9 : 32'd9;
	end
	// controller for eq_548.eq_548_in0
	// controller for eq_548.eq_548_in1
	// Insensitive connections
	always @(*) begin
		eq_548_in0 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
		eq_548_in1 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
	end
	// controller for eq_552.eq_552_in0
	// controller for eq_552.eq_552_in1
	// Insensitive connections
	always @(*) begin
		eq_552_in0 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
		eq_552_in1 = valid ? 32'd9 : 32'd9;
	end
	// controller for eq_557.eq_557_in0
	// controller for eq_557.eq_557_in1
	// Insensitive connections
	always @(*) begin
		eq_557_in0 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
		eq_557_in1 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
	end
	// controller for eq_561.eq_561_in0
	// controller for eq_561.eq_561_in1
	// Insensitive connections
	always @(*) begin
		eq_561_in0 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
		eq_561_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_563.eq_563_in0
	// controller for eq_563.eq_563_in1
	// Insensitive connections
	always @(*) begin
		eq_563_in0 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
		eq_563_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_568.eq_568_in0
	// controller for eq_568.eq_568_in1
	// Insensitive connections
	always @(*) begin
		eq_568_in0 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
		eq_568_in1 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
	end
	// controller for eq_572.eq_572_in0
	// controller for eq_572.eq_572_in1
	// Insensitive connections
	always @(*) begin
		eq_572_in0 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
		eq_572_in1 = valid ? 32'd10 : 32'd10;
	end
	// controller for eq_577.eq_577_in0
	// controller for eq_577.eq_577_in1
	// Insensitive connections
	always @(*) begin
		eq_577_in0 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
		eq_577_in1 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
	end
	// controller for eq_581.eq_581_in0
	// controller for eq_581.eq_581_in1
	// Insensitive connections
	always @(*) begin
		eq_581_in0 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
		eq_581_in1 = valid ? 32'd10 : 32'd10;
	end
	// controller for eq_586.eq_586_in0
	// controller for eq_586.eq_586_in1
	// Insensitive connections
	always @(*) begin
		eq_586_in0 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
		eq_586_in1 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
	end
	// controller for eq_590.eq_590_in0
	// controller for eq_590.eq_590_in1
	// Insensitive connections
	always @(*) begin
		eq_590_in0 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
		eq_590_in1 = valid ? 32'd10 : 32'd10;
	end
	// controller for eq_595.eq_595_in0
	// controller for eq_595.eq_595_in1
	// Insensitive connections
	always @(*) begin
		eq_595_in0 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
		eq_595_in1 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
	end
	// controller for eq_599.eq_599_in0
	// controller for eq_599.eq_599_in1
	// Insensitive connections
	always @(*) begin
		eq_599_in0 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
		eq_599_in1 = valid ? 32'd10 : 32'd10;
	end
	// controller for eq_604.eq_604_in0
	// controller for eq_604.eq_604_in1
	// Insensitive connections
	always @(*) begin
		eq_604_in0 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
		eq_604_in1 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
	end
	// controller for eq_611.eq_611_in0
	// controller for eq_611.eq_611_in1
	// Insensitive connections
	always @(*) begin
		eq_611_in0 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
		eq_611_in1 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
	end
	// controller for eq_615.eq_615_in0
	// controller for eq_615.eq_615_in1
	// Insensitive connections
	always @(*) begin
		eq_615_in0 = valid ? state_4_last_BB_reg : state_4_last_BB_reg;
		eq_615_in1 = valid ? 32'd6 : 32'd6;
	end
	// controller for eq_96.eq_96_in0
	// controller for eq_96.eq_96_in1
	// Insensitive connections
	always @(*) begin
		eq_96_in0 = valid ? 32'd0 : 32'd0;
		eq_96_in1 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
	end
	// controller for eq_97.eq_97_in0
	// controller for eq_97.eq_97_in1
	// Insensitive connections
	always @(*) begin
		eq_97_in0 = valid ? 32'd8 : 32'd8;
		eq_97_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_99.eq_99_in0
	// controller for eq_99.eq_99_in1
	// Insensitive connections
	always @(*) begin
		eq_99_in0 = valid ? 32'd0 : 32'd0;
		eq_99_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for icmp_16.cmp_in0_icmp_16
	// controller for icmp_16.cmp_in1_icmp_16
	// Insensitive connections
	always @(*) begin
		cmp_in0_icmp_16 = valid ? add_out_add_15 : add_out_add_15;
		cmp_in1_icmp_16 = valid ? 32'd4 : 32'd4;
	end
	// controller for in.in_read_valid_reg
	always @(*) begin
		if (andOp_159_out) begin 
			in_read_valid_reg = -(1'd1);
		end else begin
			in_read_valid_reg = 0;
		end
	end
	// controller for notOp_121.notOp_121_in0
	// Insensitive connections
	always @(*) begin
		notOp_121_in0 = valid ? eq_120_out : eq_120_out;
	end
	// controller for notOp_125.notOp_125_in0
	// Insensitive connections
	always @(*) begin
		notOp_125_in0 = valid ? eq_124_out : eq_124_out;
	end
	// controller for notOp_128.notOp_128_in0
	// Insensitive connections
	always @(*) begin
		notOp_128_in0 = valid ? eq_127_out : eq_127_out;
	end
	// controller for notOp_132.notOp_132_in0
	// Insensitive connections
	always @(*) begin
		notOp_132_in0 = valid ? eq_131_out : eq_131_out;
	end
	// controller for notOp_136.notOp_136_in0
	// Insensitive connections
	always @(*) begin
		notOp_136_in0 = valid ? eq_135_out : eq_135_out;
	end
	// controller for notOp_139.notOp_139_in0
	// Insensitive connections
	always @(*) begin
		notOp_139_in0 = valid ? eq_138_out : eq_138_out;
	end
	// controller for notOp_142.notOp_142_in0
	// Insensitive connections
	always @(*) begin
		notOp_142_in0 = valid ? eq_141_out : eq_141_out;
	end
	// controller for notOp_146.notOp_146_in0
	// Insensitive connections
	always @(*) begin
		notOp_146_in0 = valid ? eq_145_out : eq_145_out;
	end
	// controller for notOp_149.notOp_149_in0
	// Insensitive connections
	always @(*) begin
		notOp_149_in0 = valid ? eq_148_out : eq_148_out;
	end
	// controller for notOp_178.notOp_178_in0
	// Insensitive connections
	always @(*) begin
		notOp_178_in0 = valid ? andOp_174_out : andOp_174_out;
	end
	// controller for notOp_180.notOp_180_in0
	// Insensitive connections
	always @(*) begin
		notOp_180_in0 = valid ? andOp_62_out : andOp_62_out;
	end
	// controller for notOp_182.notOp_182_in0
	// Insensitive connections
	always @(*) begin
		notOp_182_in0 = valid ? andOp_71_out : andOp_71_out;
	end
	// controller for notOp_184.notOp_184_in0
	// Insensitive connections
	always @(*) begin
		notOp_184_in0 = valid ? andOp_60_out : andOp_60_out;
	end
	// controller for notOp_186.notOp_186_in0
	// Insensitive connections
	always @(*) begin
		notOp_186_in0 = valid ? andOp_175_out : andOp_175_out;
	end
	// controller for notOp_188.notOp_188_in0
	// Insensitive connections
	always @(*) begin
		notOp_188_in0 = valid ? andOp_176_out : andOp_176_out;
	end
	// controller for notOp_190.notOp_190_in0
	// Insensitive connections
	always @(*) begin
		notOp_190_in0 = valid ? andOp_177_out : andOp_177_out;
	end
	// controller for notOp_192.notOp_192_in0
	// Insensitive connections
	always @(*) begin
		notOp_192_in0 = valid ? andOp_83_out : andOp_83_out;
	end
	// controller for notOp_198.notOp_198_in0
	// Insensitive connections
	always @(*) begin
		notOp_198_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_203.notOp_203_in0
	// Insensitive connections
	always @(*) begin
		notOp_203_in0 = valid ? eq_201_out : eq_201_out;
	end
	// controller for notOp_209.notOp_209_in0
	// Insensitive connections
	always @(*) begin
		notOp_209_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_214.notOp_214_in0
	// Insensitive connections
	always @(*) begin
		notOp_214_in0 = valid ? eq_212_out : eq_212_out;
	end
	// controller for notOp_218.notOp_218_in0
	// Insensitive connections
	always @(*) begin
		notOp_218_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_223.notOp_223_in0
	// Insensitive connections
	always @(*) begin
		notOp_223_in0 = valid ? eq_221_out : eq_221_out;
	end
	// controller for notOp_229.notOp_229_in0
	// Insensitive connections
	always @(*) begin
		notOp_229_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_234.notOp_234_in0
	// Insensitive connections
	always @(*) begin
		notOp_234_in0 = valid ? eq_232_out : eq_232_out;
	end
	// controller for notOp_238.notOp_238_in0
	// Insensitive connections
	always @(*) begin
		notOp_238_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_243.notOp_243_in0
	// Insensitive connections
	always @(*) begin
		notOp_243_in0 = valid ? eq_241_out : eq_241_out;
	end
	// controller for notOp_247.notOp_247_in0
	// Insensitive connections
	always @(*) begin
		notOp_247_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_252.notOp_252_in0
	// Insensitive connections
	always @(*) begin
		notOp_252_in0 = valid ? eq_250_out : eq_250_out;
	end
	// controller for notOp_256.notOp_256_in0
	// Insensitive connections
	always @(*) begin
		notOp_256_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_261.notOp_261_in0
	// Insensitive connections
	always @(*) begin
		notOp_261_in0 = valid ? eq_259_out : eq_259_out;
	end
	// controller for notOp_265.notOp_265_in0
	// Insensitive connections
	always @(*) begin
		notOp_265_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_270.notOp_270_in0
	// Insensitive connections
	always @(*) begin
		notOp_270_in0 = valid ? eq_268_out : eq_268_out;
	end
	// controller for notOp_274.notOp_274_in0
	// Insensitive connections
	always @(*) begin
		notOp_274_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_279.notOp_279_in0
	// Insensitive connections
	always @(*) begin
		notOp_279_in0 = valid ? eq_277_out : eq_277_out;
	end
	// controller for notOp_285.notOp_285_in0
	// Insensitive connections
	always @(*) begin
		notOp_285_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
	end
	// controller for notOp_290.notOp_290_in0
	// Insensitive connections
	always @(*) begin
		notOp_290_in0 = valid ? eq_288_out : eq_288_out;
	end
	// controller for notOp_294.notOp_294_in0
	// Insensitive connections
	always @(*) begin
		notOp_294_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_299.notOp_299_in0
	// Insensitive connections
	always @(*) begin
		notOp_299_in0 = valid ? eq_297_out : eq_297_out;
	end
	// controller for notOp_303.notOp_303_in0
	// Insensitive connections
	always @(*) begin
		notOp_303_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
	end
	// controller for notOp_308.notOp_308_in0
	// Insensitive connections
	always @(*) begin
		notOp_308_in0 = valid ? eq_306_out : eq_306_out;
	end
	// controller for notOp_312.notOp_312_in0
	// Insensitive connections
	always @(*) begin
		notOp_312_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_317.notOp_317_in0
	// Insensitive connections
	always @(*) begin
		notOp_317_in0 = valid ? eq_315_out : eq_315_out;
	end
	// controller for notOp_321.notOp_321_in0
	// Insensitive connections
	always @(*) begin
		notOp_321_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_326.notOp_326_in0
	// Insensitive connections
	always @(*) begin
		notOp_326_in0 = valid ? eq_324_out : eq_324_out;
	end
	// controller for notOp_330.notOp_330_in0
	// Insensitive connections
	always @(*) begin
		notOp_330_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_335.notOp_335_in0
	// Insensitive connections
	always @(*) begin
		notOp_335_in0 = valid ? eq_333_out : eq_333_out;
	end
	// controller for notOp_339.notOp_339_in0
	// Insensitive connections
	always @(*) begin
		notOp_339_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_344.notOp_344_in0
	// Insensitive connections
	always @(*) begin
		notOp_344_in0 = valid ? eq_342_out : eq_342_out;
	end
	// controller for notOp_348.notOp_348_in0
	// Insensitive connections
	always @(*) begin
		notOp_348_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_353.notOp_353_in0
	// Insensitive connections
	always @(*) begin
		notOp_353_in0 = valid ? eq_351_out : eq_351_out;
	end
	// controller for notOp_357.notOp_357_in0
	// Insensitive connections
	always @(*) begin
		notOp_357_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_362.notOp_362_in0
	// Insensitive connections
	always @(*) begin
		notOp_362_in0 = valid ? eq_360_out : eq_360_out;
	end
	// controller for notOp_368.notOp_368_in0
	// Insensitive connections
	always @(*) begin
		notOp_368_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_373.notOp_373_in0
	// Insensitive connections
	always @(*) begin
		notOp_373_in0 = valid ? eq_371_out : eq_371_out;
	end
	// controller for notOp_379.notOp_379_in0
	// Insensitive connections
	always @(*) begin
		notOp_379_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
	end
	// controller for notOp_384.notOp_384_in0
	// Insensitive connections
	always @(*) begin
		notOp_384_in0 = valid ? eq_382_out : eq_382_out;
	end
	// controller for notOp_388.notOp_388_in0
	// Insensitive connections
	always @(*) begin
		notOp_388_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_393.notOp_393_in0
	// Insensitive connections
	always @(*) begin
		notOp_393_in0 = valid ? eq_391_out : eq_391_out;
	end
	// controller for notOp_399.notOp_399_in0
	// Insensitive connections
	always @(*) begin
		notOp_399_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_404.notOp_404_in0
	// Insensitive connections
	always @(*) begin
		notOp_404_in0 = valid ? eq_402_out : eq_402_out;
	end
	// controller for notOp_408.notOp_408_in0
	// Insensitive connections
	always @(*) begin
		notOp_408_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_413.notOp_413_in0
	// Insensitive connections
	always @(*) begin
		notOp_413_in0 = valid ? eq_411_out : eq_411_out;
	end
	// controller for notOp_417.notOp_417_in0
	// Insensitive connections
	always @(*) begin
		notOp_417_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_422.notOp_422_in0
	// Insensitive connections
	always @(*) begin
		notOp_422_in0 = valid ? eq_420_out : eq_420_out;
	end
	// controller for notOp_426.notOp_426_in0
	// Insensitive connections
	always @(*) begin
		notOp_426_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_431.notOp_431_in0
	// Insensitive connections
	always @(*) begin
		notOp_431_in0 = valid ? eq_429_out : eq_429_out;
	end
	// controller for notOp_435.notOp_435_in0
	// Insensitive connections
	always @(*) begin
		notOp_435_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_440.notOp_440_in0
	// Insensitive connections
	always @(*) begin
		notOp_440_in0 = valid ? eq_438_out : eq_438_out;
	end
	// controller for notOp_444.notOp_444_in0
	// Insensitive connections
	always @(*) begin
		notOp_444_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_449.notOp_449_in0
	// Insensitive connections
	always @(*) begin
		notOp_449_in0 = valid ? eq_447_out : eq_447_out;
	end
	// controller for notOp_455.notOp_455_in0
	// Insensitive connections
	always @(*) begin
		notOp_455_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_460.notOp_460_in0
	// Insensitive connections
	always @(*) begin
		notOp_460_in0 = valid ? eq_458_out : eq_458_out;
	end
	// controller for notOp_466.notOp_466_in0
	// Insensitive connections
	always @(*) begin
		notOp_466_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
	end
	// controller for notOp_47.notOp_47_in0
	// Insensitive connections
	always @(*) begin
		notOp_47_in0 = valid ? andOp_46_out : andOp_46_out;
	end
	// controller for notOp_471.notOp_471_in0
	// Insensitive connections
	always @(*) begin
		notOp_471_in0 = valid ? eq_469_out : eq_469_out;
	end
	// controller for notOp_475.notOp_475_in0
	// Insensitive connections
	always @(*) begin
		notOp_475_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_480.notOp_480_in0
	// Insensitive connections
	always @(*) begin
		notOp_480_in0 = valid ? eq_478_out : eq_478_out;
	end
	// controller for notOp_486.notOp_486_in0
	// Insensitive connections
	always @(*) begin
		notOp_486_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
	end
	// controller for notOp_491.notOp_491_in0
	// Insensitive connections
	always @(*) begin
		notOp_491_in0 = valid ? eq_489_out : eq_489_out;
	end
	// controller for notOp_493.notOp_493_in0
	// Insensitive connections
	always @(*) begin
		notOp_493_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
	end
	// controller for notOp_498.notOp_498_in0
	// Insensitive connections
	always @(*) begin
		notOp_498_in0 = valid ? eq_496_out : eq_496_out;
	end
	// controller for notOp_50.notOp_50_in0
	// Insensitive connections
	always @(*) begin
		notOp_50_in0 = valid ? andOp_49_out : andOp_49_out;
	end
	// controller for notOp_500.notOp_500_in0
	// Insensitive connections
	always @(*) begin
		notOp_500_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
	end
	// controller for notOp_505.notOp_505_in0
	// Insensitive connections
	always @(*) begin
		notOp_505_in0 = valid ? eq_503_out : eq_503_out;
	end
	// controller for notOp_507.notOp_507_in0
	// Insensitive connections
	always @(*) begin
		notOp_507_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
	end
	// controller for notOp_512.notOp_512_in0
	// Insensitive connections
	always @(*) begin
		notOp_512_in0 = valid ? eq_510_out : eq_510_out;
	end
	// controller for notOp_514.notOp_514_in0
	// Insensitive connections
	always @(*) begin
		notOp_514_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_519.notOp_519_in0
	// Insensitive connections
	always @(*) begin
		notOp_519_in0 = valid ? eq_517_out : eq_517_out;
	end
	// controller for notOp_523.notOp_523_in0
	// Insensitive connections
	always @(*) begin
		notOp_523_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_528.notOp_528_in0
	// Insensitive connections
	always @(*) begin
		notOp_528_in0 = valid ? eq_526_out : eq_526_out;
	end
	// controller for notOp_53.notOp_53_in0
	// Insensitive connections
	always @(*) begin
		notOp_53_in0 = valid ? andOp_52_out : andOp_52_out;
	end
	// controller for notOp_534.notOp_534_in0
	// Insensitive connections
	always @(*) begin
		notOp_534_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_539.notOp_539_in0
	// Insensitive connections
	always @(*) begin
		notOp_539_in0 = valid ? eq_537_out : eq_537_out;
	end
	// controller for notOp_545.notOp_545_in0
	// Insensitive connections
	always @(*) begin
		notOp_545_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_550.notOp_550_in0
	// Insensitive connections
	always @(*) begin
		notOp_550_in0 = valid ? eq_548_out : eq_548_out;
	end
	// controller for notOp_554.notOp_554_in0
	// Insensitive connections
	always @(*) begin
		notOp_554_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_559.notOp_559_in0
	// Insensitive connections
	always @(*) begin
		notOp_559_in0 = valid ? eq_557_out : eq_557_out;
	end
	// controller for notOp_56.notOp_56_in0
	// Insensitive connections
	always @(*) begin
		notOp_56_in0 = valid ? andOp_55_out : andOp_55_out;
	end
	// controller for notOp_565.notOp_565_in0
	// Insensitive connections
	always @(*) begin
		notOp_565_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
	end
	// controller for notOp_570.notOp_570_in0
	// Insensitive connections
	always @(*) begin
		notOp_570_in0 = valid ? eq_568_out : eq_568_out;
	end
	// controller for notOp_574.notOp_574_in0
	// Insensitive connections
	always @(*) begin
		notOp_574_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
	end
	// controller for notOp_579.notOp_579_in0
	// Insensitive connections
	always @(*) begin
		notOp_579_in0 = valid ? eq_577_out : eq_577_out;
	end
	// controller for notOp_583.notOp_583_in0
	// Insensitive connections
	always @(*) begin
		notOp_583_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
	end
	// controller for notOp_588.notOp_588_in0
	// Insensitive connections
	always @(*) begin
		notOp_588_in0 = valid ? eq_586_out : eq_586_out;
	end
	// controller for notOp_59.notOp_59_in0
	// Insensitive connections
	always @(*) begin
		notOp_59_in0 = valid ? andOp_58_out : andOp_58_out;
	end
	// controller for notOp_592.notOp_592_in0
	// Insensitive connections
	always @(*) begin
		notOp_592_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
	end
	// controller for notOp_597.notOp_597_in0
	// Insensitive connections
	always @(*) begin
		notOp_597_in0 = valid ? eq_595_out : eq_595_out;
	end
	// controller for notOp_601.notOp_601_in0
	// Insensitive connections
	always @(*) begin
		notOp_601_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
	end
	// controller for notOp_606.notOp_606_in0
	// Insensitive connections
	always @(*) begin
		notOp_606_in0 = valid ? eq_604_out : eq_604_out;
	end
	// controller for notOp_608.notOp_608_in0
	// Insensitive connections
	always @(*) begin
		notOp_608_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
	end
	// controller for notOp_61.notOp_61_in0
	// Insensitive connections
	always @(*) begin
		notOp_61_in0 = valid ? in_read_ready : in_read_ready;
	end
	// controller for notOp_613.notOp_613_in0
	// Insensitive connections
	always @(*) begin
		notOp_613_in0 = valid ? eq_611_out : eq_611_out;
	end
	// controller for notOp_65.notOp_65_in0
	// Insensitive connections
	always @(*) begin
		notOp_65_in0 = valid ? andOp_64_out : andOp_64_out;
	end
	// controller for notOp_68.notOp_68_in0
	// Insensitive connections
	always @(*) begin
		notOp_68_in0 = valid ? andOp_67_out : andOp_67_out;
	end
	// controller for notOp_70.notOp_70_in0
	// Insensitive connections
	always @(*) begin
		notOp_70_in0 = valid ? icmp_tmp_6 : icmp_tmp_6;
	end
	// controller for notOp_74.notOp_74_in0
	// Insensitive connections
	always @(*) begin
		notOp_74_in0 = valid ? andOp_73_out : andOp_73_out;
	end
	// controller for notOp_77.notOp_77_in0
	// Insensitive connections
	always @(*) begin
		notOp_77_in0 = valid ? andOp_76_out : andOp_76_out;
	end
	// controller for notOp_80.notOp_80_in0
	// Insensitive connections
	always @(*) begin
		notOp_80_in0 = valid ? andOp_79_out : andOp_79_out;
	end
	// controller for notOp_82.notOp_82_in0
	// Insensitive connections
	always @(*) begin
		notOp_82_in0 = valid ? out_write_ready : out_write_ready;
	end
	// controller for notOp_86.notOp_86_in0
	// Insensitive connections
	always @(*) begin
		notOp_86_in0 = valid ? andOp_85_out : andOp_85_out;
	end
	// controller for notOp_89.notOp_89_in0
	// Insensitive connections
	always @(*) begin
		notOp_89_in0 = valid ? andOp_88_out : andOp_88_out;
	end
	// controller for notOp_91.notOp_91_in0
	// Insensitive connections
	always @(*) begin
		notOp_91_in0 = valid ? icmp_tmp_6 : icmp_tmp_6;
	end
	// controller for notOp_95.notOp_95_in0
	// Insensitive connections
	always @(*) begin
		notOp_95_in0 = valid ? andOp_94_out : andOp_94_out;
	end
	// controller for orOp_101.orOp_101_in0
	// controller for orOp_101.orOp_101_in1
	// Insensitive connections
	always @(*) begin
		orOp_101_in0 = valid ? eq_100_out : eq_100_out;
		orOp_101_in1 = valid ? andOp_46_out : andOp_46_out;
	end
	// controller for orOp_103.orOp_103_in0
	// controller for orOp_103.orOp_103_in1
	// Insensitive connections
	always @(*) begin
		orOp_103_in0 = valid ? eq_102_out : eq_102_out;
		orOp_103_in1 = valid ? andOp_49_out : andOp_49_out;
	end
	// controller for orOp_106.orOp_106_in0
	// controller for orOp_106.orOp_106_in1
	// Insensitive connections
	always @(*) begin
		orOp_106_in0 = valid ? eq_105_out : eq_105_out;
		orOp_106_in1 = valid ? andOp_64_out : andOp_64_out;
	end
	// controller for orOp_109.orOp_109_in0
	// controller for orOp_109.orOp_109_in1
	// Insensitive connections
	always @(*) begin
		orOp_109_in0 = valid ? eq_108_out : eq_108_out;
		orOp_109_in1 = valid ? andOp_94_out : andOp_94_out;
	end
	// controller for orOp_111.orOp_111_in0
	// controller for orOp_111.orOp_111_in1
	// Insensitive connections
	always @(*) begin
		orOp_111_in0 = valid ? eq_110_out : eq_110_out;
		orOp_111_in1 = valid ? andOp_76_out : andOp_76_out;
	end
	// controller for orOp_113.orOp_113_in0
	// controller for orOp_113.orOp_113_in1
	// Insensitive connections
	always @(*) begin
		orOp_113_in0 = valid ? eq_112_out : eq_112_out;
		orOp_113_in1 = valid ? andOp_81_out : andOp_81_out;
	end
	// controller for orOp_116.orOp_116_in0
	// controller for orOp_116.orOp_116_in1
	// Insensitive connections
	always @(*) begin
		orOp_116_in0 = valid ? eq_115_out : eq_115_out;
		orOp_116_in1 = valid ? andOp_85_out : andOp_85_out;
	end
	// controller for orOp_118.orOp_118_in0
	// controller for orOp_118.orOp_118_in1
	// Insensitive connections
	always @(*) begin
		orOp_118_in0 = valid ? eq_117_out : eq_117_out;
		orOp_118_in1 = valid ? andOp_69_out : andOp_69_out;
	end
	// controller for orOp_98.orOp_98_in0
	// controller for orOp_98.orOp_98_in1
	// Insensitive connections
	always @(*) begin
		orOp_98_in0 = valid ? eq_97_out : eq_97_out;
		orOp_98_in1 = valid ? andOp_55_out : andOp_55_out;
	end
	// controller for out.out_in_data_reg
	always @(*) begin
		if (andOp_171_out) begin 
			out_in_data_reg = rdata_ram_0;
		end else begin
			out_in_data_reg = 0;
		end
	end
	// controller for out.out_write_valid_reg
	always @(*) begin
		if (andOp_172_out) begin 
			out_write_valid_reg = -(1'd1);
		end else begin
			out_write_valid_reg = 0;
		end
	end
	// controller for phi_7.phi_in_phi_7
	// controller for phi_7.phi_last_block_phi_7
	// controller for phi_7.phi_s_phi_7
	// Insensitive connections
	always @(*) begin
		phi_in_phi_7 = valid ? concat_162_out : concat_162_out;
		phi_last_block_phi_7 = valid ? bb_3_predecessor_in_state_1_out_data : bb_3_predecessor_in_state_1_out_data;
		phi_s_phi_7 = valid ? concat_163_out : concat_163_out;
	end
	// controller for ram_0.raddr_ram_0_reg
	always @(*) begin
		if (andOp_155_out) begin 
			raddr_ram_0_reg = 32'd0;
		end else if (andOp_157_out) begin 
			raddr_ram_0_reg = 32'd0;
		end else begin
			raddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.waddr_ram_0_reg
	always @(*) begin
		if (andOp_154_out) begin 
			waddr_ram_0_reg = 32'd0;
		end else if (andOp_156_out) begin 
			waddr_ram_0_reg = 32'd0;
		end else begin
			waddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wdata_ram_0_reg
	always @(*) begin
		if (andOp_154_out) begin 
			wdata_ram_0_reg = 32'd0;
		end else if (andOp_156_out) begin 
			wdata_ram_0_reg = add_out_add_13;
		end else begin
			wdata_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wen_ram_0_reg
	always @(*) begin
		if (andOp_154_out) begin 
			wen_ram_0_reg = 1'd1;
		end else if (andOp_156_out) begin 
			wen_ram_0_reg = 1'd1;
		end else begin
			wen_ram_0_reg = 0;
		end
	end
	// controller for ret_21.valid_reg
	always @(*) begin
		if (andOp_170_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// controller for tmp_output_165.tmp_output_165_in_data
	always @(*) begin
		if (eq_166_out) begin 
			tmp_output_165_in_data = in_out_data;
		end else begin
			tmp_output_165_in_data = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			add_tmp_5 <= 0;
		end else begin
			if (andOp_196_out) begin
				add_tmp_5 <= add_out_add_15;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			call_tmp_2 <= 0;
		end else begin
			if (andOp_195_out) begin
				call_tmp_2 <= in_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_0 <= 0;
		end else begin
			if (andOp_200_out) begin
				data_store_0_0 <= in_read_ready;
			end
			if (andOp_206_out) begin
				data_store_0_0 <= data_store_1_9;
			end
			if (andOp_208_out) begin
				data_store_0_0 <= data_store_1_9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_1 <= 0;
		end else begin
			if (andOp_211_out) begin
				data_store_0_1 <= in_out_data;
			end
			if (andOp_217_out) begin
				data_store_0_1 <= data_store_1_10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_2 <= 0;
		end else begin
			if (andOp_220_out) begin
				data_store_0_2 <= phi_out_phi_7;
			end
			if (andOp_226_out) begin
				data_store_0_2 <= data_store_4_38;
			end
			if (andOp_228_out) begin
				data_store_0_2 <= data_store_1_11;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_3 <= 0;
		end else begin
			if (andOp_231_out) begin
				data_store_0_3 <= rdata_ram_0;
			end
			if (andOp_237_out) begin
				data_store_0_3 <= data_store_3_30;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_4 <= 0;
		end else begin
			if (andOp_240_out) begin
				data_store_0_4 <= add_out_add_13;
			end
			if (andOp_246_out) begin
				data_store_0_4 <= data_store_3_31;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_5 <= 0;
		end else begin
			if (andOp_249_out) begin
				data_store_0_5 <= add_out_add_15;
			end
			if (andOp_255_out) begin
				data_store_0_5 <= data_store_3_32;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_6 <= 0;
		end else begin
			if (andOp_258_out) begin
				data_store_0_6 <= cmp_out_icmp_16;
			end
			if (andOp_264_out) begin
				data_store_0_6 <= data_store_3_33;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_7 <= 0;
		end else begin
			if (andOp_267_out) begin
				data_store_0_7 <= rdata_ram_0;
			end
			if (andOp_273_out) begin
				data_store_0_7 <= data_store_4_43;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_8 <= 0;
		end else begin
			if (andOp_276_out) begin
				data_store_0_8 <= out_write_ready;
			end
			if (andOp_282_out) begin
				data_store_0_8 <= data_store_4_44;
			end
			if (andOp_284_out) begin
				data_store_0_8 <= data_store_4_44;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_10 <= 0;
		end else begin
			if (andOp_296_out) begin
				data_store_1_10 <= in_out_data;
			end
			if (andOp_298_out) begin
				data_store_1_10 <= data_store_0_1;
			end
			if (andOp_302_out) begin
				data_store_1_10 <= data_store_1_10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_11 <= 0;
		end else begin
			if (andOp_305_out) begin
				data_store_1_11 <= phi_out_phi_7;
			end
			if (andOp_307_out) begin
				data_store_1_11 <= data_store_0_2;
			end
			if (andOp_311_out) begin
				data_store_1_11 <= data_store_4_38;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_12 <= 0;
		end else begin
			if (andOp_314_out) begin
				data_store_1_12 <= rdata_ram_0;
			end
			if (andOp_316_out) begin
				data_store_1_12 <= data_store_0_3;
			end
			if (andOp_320_out) begin
				data_store_1_12 <= data_store_3_30;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_13 <= 0;
		end else begin
			if (andOp_323_out) begin
				data_store_1_13 <= add_out_add_13;
			end
			if (andOp_325_out) begin
				data_store_1_13 <= data_store_0_4;
			end
			if (andOp_329_out) begin
				data_store_1_13 <= data_store_3_31;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_14 <= 0;
		end else begin
			if (andOp_332_out) begin
				data_store_1_14 <= add_out_add_15;
			end
			if (andOp_334_out) begin
				data_store_1_14 <= data_store_0_5;
			end
			if (andOp_338_out) begin
				data_store_1_14 <= data_store_3_32;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_15 <= 0;
		end else begin
			if (andOp_341_out) begin
				data_store_1_15 <= cmp_out_icmp_16;
			end
			if (andOp_343_out) begin
				data_store_1_15 <= data_store_0_6;
			end
			if (andOp_347_out) begin
				data_store_1_15 <= data_store_3_33;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_16 <= 0;
		end else begin
			if (andOp_350_out) begin
				data_store_1_16 <= rdata_ram_0;
			end
			if (andOp_352_out) begin
				data_store_1_16 <= data_store_0_7;
			end
			if (andOp_356_out) begin
				data_store_1_16 <= data_store_4_43;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_17 <= 0;
		end else begin
			if (andOp_359_out) begin
				data_store_1_17 <= out_write_ready;
			end
			if (andOp_361_out) begin
				data_store_1_17 <= data_store_0_8;
			end
			if (andOp_365_out) begin
				data_store_1_17 <= data_store_4_44;
			end
			if (andOp_367_out) begin
				data_store_1_17 <= data_store_4_44;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_9 <= 0;
		end else begin
			if (andOp_287_out) begin
				data_store_1_9 <= in_read_ready;
			end
			if (andOp_289_out) begin
				data_store_1_9 <= data_store_0_0;
			end
			if (andOp_293_out) begin
				data_store_1_9 <= data_store_1_9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_18 <= 0;
		end else begin
			if (andOp_370_out) begin
				data_store_2_18 <= in_read_ready;
			end
			if (andOp_372_out) begin
				data_store_2_18 <= data_store_1_9;
			end
			if (andOp_376_out) begin
				data_store_2_18 <= data_store_1_9;
			end
			if (andOp_378_out) begin
				data_store_2_18 <= data_store_1_9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_19 <= 0;
		end else begin
			if (andOp_381_out) begin
				data_store_2_19 <= in_out_data;
			end
			if (andOp_383_out) begin
				data_store_2_19 <= data_store_1_10;
			end
			if (andOp_387_out) begin
				data_store_2_19 <= data_store_1_10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_20 <= 0;
		end else begin
			if (andOp_390_out) begin
				data_store_2_20 <= phi_out_phi_7;
			end
			if (andOp_392_out) begin
				data_store_2_20 <= data_store_1_11;
			end
			if (andOp_396_out) begin
				data_store_2_20 <= data_store_4_38;
			end
			if (andOp_398_out) begin
				data_store_2_20 <= data_store_1_11;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_21 <= 0;
		end else begin
			if (andOp_401_out) begin
				data_store_2_21 <= rdata_ram_0;
			end
			if (andOp_403_out) begin
				data_store_2_21 <= data_store_1_12;
			end
			if (andOp_407_out) begin
				data_store_2_21 <= data_store_3_30;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_22 <= 0;
		end else begin
			if (andOp_410_out) begin
				data_store_2_22 <= add_out_add_13;
			end
			if (andOp_412_out) begin
				data_store_2_22 <= data_store_1_13;
			end
			if (andOp_416_out) begin
				data_store_2_22 <= data_store_3_31;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_23 <= 0;
		end else begin
			if (andOp_419_out) begin
				data_store_2_23 <= add_out_add_15;
			end
			if (andOp_421_out) begin
				data_store_2_23 <= data_store_1_14;
			end
			if (andOp_425_out) begin
				data_store_2_23 <= data_store_3_32;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_24 <= 0;
		end else begin
			if (andOp_428_out) begin
				data_store_2_24 <= cmp_out_icmp_16;
			end
			if (andOp_430_out) begin
				data_store_2_24 <= data_store_1_15;
			end
			if (andOp_434_out) begin
				data_store_2_24 <= data_store_3_33;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_25 <= 0;
		end else begin
			if (andOp_437_out) begin
				data_store_2_25 <= rdata_ram_0;
			end
			if (andOp_439_out) begin
				data_store_2_25 <= data_store_1_16;
			end
			if (andOp_443_out) begin
				data_store_2_25 <= data_store_4_43;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_26 <= 0;
		end else begin
			if (andOp_446_out) begin
				data_store_2_26 <= out_write_ready;
			end
			if (andOp_448_out) begin
				data_store_2_26 <= data_store_1_17;
			end
			if (andOp_452_out) begin
				data_store_2_26 <= data_store_4_44;
			end
			if (andOp_454_out) begin
				data_store_2_26 <= data_store_4_44;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_27 <= 0;
		end else begin
			if (andOp_457_out) begin
				data_store_3_27 <= in_read_ready;
			end
			if (andOp_459_out) begin
				data_store_3_27 <= data_store_2_18;
			end
			if (andOp_463_out) begin
				data_store_3_27 <= data_store_1_9;
			end
			if (andOp_465_out) begin
				data_store_3_27 <= data_store_1_9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_28 <= 0;
		end else begin
			if (andOp_468_out) begin
				data_store_3_28 <= in_out_data;
			end
			if (andOp_470_out) begin
				data_store_3_28 <= data_store_2_19;
			end
			if (andOp_474_out) begin
				data_store_3_28 <= data_store_1_10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_29 <= 0;
		end else begin
			if (andOp_477_out) begin
				data_store_3_29 <= phi_out_phi_7;
			end
			if (andOp_479_out) begin
				data_store_3_29 <= data_store_2_20;
			end
			if (andOp_483_out) begin
				data_store_3_29 <= data_store_4_38;
			end
			if (andOp_485_out) begin
				data_store_3_29 <= data_store_1_11;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_30 <= 0;
		end else begin
			if (andOp_488_out) begin
				data_store_3_30 <= rdata_ram_0;
			end
			if (andOp_490_out) begin
				data_store_3_30 <= data_store_2_21;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_31 <= 0;
		end else begin
			if (andOp_495_out) begin
				data_store_3_31 <= add_out_add_13;
			end
			if (andOp_497_out) begin
				data_store_3_31 <= data_store_2_22;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_32 <= 0;
		end else begin
			if (andOp_502_out) begin
				data_store_3_32 <= add_out_add_15;
			end
			if (andOp_504_out) begin
				data_store_3_32 <= data_store_2_23;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_33 <= 0;
		end else begin
			if (andOp_509_out) begin
				data_store_3_33 <= cmp_out_icmp_16;
			end
			if (andOp_511_out) begin
				data_store_3_33 <= data_store_2_24;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_34 <= 0;
		end else begin
			if (andOp_516_out) begin
				data_store_3_34 <= rdata_ram_0;
			end
			if (andOp_518_out) begin
				data_store_3_34 <= data_store_2_25;
			end
			if (andOp_522_out) begin
				data_store_3_34 <= data_store_4_43;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_35 <= 0;
		end else begin
			if (andOp_525_out) begin
				data_store_3_35 <= out_write_ready;
			end
			if (andOp_527_out) begin
				data_store_3_35 <= data_store_2_26;
			end
			if (andOp_531_out) begin
				data_store_3_35 <= data_store_4_44;
			end
			if (andOp_533_out) begin
				data_store_3_35 <= data_store_4_44;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_36 <= 0;
		end else begin
			if (andOp_536_out) begin
				data_store_4_36 <= in_read_ready;
			end
			if (andOp_538_out) begin
				data_store_4_36 <= data_store_3_27;
			end
			if (andOp_542_out) begin
				data_store_4_36 <= data_store_1_9;
			end
			if (andOp_544_out) begin
				data_store_4_36 <= data_store_1_9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_37 <= 0;
		end else begin
			if (andOp_547_out) begin
				data_store_4_37 <= in_out_data;
			end
			if (andOp_549_out) begin
				data_store_4_37 <= data_store_3_28;
			end
			if (andOp_553_out) begin
				data_store_4_37 <= data_store_1_10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_38 <= 0;
		end else begin
			if (andOp_556_out) begin
				data_store_4_38 <= phi_out_phi_7;
			end
			if (andOp_558_out) begin
				data_store_4_38 <= data_store_3_29;
			end
			if (andOp_562_out) begin
				data_store_4_38 <= data_store_4_38;
			end
			if (andOp_564_out) begin
				data_store_4_38 <= data_store_1_11;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_39 <= 0;
		end else begin
			if (andOp_567_out) begin
				data_store_4_39 <= rdata_ram_0;
			end
			if (andOp_569_out) begin
				data_store_4_39 <= data_store_3_30;
			end
			if (andOp_573_out) begin
				data_store_4_39 <= data_store_3_30;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_40 <= 0;
		end else begin
			if (andOp_576_out) begin
				data_store_4_40 <= add_out_add_13;
			end
			if (andOp_578_out) begin
				data_store_4_40 <= data_store_3_31;
			end
			if (andOp_582_out) begin
				data_store_4_40 <= data_store_3_31;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_41 <= 0;
		end else begin
			if (andOp_585_out) begin
				data_store_4_41 <= add_out_add_15;
			end
			if (andOp_587_out) begin
				data_store_4_41 <= data_store_3_32;
			end
			if (andOp_591_out) begin
				data_store_4_41 <= data_store_3_32;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_42 <= 0;
		end else begin
			if (andOp_594_out) begin
				data_store_4_42 <= cmp_out_icmp_16;
			end
			if (andOp_596_out) begin
				data_store_4_42 <= data_store_3_33;
			end
			if (andOp_600_out) begin
				data_store_4_42 <= data_store_3_33;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_43 <= 0;
		end else begin
			if (andOp_603_out) begin
				data_store_4_43 <= rdata_ram_0;
			end
			if (andOp_605_out) begin
				data_store_4_43 <= data_store_3_34;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_44 <= 0;
		end else begin
			if (andOp_610_out) begin
				data_store_4_44 <= out_write_ready;
			end
			if (andOp_612_out) begin
				data_store_4_44 <= data_store_3_35;
			end
			if (andOp_616_out) begin
				data_store_4_44 <= data_store_4_44;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_174_out) begin
				global_state <= 32'd1;
			end
			if (andOp_175_out) begin
				global_state <= 32'd3;
			end
			if (andOp_176_out) begin
				global_state <= 32'd4;
			end
			if (andOp_177_out) begin
				global_state <= 32'd4;
			end
			if (andOp_60_out) begin
				global_state <= 32'd2;
			end
			if (andOp_62_out) begin
				global_state <= 32'd1;
			end
			if (andOp_71_out) begin
				global_state <= 32'd1;
			end
			if (andOp_83_out) begin
				global_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			icmp_tmp_6 <= 0;
		end else begin
			if (andOp_197_out) begin
				icmp_tmp_6 <= cmp_out_icmp_16;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			phi_tmp_1 <= 0;
		end else begin
			if (andOp_194_out) begin
				phi_tmp_1 <= phi_out_phi_7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (1'd1) begin
				state_0_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_174_out) begin
				state_1_entry_BB_reg <= 32'd0;
			end
			if (andOp_62_out) begin
				state_1_entry_BB_reg <= 32'd9;
			end
			if (andOp_71_out) begin
				state_1_entry_BB_reg <= 32'd3;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_174_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_183_out) begin
				state_1_is_active <= 1'd0;
			end
			if (andOp_62_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_71_out) begin
				state_1_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_62_out) begin
				state_1_last_BB_reg <= 32'd9;
			end
			if (andOp_71_out) begin
				state_1_last_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_60_out) begin
				state_2_entry_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_185_out) begin
				state_2_is_active <= 1'd0;
			end
			if (andOp_60_out) begin
				state_2_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_60_out) begin
				state_2_last_BB_reg <= 32'd9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_175_out) begin
				state_3_entry_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_175_out) begin
				state_3_is_active <= 1'd1;
			end
			if (andOp_187_out) begin
				state_3_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_64_out) begin
				state_3_last_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_176_out) begin
				state_4_entry_BB_reg <= 32'd4;
			end
			if (andOp_177_out) begin
				state_4_entry_BB_reg <= 32'd2;
			end
			if (andOp_83_out) begin
				state_4_entry_BB_reg <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_176_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_177_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_193_out) begin
				state_4_is_active <= 1'd0;
			end
			if (andOp_83_out) begin
				state_4_is_active <= 1'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_83_out) begin
				state_4_last_BB_reg <= 32'd6;
			end
			if (andOp_85_out) begin
				state_4_last_BB_reg <= 32'd7;
			end
		end
	end

endmodule

