module channel_reduce_4(input [0:0] clk, input [0:0] rst, output [0:0] valid, output [31:0] in_in_data, output [0:0] in_read_valid, output [0:0] in_rst, output [0:0] in_write_valid, input [31:0] in_out_data, input [0:0] in_read_ready, input [0:0] in_write_ready, output [31:0] out_in_data, output [0:0] out_read_valid, output [0:0] out_rst, output [0:0] out_write_valid, input [31:0] out_out_data, input [0:0] out_read_ready, input [0:0] out_write_ready);

	reg [0:0] valid_reg;
	reg [31:0] in_in_data_reg;
	reg [0:0] in_read_valid_reg;
	reg [0:0] in_rst_reg;
	reg [0:0] in_write_valid_reg;
	reg [31:0] out_in_data_reg;
	reg [0:0] out_read_valid_reg;
	reg [0:0] out_rst_reg;
	reg [0:0] out_write_valid_reg;

	assign valid = valid_reg;
	assign in_in_data = in_in_data_reg;
	assign in_read_valid = in_read_valid_reg;
	assign in_rst = in_rst_reg;
	assign in_write_valid = in_write_valid_reg;
	assign out_in_data = out_in_data_reg;
	assign out_read_valid = out_read_valid_reg;
	assign out_rst = out_rst_reg;
	assign out_write_valid = out_write_valid_reg;

	// Start debug wires and ports

	initial begin
	end





	// End debug wires and ports

	// Start Functional Units
	br_dummy br_unit();

	reg [31:0] raddr_ram_0_reg;
	reg [31:0] waddr_ram_0_reg;
	reg [31:0] wdata_ram_0_reg;
	reg [0:0] wen_ram_0_reg;
	wire [31:0] rdata_ram_0;
	register #(.WIDTH(32)) ram_0(.clk(clk), .raddr(raddr_ram_0_reg), .rdata(rdata_ram_0), .rst(rst), .waddr(waddr_ram_0_reg), .wdata(wdata_ram_0_reg), .wen(wen_ram_0_reg));

	reg [31:0] add_in0_add_12;
	reg [31:0] add_in1_add_12;
	wire [31:0] add_out_add_12;
	add #(.WIDTH(32)) add_add_12(.in0(add_in0_add_12), .in1(add_in1_add_12), .out(add_out_add_12));

	reg [31:0] add_in0_add_14;
	reg [31:0] add_in1_add_14;
	wire [31:0] add_out_add_14;
	add #(.WIDTH(32)) add_add_14(.in0(add_in0_add_14), .in1(add_in1_add_14), .out(add_out_add_14));

	reg [31:0] cmp_in0_icmp_15;
	reg [31:0] cmp_in1_icmp_15;
	wire [0:0] cmp_out_icmp_15;
	eq #(.WIDTH(32)) icmp_15(.in0(cmp_in0_icmp_15), .in1(cmp_in1_icmp_15), .out(cmp_out_icmp_15));

	add call_20();

	reg [63:0] phi_in_phi_6;
	reg [31:0] phi_last_block_phi_6;
	reg [63:0] phi_s_phi_6;
	wire [31:0] phi_out_phi_6;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_6(.in(phi_in_phi_6), .last_block(phi_last_block_phi_6), .out(phi_out_phi_6), .s(phi_s_phi_6));

	add alloca_1();

	add bitcast_2();

	add call_3();

	reg [0:0] bb_0_active_in_data;
	wire [0:0] bb_0_active_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active(.in_data(bb_0_active_in_data), .out_data(bb_0_active_out_data));

	reg [31:0] eq_0_in0;
	reg [31:0] eq_0_in1;
	wire [0:0] eq_0_out;
	eq #(.WIDTH(32)) eq_0(.in0(eq_0_in0), .in1(eq_0_in1), .out(eq_0_out));

	reg [0:0] andOp_1_in0;
	reg [0:0] andOp_1_in1;
	wire [0:0] andOp_1_out;
	andOp #(.WIDTH(1)) andOp_1(.in0(andOp_1_in0), .in1(andOp_1_in1), .out(andOp_1_out));

	reg [0:0] andOp_2_in0;
	reg [0:0] andOp_2_in1;
	wire [0:0] andOp_2_out;
	andOp #(.WIDTH(1)) andOp_2(.in0(andOp_2_in0), .in1(andOp_2_in1), .out(andOp_2_out));

	reg [0:0] br_0_happened_in_data;
	wire [0:0] br_0_happened_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened(.in_data(br_0_happened_in_data), .out_data(br_0_happened_out_data));

	reg [0:0] notOp_3_in0;
	wire [0:0] notOp_3_out;
	notOp #(.WIDTH(1)) notOp_3(.in(notOp_3_in0), .out(notOp_3_out));

	reg [0:0] bb_1_active_in_data;
	wire [0:0] bb_1_active_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active(.in_data(bb_1_active_in_data), .out_data(bb_1_active_out_data));

	reg [31:0] eq_4_in0;
	reg [31:0] eq_4_in1;
	wire [0:0] eq_4_out;
	eq #(.WIDTH(32)) eq_4(.in0(eq_4_in0), .in1(eq_4_in1), .out(eq_4_out));

	reg [0:0] andOp_5_in0;
	reg [0:0] andOp_5_in1;
	wire [0:0] andOp_5_out;
	andOp #(.WIDTH(1)) andOp_5(.in0(andOp_5_in0), .in1(andOp_5_in1), .out(andOp_5_out));

	reg [0:0] andOp_6_in0;
	reg [0:0] andOp_6_in1;
	wire [0:0] andOp_6_out;
	andOp #(.WIDTH(1)) andOp_6(.in0(andOp_6_in0), .in1(andOp_6_in1), .out(andOp_6_out));

	reg [0:0] br_1_happened_in_data;
	wire [0:0] br_1_happened_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened(.in_data(br_1_happened_in_data), .out_data(br_1_happened_out_data));

	reg [0:0] notOp_7_in0;
	wire [0:0] notOp_7_out;
	notOp #(.WIDTH(1)) notOp_7(.in(notOp_7_in0), .out(notOp_7_out));

	reg [0:0] bb_2_active_in_data;
	wire [0:0] bb_2_active_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active(.in_data(bb_2_active_in_data), .out_data(bb_2_active_out_data));

	reg [0:0] bb_3_active_in_data;
	wire [0:0] bb_3_active_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active(.in_data(bb_3_active_in_data), .out_data(bb_3_active_out_data));

	reg [31:0] eq_8_in0;
	reg [31:0] eq_8_in1;
	wire [0:0] eq_8_out;
	eq #(.WIDTH(32)) eq_8(.in0(eq_8_in0), .in1(eq_8_in1), .out(eq_8_out));

	reg [0:0] andOp_9_in0;
	reg [0:0] andOp_9_in1;
	wire [0:0] andOp_9_out;
	andOp #(.WIDTH(1)) andOp_9(.in0(andOp_9_in0), .in1(andOp_9_in1), .out(andOp_9_out));

	reg [0:0] andOp_10_in0;
	reg [0:0] andOp_10_in1;
	wire [0:0] andOp_10_out;
	andOp #(.WIDTH(1)) andOp_10(.in0(andOp_10_in0), .in1(andOp_10_in1), .out(andOp_10_out));

	reg [0:0] br_3_happened_in_data;
	wire [0:0] br_3_happened_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened(.in_data(br_3_happened_in_data), .out_data(br_3_happened_out_data));

	reg [0:0] notOp_11_in0;
	wire [0:0] notOp_11_out;
	notOp #(.WIDTH(1)) notOp_11(.in(notOp_11_in0), .out(notOp_11_out));

	reg [0:0] bb_4_active_in_data;
	wire [0:0] bb_4_active_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active(.in_data(bb_4_active_in_data), .out_data(bb_4_active_out_data));

	reg [31:0] eq_12_in0;
	reg [31:0] eq_12_in1;
	wire [0:0] eq_12_out;
	eq #(.WIDTH(32)) eq_12(.in0(eq_12_in0), .in1(eq_12_in1), .out(eq_12_out));

	reg [0:0] andOp_13_in0;
	reg [0:0] andOp_13_in1;
	wire [0:0] andOp_13_out;
	andOp #(.WIDTH(1)) andOp_13(.in0(andOp_13_in0), .in1(andOp_13_in1), .out(andOp_13_out));

	reg [0:0] andOp_14_in0;
	reg [0:0] andOp_14_in1;
	wire [0:0] andOp_14_out;
	andOp #(.WIDTH(1)) andOp_14(.in0(andOp_14_in0), .in1(andOp_14_in1), .out(andOp_14_out));

	reg [0:0] br_4_happened_in_data;
	wire [0:0] br_4_happened_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened(.in_data(br_4_happened_in_data), .out_data(br_4_happened_out_data));

	reg [0:0] notOp_15_in0;
	wire [0:0] notOp_15_out;
	notOp #(.WIDTH(1)) notOp_15(.in(notOp_15_in0), .out(notOp_15_out));

	reg [0:0] andOp_16_in0;
	reg [0:0] andOp_16_in1;
	wire [0:0] andOp_16_out;
	andOp #(.WIDTH(1)) andOp_16(.in0(andOp_16_in0), .in1(andOp_16_in1), .out(andOp_16_out));

	reg [0:0] notOp_17_in0;
	wire [0:0] notOp_17_out;
	notOp #(.WIDTH(1)) notOp_17(.in(notOp_17_in0), .out(notOp_17_out));

	reg [0:0] andOp_18_in0;
	reg [0:0] andOp_18_in1;
	wire [0:0] andOp_18_out;
	andOp #(.WIDTH(1)) andOp_18(.in0(andOp_18_in0), .in1(andOp_18_in1), .out(andOp_18_out));

	reg [0:0] bb_5_active_in_data;
	wire [0:0] bb_5_active_out_data;
	hls_wire #(.WIDTH(1)) bb_5_active(.in_data(bb_5_active_in_data), .out_data(bb_5_active_out_data));

	reg [31:0] eq_19_in0;
	reg [31:0] eq_19_in1;
	wire [0:0] eq_19_out;
	eq #(.WIDTH(32)) eq_19(.in0(eq_19_in0), .in1(eq_19_in1), .out(eq_19_out));

	reg [0:0] andOp_20_in0;
	reg [0:0] andOp_20_in1;
	wire [0:0] andOp_20_out;
	andOp #(.WIDTH(1)) andOp_20(.in0(andOp_20_in0), .in1(andOp_20_in1), .out(andOp_20_out));

	reg [0:0] andOp_21_in0;
	reg [0:0] andOp_21_in1;
	wire [0:0] andOp_21_out;
	andOp #(.WIDTH(1)) andOp_21(.in0(andOp_21_in0), .in1(andOp_21_in1), .out(andOp_21_out));

	reg [0:0] br_5_happened_in_data;
	wire [0:0] br_5_happened_out_data;
	hls_wire #(.WIDTH(1)) br_5_happened(.in_data(br_5_happened_in_data), .out_data(br_5_happened_out_data));

	reg [0:0] notOp_22_in0;
	wire [0:0] notOp_22_out;
	notOp #(.WIDTH(1)) notOp_22(.in(notOp_22_in0), .out(notOp_22_out));

	reg [0:0] bb_6_active_in_data;
	wire [0:0] bb_6_active_out_data;
	hls_wire #(.WIDTH(1)) bb_6_active(.in_data(bb_6_active_in_data), .out_data(bb_6_active_out_data));

	reg [31:0] eq_23_in0;
	reg [31:0] eq_23_in1;
	wire [0:0] eq_23_out;
	eq #(.WIDTH(32)) eq_23(.in0(eq_23_in0), .in1(eq_23_in1), .out(eq_23_out));

	reg [0:0] andOp_24_in0;
	reg [0:0] andOp_24_in1;
	wire [0:0] andOp_24_out;
	andOp #(.WIDTH(1)) andOp_24(.in0(andOp_24_in0), .in1(andOp_24_in1), .out(andOp_24_out));

	reg [0:0] andOp_25_in0;
	reg [0:0] andOp_25_in1;
	wire [0:0] andOp_25_out;
	andOp #(.WIDTH(1)) andOp_25(.in0(andOp_25_in0), .in1(andOp_25_in1), .out(andOp_25_out));

	reg [0:0] br_6_happened_in_data;
	wire [0:0] br_6_happened_out_data;
	hls_wire #(.WIDTH(1)) br_6_happened(.in_data(br_6_happened_in_data), .out_data(br_6_happened_out_data));

	reg [0:0] notOp_26_in0;
	wire [0:0] notOp_26_out;
	notOp #(.WIDTH(1)) notOp_26(.in(notOp_26_in0), .out(notOp_26_out));

	reg [0:0] andOp_27_in0;
	reg [0:0] andOp_27_in1;
	wire [0:0] andOp_27_out;
	andOp #(.WIDTH(1)) andOp_27(.in0(andOp_27_in0), .in1(andOp_27_in1), .out(andOp_27_out));

	reg [0:0] notOp_28_in0;
	wire [0:0] notOp_28_out;
	notOp #(.WIDTH(1)) notOp_28(.in(notOp_28_in0), .out(notOp_28_out));

	reg [0:0] andOp_29_in0;
	reg [0:0] andOp_29_in1;
	wire [0:0] andOp_29_out;
	andOp #(.WIDTH(1)) andOp_29(.in0(andOp_29_in0), .in1(andOp_29_in1), .out(andOp_29_out));

	reg [0:0] bb_7_active_in_data;
	wire [0:0] bb_7_active_out_data;
	hls_wire #(.WIDTH(1)) bb_7_active(.in_data(bb_7_active_in_data), .out_data(bb_7_active_out_data));

	reg [31:0] eq_30_in0;
	reg [31:0] eq_30_in1;
	wire [0:0] eq_30_out;
	eq #(.WIDTH(32)) eq_30(.in0(eq_30_in0), .in1(eq_30_in1), .out(eq_30_out));

	reg [0:0] andOp_31_in0;
	reg [0:0] andOp_31_in1;
	wire [0:0] andOp_31_out;
	andOp #(.WIDTH(1)) andOp_31(.in0(andOp_31_in0), .in1(andOp_31_in1), .out(andOp_31_out));

	reg [0:0] andOp_32_in0;
	reg [0:0] andOp_32_in1;
	wire [0:0] andOp_32_out;
	andOp #(.WIDTH(1)) andOp_32(.in0(andOp_32_in0), .in1(andOp_32_in1), .out(andOp_32_out));

	reg [0:0] br_7_happened_in_data;
	wire [0:0] br_7_happened_out_data;
	hls_wire #(.WIDTH(1)) br_7_happened(.in_data(br_7_happened_in_data), .out_data(br_7_happened_out_data));

	reg [0:0] notOp_33_in0;
	wire [0:0] notOp_33_out;
	notOp #(.WIDTH(1)) notOp_33(.in(notOp_33_in0), .out(notOp_33_out));

	reg [0:0] bb_8_active_in_data;
	wire [0:0] bb_8_active_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active(.in_data(bb_8_active_in_data), .out_data(bb_8_active_out_data));

	reg [31:0] eq_34_in0;
	reg [31:0] eq_34_in1;
	wire [0:0] eq_34_out;
	eq #(.WIDTH(32)) eq_34(.in0(eq_34_in0), .in1(eq_34_in1), .out(eq_34_out));

	reg [0:0] andOp_35_in0;
	reg [0:0] andOp_35_in1;
	wire [0:0] andOp_35_out;
	andOp #(.WIDTH(1)) andOp_35(.in0(andOp_35_in0), .in1(andOp_35_in1), .out(andOp_35_out));

	reg [0:0] andOp_36_in0;
	reg [0:0] andOp_36_in1;
	wire [0:0] andOp_36_out;
	andOp #(.WIDTH(1)) andOp_36(.in0(andOp_36_in0), .in1(andOp_36_in1), .out(andOp_36_out));

	reg [0:0] br_8_happened_in_data;
	wire [0:0] br_8_happened_out_data;
	hls_wire #(.WIDTH(1)) br_8_happened(.in_data(br_8_happened_in_data), .out_data(br_8_happened_out_data));

	reg [0:0] notOp_37_in0;
	wire [0:0] notOp_37_out;
	notOp #(.WIDTH(1)) notOp_37(.in(notOp_37_in0), .out(notOp_37_out));

	reg [0:0] bb_9_active_in_data;
	wire [0:0] bb_9_active_out_data;
	hls_wire #(.WIDTH(1)) bb_9_active(.in_data(bb_9_active_in_data), .out_data(bb_9_active_out_data));

	reg [31:0] eq_38_in0;
	reg [31:0] eq_38_in1;
	wire [0:0] eq_38_out;
	eq #(.WIDTH(32)) eq_38(.in0(eq_38_in0), .in1(eq_38_in1), .out(eq_38_out));

	reg [0:0] andOp_39_in0;
	reg [0:0] andOp_39_in1;
	wire [0:0] andOp_39_out;
	andOp #(.WIDTH(1)) andOp_39(.in0(andOp_39_in0), .in1(andOp_39_in1), .out(andOp_39_out));

	reg [0:0] andOp_40_in0;
	reg [0:0] andOp_40_in1;
	wire [0:0] andOp_40_out;
	andOp #(.WIDTH(1)) andOp_40(.in0(andOp_40_in0), .in1(andOp_40_in1), .out(andOp_40_out));

	reg [0:0] br_9_happened_in_data;
	wire [0:0] br_9_happened_out_data;
	hls_wire #(.WIDTH(1)) br_9_happened(.in_data(br_9_happened_in_data), .out_data(br_9_happened_out_data));

	reg [0:0] notOp_41_in0;
	wire [0:0] notOp_41_out;
	notOp #(.WIDTH(1)) notOp_41(.in(notOp_41_in0), .out(notOp_41_out));

	reg [0:0] andOp_42_in0;
	reg [0:0] andOp_42_in1;
	wire [0:0] andOp_42_out;
	andOp #(.WIDTH(1)) andOp_42(.in0(andOp_42_in0), .in1(andOp_42_in1), .out(andOp_42_out));

	reg [0:0] notOp_43_in0;
	wire [0:0] notOp_43_out;
	notOp #(.WIDTH(1)) notOp_43(.in(notOp_43_in0), .out(notOp_43_out));

	reg [0:0] andOp_44_in0;
	reg [0:0] andOp_44_in1;
	wire [0:0] andOp_44_out;
	andOp #(.WIDTH(1)) andOp_44(.in0(andOp_44_in0), .in1(andOp_44_in1), .out(andOp_44_out));

	reg [0:0] bb_10_active_in_data;
	wire [0:0] bb_10_active_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active(.in_data(bb_10_active_in_data), .out_data(bb_10_active_out_data));

	reg [31:0] eq_45_in0;
	reg [31:0] eq_45_in1;
	wire [0:0] eq_45_out;
	eq #(.WIDTH(32)) eq_45(.in0(eq_45_in0), .in1(eq_45_in1), .out(eq_45_out));

	reg [0:0] andOp_46_in0;
	reg [0:0] andOp_46_in1;
	wire [0:0] andOp_46_out;
	andOp #(.WIDTH(1)) andOp_46(.in0(andOp_46_in0), .in1(andOp_46_in1), .out(andOp_46_out));

	reg [0:0] andOp_47_in0;
	reg [0:0] andOp_47_in1;
	wire [0:0] andOp_47_out;
	andOp #(.WIDTH(1)) andOp_47(.in0(andOp_47_in0), .in1(andOp_47_in1), .out(andOp_47_out));

	reg [0:0] br_10_happened_in_data;
	wire [0:0] br_10_happened_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened(.in_data(br_10_happened_in_data), .out_data(br_10_happened_out_data));

	reg [0:0] notOp_48_in0;
	wire [0:0] notOp_48_out;
	notOp #(.WIDTH(1)) notOp_48(.in(notOp_48_in0), .out(notOp_48_out));

	reg [31:0] eq_49_in0;
	reg [31:0] eq_49_in1;
	wire [0:0] eq_49_out;
	eq #(.WIDTH(32)) eq_49(.in0(eq_49_in0), .in1(eq_49_in1), .out(eq_49_out));

	reg [31:0] eq_50_in0;
	reg [31:0] eq_50_in1;
	wire [0:0] eq_50_out;
	eq #(.WIDTH(32)) eq_50(.in0(eq_50_in0), .in1(eq_50_in1), .out(eq_50_out));

	reg [0:0] orOp_51_in0;
	reg [0:0] orOp_51_in1;
	wire [0:0] orOp_51_out;
	orOp #(.WIDTH(1)) orOp_51(.in0(orOp_51_in0), .in1(orOp_51_in1), .out(orOp_51_out));

	reg [31:0] eq_52_in0;
	reg [31:0] eq_52_in1;
	wire [0:0] eq_52_out;
	eq #(.WIDTH(32)) eq_52(.in0(eq_52_in0), .in1(eq_52_in1), .out(eq_52_out));

	reg [0:0] orOp_53_in0;
	reg [0:0] orOp_53_in1;
	wire [0:0] orOp_53_out;
	orOp #(.WIDTH(1)) orOp_53(.in0(orOp_53_in0), .in1(orOp_53_in1), .out(orOp_53_out));

	reg [31:0] eq_54_in0;
	reg [31:0] eq_54_in1;
	wire [0:0] eq_54_out;
	eq #(.WIDTH(32)) eq_54(.in0(eq_54_in0), .in1(eq_54_in1), .out(eq_54_out));

	reg [0:0] orOp_55_in0;
	reg [0:0] orOp_55_in1;
	wire [0:0] orOp_55_out;
	orOp #(.WIDTH(1)) orOp_55(.in0(orOp_55_in0), .in1(orOp_55_in1), .out(orOp_55_out));

	reg [31:0] eq_56_in0;
	reg [31:0] eq_56_in1;
	wire [0:0] eq_56_out;
	eq #(.WIDTH(32)) eq_56(.in0(eq_56_in0), .in1(eq_56_in1), .out(eq_56_out));

	reg [0:0] orOp_57_in0;
	reg [0:0] orOp_57_in1;
	wire [0:0] orOp_57_out;
	orOp #(.WIDTH(1)) orOp_57(.in0(orOp_57_in0), .in1(orOp_57_in1), .out(orOp_57_out));

	reg [31:0] eq_58_in0;
	reg [31:0] eq_58_in1;
	wire [0:0] eq_58_out;
	eq #(.WIDTH(32)) eq_58(.in0(eq_58_in0), .in1(eq_58_in1), .out(eq_58_out));

	reg [0:0] orOp_59_in0;
	reg [0:0] orOp_59_in1;
	wire [0:0] orOp_59_out;
	orOp #(.WIDTH(1)) orOp_59(.in0(orOp_59_in0), .in1(orOp_59_in1), .out(orOp_59_out));

	reg [31:0] eq_60_in0;
	reg [31:0] eq_60_in1;
	wire [0:0] eq_60_out;
	eq #(.WIDTH(32)) eq_60(.in0(eq_60_in0), .in1(eq_60_in1), .out(eq_60_out));

	reg [0:0] orOp_61_in0;
	reg [0:0] orOp_61_in1;
	wire [0:0] orOp_61_out;
	orOp #(.WIDTH(1)) orOp_61(.in0(orOp_61_in0), .in1(orOp_61_in1), .out(orOp_61_out));

	reg [31:0] eq_62_in0;
	reg [31:0] eq_62_in1;
	wire [0:0] eq_62_out;
	eq #(.WIDTH(32)) eq_62(.in0(eq_62_in0), .in1(eq_62_in1), .out(eq_62_out));

	reg [0:0] orOp_63_in0;
	reg [0:0] orOp_63_in1;
	wire [0:0] orOp_63_out;
	orOp #(.WIDTH(1)) orOp_63(.in0(orOp_63_in0), .in1(orOp_63_in1), .out(orOp_63_out));

	reg [31:0] eq_64_in0;
	reg [31:0] eq_64_in1;
	wire [0:0] eq_64_out;
	eq #(.WIDTH(32)) eq_64(.in0(eq_64_in0), .in1(eq_64_in1), .out(eq_64_out));

	reg [0:0] orOp_65_in0;
	reg [0:0] orOp_65_in1;
	wire [0:0] orOp_65_out;
	orOp #(.WIDTH(1)) orOp_65(.in0(orOp_65_in0), .in1(orOp_65_in1), .out(orOp_65_out));

	reg [31:0] eq_66_in0;
	reg [31:0] eq_66_in1;
	wire [0:0] eq_66_out;
	eq #(.WIDTH(32)) eq_66(.in0(eq_66_in0), .in1(eq_66_in1), .out(eq_66_out));

	reg [0:0] orOp_67_in0;
	reg [0:0] orOp_67_in1;
	wire [0:0] orOp_67_out;
	orOp #(.WIDTH(1)) orOp_67(.in0(orOp_67_in0), .in1(orOp_67_in1), .out(orOp_67_out));

	reg [31:0] eq_68_in0;
	reg [31:0] eq_68_in1;
	wire [0:0] eq_68_out;
	eq #(.WIDTH(32)) eq_68(.in0(eq_68_in0), .in1(eq_68_in1), .out(eq_68_out));

	reg [0:0] orOp_69_in0;
	reg [0:0] orOp_69_in1;
	wire [0:0] orOp_69_out;
	orOp #(.WIDTH(1)) orOp_69(.in0(orOp_69_in0), .in1(orOp_69_in1), .out(orOp_69_out));

	reg [31:0] eq_70_in0;
	reg [31:0] eq_70_in1;
	wire [0:0] eq_70_out;
	eq #(.WIDTH(32)) eq_70(.in0(eq_70_in0), .in1(eq_70_in1), .out(eq_70_out));

	reg [0:0] andOp_71_in0;
	reg [0:0] andOp_71_in1;
	wire [0:0] andOp_71_out;
	andOp #(.WIDTH(1)) andOp_71(.in0(andOp_71_in0), .in1(andOp_71_in1), .out(andOp_71_out));

	reg [31:0] eq_72_in0;
	reg [31:0] eq_72_in1;
	wire [0:0] eq_72_out;
	eq #(.WIDTH(32)) eq_72(.in0(eq_72_in0), .in1(eq_72_in1), .out(eq_72_out));

	reg [0:0] andOp_73_in0;
	reg [0:0] andOp_73_in1;
	wire [0:0] andOp_73_out;
	andOp #(.WIDTH(1)) andOp_73(.in0(andOp_73_in0), .in1(andOp_73_in1), .out(andOp_73_out));

	reg [31:0] eq_74_in0;
	reg [31:0] eq_74_in1;
	wire [0:0] eq_74_out;
	eq #(.WIDTH(32)) eq_74(.in0(eq_74_in0), .in1(eq_74_in1), .out(eq_74_out));

	reg [0:0] andOp_75_in0;
	reg [0:0] andOp_75_in1;
	wire [0:0] andOp_75_out;
	andOp #(.WIDTH(1)) andOp_75(.in0(andOp_75_in0), .in1(andOp_75_in1), .out(andOp_75_out));

	reg [31:0] eq_76_in0;
	reg [31:0] eq_76_in1;
	wire [0:0] eq_76_out;
	eq #(.WIDTH(32)) eq_76(.in0(eq_76_in0), .in1(eq_76_in1), .out(eq_76_out));

	reg [0:0] andOp_77_in0;
	reg [0:0] andOp_77_in1;
	wire [0:0] andOp_77_out;
	andOp #(.WIDTH(1)) andOp_77(.in0(andOp_77_in0), .in1(andOp_77_in1), .out(andOp_77_out));

	reg [31:0] eq_78_in0;
	reg [31:0] eq_78_in1;
	wire [0:0] eq_78_out;
	eq #(.WIDTH(32)) eq_78(.in0(eq_78_in0), .in1(eq_78_in1), .out(eq_78_out));

	reg [0:0] andOp_79_in0;
	reg [0:0] andOp_79_in1;
	wire [0:0] andOp_79_out;
	andOp #(.WIDTH(1)) andOp_79(.in0(andOp_79_in0), .in1(andOp_79_in1), .out(andOp_79_out));

	reg [31:0] bb_0_predecessor_in_data;
	wire [31:0] bb_0_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor(.in_data(bb_0_predecessor_in_data), .out_data(bb_0_predecessor_out_data));

	reg [31:0] eq_80_in0;
	reg [31:0] eq_80_in1;
	wire [0:0] eq_80_out;
	eq #(.WIDTH(32)) eq_80(.in0(eq_80_in0), .in1(eq_80_in1), .out(eq_80_out));

	reg [31:0] bb_1_predecessor_in_data;
	wire [31:0] bb_1_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor(.in_data(bb_1_predecessor_in_data), .out_data(bb_1_predecessor_out_data));

	reg [31:0] eq_81_in0;
	reg [31:0] eq_81_in1;
	wire [0:0] eq_81_out;
	eq #(.WIDTH(32)) eq_81(.in0(eq_81_in0), .in1(eq_81_in1), .out(eq_81_out));

	reg [0:0] notOp_82_in0;
	wire [0:0] notOp_82_out;
	notOp #(.WIDTH(1)) notOp_82(.in(notOp_82_in0), .out(notOp_82_out));

	reg [0:0] andOp_83_in0;
	reg [0:0] andOp_83_in1;
	wire [0:0] andOp_83_out;
	andOp #(.WIDTH(1)) andOp_83(.in0(andOp_83_in0), .in1(andOp_83_in1), .out(andOp_83_out));

	reg [31:0] bb_2_predecessor_in_data;
	wire [31:0] bb_2_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor(.in_data(bb_2_predecessor_in_data), .out_data(bb_2_predecessor_out_data));

	reg [31:0] eq_84_in0;
	reg [31:0] eq_84_in1;
	wire [0:0] eq_84_out;
	eq #(.WIDTH(32)) eq_84(.in0(eq_84_in0), .in1(eq_84_in1), .out(eq_84_out));

	reg [0:0] notOp_85_in0;
	wire [0:0] notOp_85_out;
	notOp #(.WIDTH(1)) notOp_85(.in(notOp_85_in0), .out(notOp_85_out));

	reg [0:0] andOp_86_in0;
	reg [0:0] andOp_86_in1;
	wire [0:0] andOp_86_out;
	andOp #(.WIDTH(1)) andOp_86(.in0(andOp_86_in0), .in1(andOp_86_in1), .out(andOp_86_out));

	reg [31:0] bb_3_predecessor_in_data;
	wire [31:0] bb_3_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor(.in_data(bb_3_predecessor_in_data), .out_data(bb_3_predecessor_out_data));

	reg [31:0] eq_87_in0;
	reg [31:0] eq_87_in1;
	wire [0:0] eq_87_out;
	eq #(.WIDTH(32)) eq_87(.in0(eq_87_in0), .in1(eq_87_in1), .out(eq_87_out));

	reg [0:0] notOp_88_in0;
	wire [0:0] notOp_88_out;
	notOp #(.WIDTH(1)) notOp_88(.in(notOp_88_in0), .out(notOp_88_out));

	reg [0:0] andOp_89_in0;
	reg [0:0] andOp_89_in1;
	wire [0:0] andOp_89_out;
	andOp #(.WIDTH(1)) andOp_89(.in0(andOp_89_in0), .in1(andOp_89_in1), .out(andOp_89_out));

	reg [31:0] bb_4_predecessor_in_data;
	wire [31:0] bb_4_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor(.in_data(bb_4_predecessor_in_data), .out_data(bb_4_predecessor_out_data));

	reg [31:0] eq_90_in0;
	reg [31:0] eq_90_in1;
	wire [0:0] eq_90_out;
	eq #(.WIDTH(32)) eq_90(.in0(eq_90_in0), .in1(eq_90_in1), .out(eq_90_out));

	reg [0:0] notOp_91_in0;
	wire [0:0] notOp_91_out;
	notOp #(.WIDTH(1)) notOp_91(.in(notOp_91_in0), .out(notOp_91_out));

	reg [0:0] andOp_92_in0;
	reg [0:0] andOp_92_in1;
	wire [0:0] andOp_92_out;
	andOp #(.WIDTH(1)) andOp_92(.in0(andOp_92_in0), .in1(andOp_92_in1), .out(andOp_92_out));

	reg [31:0] bb_5_predecessor_in_data;
	wire [31:0] bb_5_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_5_predecessor(.in_data(bb_5_predecessor_in_data), .out_data(bb_5_predecessor_out_data));

	reg [31:0] eq_93_in0;
	reg [31:0] eq_93_in1;
	wire [0:0] eq_93_out;
	eq #(.WIDTH(32)) eq_93(.in0(eq_93_in0), .in1(eq_93_in1), .out(eq_93_out));

	reg [0:0] notOp_94_in0;
	wire [0:0] notOp_94_out;
	notOp #(.WIDTH(1)) notOp_94(.in(notOp_94_in0), .out(notOp_94_out));

	reg [0:0] andOp_95_in0;
	reg [0:0] andOp_95_in1;
	wire [0:0] andOp_95_out;
	andOp #(.WIDTH(1)) andOp_95(.in0(andOp_95_in0), .in1(andOp_95_in1), .out(andOp_95_out));

	reg [31:0] bb_6_predecessor_in_data;
	wire [31:0] bb_6_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_6_predecessor(.in_data(bb_6_predecessor_in_data), .out_data(bb_6_predecessor_out_data));

	reg [31:0] eq_96_in0;
	reg [31:0] eq_96_in1;
	wire [0:0] eq_96_out;
	eq #(.WIDTH(32)) eq_96(.in0(eq_96_in0), .in1(eq_96_in1), .out(eq_96_out));

	reg [0:0] notOp_97_in0;
	wire [0:0] notOp_97_out;
	notOp #(.WIDTH(1)) notOp_97(.in(notOp_97_in0), .out(notOp_97_out));

	reg [0:0] andOp_98_in0;
	reg [0:0] andOp_98_in1;
	wire [0:0] andOp_98_out;
	andOp #(.WIDTH(1)) andOp_98(.in0(andOp_98_in0), .in1(andOp_98_in1), .out(andOp_98_out));

	reg [31:0] bb_7_predecessor_in_data;
	wire [31:0] bb_7_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_7_predecessor(.in_data(bb_7_predecessor_in_data), .out_data(bb_7_predecessor_out_data));

	reg [31:0] eq_99_in0;
	reg [31:0] eq_99_in1;
	wire [0:0] eq_99_out;
	eq #(.WIDTH(32)) eq_99(.in0(eq_99_in0), .in1(eq_99_in1), .out(eq_99_out));

	reg [0:0] notOp_100_in0;
	wire [0:0] notOp_100_out;
	notOp #(.WIDTH(1)) notOp_100(.in(notOp_100_in0), .out(notOp_100_out));

	reg [0:0] andOp_101_in0;
	reg [0:0] andOp_101_in1;
	wire [0:0] andOp_101_out;
	andOp #(.WIDTH(1)) andOp_101(.in0(andOp_101_in0), .in1(andOp_101_in1), .out(andOp_101_out));

	reg [31:0] bb_8_predecessor_in_data;
	wire [31:0] bb_8_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor(.in_data(bb_8_predecessor_in_data), .out_data(bb_8_predecessor_out_data));

	reg [31:0] eq_102_in0;
	reg [31:0] eq_102_in1;
	wire [0:0] eq_102_out;
	eq #(.WIDTH(32)) eq_102(.in0(eq_102_in0), .in1(eq_102_in1), .out(eq_102_out));

	reg [0:0] notOp_103_in0;
	wire [0:0] notOp_103_out;
	notOp #(.WIDTH(1)) notOp_103(.in(notOp_103_in0), .out(notOp_103_out));

	reg [0:0] andOp_104_in0;
	reg [0:0] andOp_104_in1;
	wire [0:0] andOp_104_out;
	andOp #(.WIDTH(1)) andOp_104(.in0(andOp_104_in0), .in1(andOp_104_in1), .out(andOp_104_out));

	reg [31:0] bb_9_predecessor_in_data;
	wire [31:0] bb_9_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_9_predecessor(.in_data(bb_9_predecessor_in_data), .out_data(bb_9_predecessor_out_data));

	reg [31:0] eq_105_in0;
	reg [31:0] eq_105_in1;
	wire [0:0] eq_105_out;
	eq #(.WIDTH(32)) eq_105(.in0(eq_105_in0), .in1(eq_105_in1), .out(eq_105_out));

	reg [0:0] notOp_106_in0;
	wire [0:0] notOp_106_out;
	notOp #(.WIDTH(1)) notOp_106(.in(notOp_106_in0), .out(notOp_106_out));

	reg [0:0] andOp_107_in0;
	reg [0:0] andOp_107_in1;
	wire [0:0] andOp_107_out;
	andOp #(.WIDTH(1)) andOp_107(.in0(andOp_107_in0), .in1(andOp_107_in1), .out(andOp_107_out));

	reg [31:0] bb_10_predecessor_in_data;
	wire [31:0] bb_10_predecessor_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor(.in_data(bb_10_predecessor_in_data), .out_data(bb_10_predecessor_out_data));

	reg [31:0] eq_108_in0;
	reg [31:0] eq_108_in1;
	wire [0:0] eq_108_out;
	eq #(.WIDTH(32)) eq_108(.in0(eq_108_in0), .in1(eq_108_in1), .out(eq_108_out));

	reg [0:0] notOp_109_in0;
	wire [0:0] notOp_109_out;
	notOp #(.WIDTH(1)) notOp_109(.in(notOp_109_in0), .out(notOp_109_out));

	reg [0:0] andOp_110_in0;
	reg [0:0] andOp_110_in1;
	wire [0:0] andOp_110_out;
	andOp #(.WIDTH(1)) andOp_110(.in0(andOp_110_in0), .in1(andOp_110_in1), .out(andOp_110_out));

	reg [31:0] eq_111_in0;
	reg [31:0] eq_111_in1;
	wire [0:0] eq_111_out;
	eq #(.WIDTH(32)) eq_111(.in0(eq_111_in0), .in1(eq_111_in1), .out(eq_111_out));

	reg [0:0] andOp_112_in0;
	reg [0:0] andOp_112_in1;
	wire [0:0] andOp_112_out;
	andOp #(.WIDTH(1)) andOp_112(.in0(andOp_112_in0), .in1(andOp_112_in1), .out(andOp_112_out));

	reg [31:0] eq_113_in0;
	reg [31:0] eq_113_in1;
	wire [0:0] eq_113_out;
	eq #(.WIDTH(32)) eq_113(.in0(eq_113_in0), .in1(eq_113_in1), .out(eq_113_out));

	reg [0:0] andOp_114_in0;
	reg [0:0] andOp_114_in1;
	wire [0:0] andOp_114_out;
	andOp #(.WIDTH(1)) andOp_114(.in0(andOp_114_in0), .in1(andOp_114_in1), .out(andOp_114_out));

	reg [31:0] eq_115_in0;
	reg [31:0] eq_115_in1;
	wire [0:0] eq_115_out;
	eq #(.WIDTH(32)) eq_115(.in0(eq_115_in0), .in1(eq_115_in1), .out(eq_115_out));

	reg [0:0] andOp_116_in0;
	reg [0:0] andOp_116_in1;
	wire [0:0] andOp_116_out;
	andOp #(.WIDTH(1)) andOp_116(.in0(andOp_116_in0), .in1(andOp_116_in1), .out(andOp_116_out));

	reg [31:0] eq_117_in0;
	reg [31:0] eq_117_in1;
	wire [0:0] eq_117_out;
	eq #(.WIDTH(32)) eq_117(.in0(eq_117_in0), .in1(eq_117_in1), .out(eq_117_out));

	reg [0:0] andOp_118_in0;
	reg [0:0] andOp_118_in1;
	wire [0:0] andOp_118_out;
	andOp #(.WIDTH(1)) andOp_118(.in0(andOp_118_in0), .in1(andOp_118_in1), .out(andOp_118_out));

	reg [31:0] eq_119_in0;
	reg [31:0] eq_119_in1;
	wire [0:0] eq_119_out;
	eq #(.WIDTH(32)) eq_119(.in0(eq_119_in0), .in1(eq_119_in1), .out(eq_119_out));

	reg [0:0] andOp_120_in0;
	reg [0:0] andOp_120_in1;
	wire [0:0] andOp_120_out;
	andOp #(.WIDTH(1)) andOp_120(.in0(andOp_120_in0), .in1(andOp_120_in1), .out(andOp_120_out));

	reg [31:0] eq_121_in0;
	reg [31:0] eq_121_in1;
	wire [0:0] eq_121_out;
	eq #(.WIDTH(32)) eq_121(.in0(eq_121_in0), .in1(eq_121_in1), .out(eq_121_out));

	reg [0:0] andOp_122_in0;
	reg [0:0] andOp_122_in1;
	wire [0:0] andOp_122_out;
	andOp #(.WIDTH(1)) andOp_122(.in0(andOp_122_in0), .in1(andOp_122_in1), .out(andOp_122_out));

	reg [31:0] eq_123_in0;
	reg [31:0] eq_123_in1;
	wire [0:0] eq_123_out;
	eq #(.WIDTH(32)) eq_123(.in0(eq_123_in0), .in1(eq_123_in1), .out(eq_123_out));

	reg [0:0] andOp_124_in0;
	reg [0:0] andOp_124_in1;
	wire [0:0] andOp_124_out;
	andOp #(.WIDTH(1)) andOp_124(.in0(andOp_124_in0), .in1(andOp_124_in1), .out(andOp_124_out));

	reg [31:0] eq_125_in0;
	reg [31:0] eq_125_in1;
	wire [0:0] eq_125_out;
	eq #(.WIDTH(32)) eq_125(.in0(eq_125_in0), .in1(eq_125_in1), .out(eq_125_out));

	reg [0:0] andOp_126_in0;
	reg [0:0] andOp_126_in1;
	wire [0:0] andOp_126_out;
	andOp #(.WIDTH(1)) andOp_126(.in0(andOp_126_in0), .in1(andOp_126_in1), .out(andOp_126_out));

	reg [31:0] eq_127_in0;
	reg [31:0] eq_127_in1;
	wire [0:0] eq_127_out;
	eq #(.WIDTH(32)) eq_127(.in0(eq_127_in0), .in1(eq_127_in1), .out(eq_127_out));

	reg [0:0] andOp_128_in0;
	reg [0:0] andOp_128_in1;
	wire [0:0] andOp_128_out;
	andOp #(.WIDTH(1)) andOp_128(.in0(andOp_128_in0), .in1(andOp_128_in1), .out(andOp_128_out));

	reg [31:0] eq_129_in0;
	reg [31:0] eq_129_in1;
	wire [0:0] eq_129_out;
	eq #(.WIDTH(32)) eq_129(.in0(eq_129_in0), .in1(eq_129_in1), .out(eq_129_out));

	reg [0:0] andOp_130_in0;
	reg [0:0] andOp_130_in1;
	wire [0:0] andOp_130_out;
	andOp #(.WIDTH(1)) andOp_130(.in0(andOp_130_in0), .in1(andOp_130_in1), .out(andOp_130_out));

	reg [31:0] eq_131_in0;
	reg [31:0] eq_131_in1;
	wire [0:0] eq_131_out;
	eq #(.WIDTH(32)) eq_131(.in0(eq_131_in0), .in1(eq_131_in1), .out(eq_131_out));

	reg [0:0] andOp_132_in0;
	reg [0:0] andOp_132_in1;
	wire [0:0] andOp_132_out;
	andOp #(.WIDTH(1)) andOp_132(.in0(andOp_132_in0), .in1(andOp_132_in1), .out(andOp_132_out));

	reg [31:0] eq_133_in0;
	reg [31:0] eq_133_in1;
	wire [0:0] eq_133_out;
	eq #(.WIDTH(32)) eq_133(.in0(eq_133_in0), .in1(eq_133_in1), .out(eq_133_out));

	reg [0:0] andOp_134_in0;
	reg [0:0] andOp_134_in1;
	wire [0:0] andOp_134_out;
	andOp #(.WIDTH(1)) andOp_134(.in0(andOp_134_in0), .in1(andOp_134_in1), .out(andOp_134_out));

	reg [31:0] tmp_output_135_in_data;
	wire [31:0] tmp_output_135_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_135(.in_data(tmp_output_135_in_data), .out_data(tmp_output_135_out_data));

	reg [31:0] eq_136_in0;
	reg [31:0] eq_136_in1;
	wire [0:0] eq_136_out;
	eq #(.WIDTH(32)) eq_136(.in0(eq_136_in0), .in1(eq_136_in1), .out(eq_136_out));

	reg [31:0] eq_137_in0;
	reg [31:0] eq_137_in1;
	wire [0:0] eq_137_out;
	eq #(.WIDTH(32)) eq_137(.in0(eq_137_in0), .in1(eq_137_in1), .out(eq_137_out));

	reg [0:0] andOp_138_in0;
	reg [0:0] andOp_138_in1;
	wire [0:0] andOp_138_out;
	andOp #(.WIDTH(1)) andOp_138(.in0(andOp_138_in0), .in1(andOp_138_in1), .out(andOp_138_out));

	reg [31:0] eq_139_in0;
	reg [31:0] eq_139_in1;
	wire [0:0] eq_139_out;
	eq #(.WIDTH(32)) eq_139(.in0(eq_139_in0), .in1(eq_139_in1), .out(eq_139_out));

	reg [0:0] andOp_140_in0;
	reg [0:0] andOp_140_in1;
	wire [0:0] andOp_140_out;
	andOp #(.WIDTH(1)) andOp_140(.in0(andOp_140_in0), .in1(andOp_140_in1), .out(andOp_140_out));

	reg [31:0] eq_141_in0;
	reg [31:0] eq_141_in1;
	wire [0:0] eq_141_out;
	eq #(.WIDTH(32)) eq_141(.in0(eq_141_in0), .in1(eq_141_in1), .out(eq_141_out));

	reg [0:0] andOp_142_in0;
	reg [0:0] andOp_142_in1;
	wire [0:0] andOp_142_out;
	andOp #(.WIDTH(1)) andOp_142(.in0(andOp_142_in0), .in1(andOp_142_in1), .out(andOp_142_out));

	reg [31:0] eq_143_in0;
	reg [31:0] eq_143_in1;
	wire [0:0] eq_143_out;
	eq #(.WIDTH(32)) eq_143(.in0(eq_143_in0), .in1(eq_143_in1), .out(eq_143_out));

	reg [0:0] andOp_144_in0;
	reg [0:0] andOp_144_in1;
	wire [0:0] andOp_144_out;
	andOp #(.WIDTH(1)) andOp_144(.in0(andOp_144_in0), .in1(andOp_144_in1), .out(andOp_144_out));

	reg [31:0] eq_145_in0;
	reg [31:0] eq_145_in1;
	wire [0:0] eq_145_out;
	eq #(.WIDTH(32)) eq_145(.in0(eq_145_in0), .in1(eq_145_in1), .out(eq_145_out));

	reg [0:0] andOp_146_in0;
	reg [0:0] andOp_146_in1;
	wire [0:0] andOp_146_out;
	andOp #(.WIDTH(1)) andOp_146(.in0(andOp_146_in0), .in1(andOp_146_in1), .out(andOp_146_out));

	reg [31:0] eq_147_in0;
	reg [31:0] eq_147_in1;
	wire [0:0] eq_147_out;
	eq #(.WIDTH(32)) eq_147(.in0(eq_147_in0), .in1(eq_147_in1), .out(eq_147_out));

	reg [0:0] andOp_148_in0;
	reg [0:0] andOp_148_in1;
	wire [0:0] andOp_148_out;
	andOp #(.WIDTH(1)) andOp_148(.in0(andOp_148_in0), .in1(andOp_148_in1), .out(andOp_148_out));

	reg [31:0] eq_149_in0;
	reg [31:0] eq_149_in1;
	wire [0:0] eq_149_out;
	eq #(.WIDTH(32)) eq_149(.in0(eq_149_in0), .in1(eq_149_in1), .out(eq_149_out));

	reg [0:0] andOp_150_in0;
	reg [0:0] andOp_150_in1;
	wire [0:0] andOp_150_out;
	andOp #(.WIDTH(1)) andOp_150(.in0(andOp_150_in0), .in1(andOp_150_in1), .out(andOp_150_out));

	reg [31:0] eq_151_in0;
	reg [31:0] eq_151_in1;
	wire [0:0] eq_151_out;
	eq #(.WIDTH(32)) eq_151(.in0(eq_151_in0), .in1(eq_151_in1), .out(eq_151_out));

	reg [0:0] andOp_152_in0;
	reg [0:0] andOp_152_in1;
	wire [0:0] andOp_152_out;
	andOp #(.WIDTH(1)) andOp_152(.in0(andOp_152_in0), .in1(andOp_152_in1), .out(andOp_152_out));

	reg [31:0] eq_153_in0;
	reg [31:0] eq_153_in1;
	wire [0:0] eq_153_out;
	eq #(.WIDTH(32)) eq_153(.in0(eq_153_in0), .in1(eq_153_in1), .out(eq_153_out));

	reg [0:0] andOp_154_in0;
	reg [0:0] andOp_154_in1;
	wire [0:0] andOp_154_out;
	andOp #(.WIDTH(1)) andOp_154(.in0(andOp_154_in0), .in1(andOp_154_in1), .out(andOp_154_out));

	reg [0:0] notOp_155_in0;
	wire [0:0] notOp_155_out;
	notOp #(.WIDTH(1)) notOp_155(.in(notOp_155_in0), .out(notOp_155_out));

	reg [0:0] andOp_156_in0;
	reg [0:0] andOp_156_in1;
	wire [0:0] andOp_156_out;
	andOp #(.WIDTH(1)) andOp_156(.in0(andOp_156_in0), .in1(andOp_156_in1), .out(andOp_156_out));

	reg [31:0] eq_157_in0;
	reg [31:0] eq_157_in1;
	wire [0:0] eq_157_out;
	eq #(.WIDTH(32)) eq_157(.in0(eq_157_in0), .in1(eq_157_in1), .out(eq_157_out));

	reg [0:0] andOp_158_in0;
	reg [0:0] andOp_158_in1;
	wire [0:0] andOp_158_out;
	andOp #(.WIDTH(1)) andOp_158(.in0(andOp_158_in0), .in1(andOp_158_in1), .out(andOp_158_out));

	reg [31:0] eq_159_in0;
	reg [31:0] eq_159_in1;
	wire [0:0] eq_159_out;
	eq #(.WIDTH(32)) eq_159(.in0(eq_159_in0), .in1(eq_159_in1), .out(eq_159_out));

	reg [0:0] andOp_160_in0;
	reg [0:0] andOp_160_in1;
	wire [0:0] andOp_160_out;
	andOp #(.WIDTH(1)) andOp_160(.in0(andOp_160_in0), .in1(andOp_160_in1), .out(andOp_160_out));

	reg [0:0] notOp_161_in0;
	wire [0:0] notOp_161_out;
	notOp #(.WIDTH(1)) notOp_161(.in(notOp_161_in0), .out(notOp_161_out));

	reg [0:0] andOp_162_in0;
	reg [0:0] andOp_162_in1;
	wire [0:0] andOp_162_out;
	andOp #(.WIDTH(1)) andOp_162(.in0(andOp_162_in0), .in1(andOp_162_in1), .out(andOp_162_out));

	reg [31:0] eq_163_in0;
	reg [31:0] eq_163_in1;
	wire [0:0] eq_163_out;
	eq #(.WIDTH(32)) eq_163(.in0(eq_163_in0), .in1(eq_163_in1), .out(eq_163_out));

	reg [0:0] andOp_164_in0;
	reg [0:0] andOp_164_in1;
	wire [0:0] andOp_164_out;
	andOp #(.WIDTH(1)) andOp_164(.in0(andOp_164_in0), .in1(andOp_164_in1), .out(andOp_164_out));

	reg [31:0] eq_165_in0;
	reg [31:0] eq_165_in1;
	wire [0:0] eq_165_out;
	eq #(.WIDTH(32)) eq_165(.in0(eq_165_in0), .in1(eq_165_in1), .out(eq_165_out));

	reg [0:0] andOp_166_in0;
	reg [0:0] andOp_166_in1;
	wire [0:0] andOp_166_out;
	andOp #(.WIDTH(1)) andOp_166(.in0(andOp_166_in0), .in1(andOp_166_in1), .out(andOp_166_out));

	reg [0:0] notOp_167_in0;
	wire [0:0] notOp_167_out;
	notOp #(.WIDTH(1)) notOp_167(.in(notOp_167_in0), .out(notOp_167_out));

	reg [0:0] andOp_168_in0;
	reg [0:0] andOp_168_in1;
	wire [0:0] andOp_168_out;
	andOp #(.WIDTH(1)) andOp_168(.in0(andOp_168_in0), .in1(andOp_168_in1), .out(andOp_168_out));

	reg [31:0] eq_169_in0;
	reg [31:0] eq_169_in1;
	wire [0:0] eq_169_out;
	eq #(.WIDTH(32)) eq_169(.in0(eq_169_in0), .in1(eq_169_in1), .out(eq_169_out));

	reg [0:0] andOp_170_in0;
	reg [0:0] andOp_170_in1;
	wire [0:0] andOp_170_out;
	andOp #(.WIDTH(1)) andOp_170(.in0(andOp_170_in0), .in1(andOp_170_in1), .out(andOp_170_out));

	reg [31:0] eq_171_in0;
	reg [31:0] eq_171_in1;
	wire [0:0] eq_171_out;
	eq #(.WIDTH(32)) eq_171(.in0(eq_171_in0), .in1(eq_171_in1), .out(eq_171_out));

	reg [0:0] andOp_172_in0;
	reg [0:0] andOp_172_in1;
	wire [0:0] andOp_172_out;
	andOp #(.WIDTH(1)) andOp_172(.in0(andOp_172_in0), .in1(andOp_172_in1), .out(andOp_172_out));

	reg [0:0] notOp_173_in0;
	wire [0:0] notOp_173_out;
	notOp #(.WIDTH(1)) notOp_173(.in(notOp_173_in0), .out(notOp_173_out));

	reg [0:0] andOp_174_in0;
	reg [0:0] andOp_174_in1;
	wire [0:0] andOp_174_out;
	andOp #(.WIDTH(1)) andOp_174(.in0(andOp_174_in0), .in1(andOp_174_in1), .out(andOp_174_out));

	reg [31:0] eq_175_in0;
	reg [31:0] eq_175_in1;
	wire [0:0] eq_175_out;
	eq #(.WIDTH(32)) eq_175(.in0(eq_175_in0), .in1(eq_175_in1), .out(eq_175_out));

	reg [0:0] andOp_176_in0;
	reg [0:0] andOp_176_in1;
	wire [0:0] andOp_176_out;
	andOp #(.WIDTH(1)) andOp_176(.in0(andOp_176_in0), .in1(andOp_176_in1), .out(andOp_176_out));

	reg [31:0] eq_177_in0;
	reg [31:0] eq_177_in1;
	wire [0:0] eq_177_out;
	eq #(.WIDTH(32)) eq_177(.in0(eq_177_in0), .in1(eq_177_in1), .out(eq_177_out));

	reg [0:0] andOp_178_in0;
	reg [0:0] andOp_178_in1;
	wire [0:0] andOp_178_out;
	andOp #(.WIDTH(1)) andOp_178(.in0(andOp_178_in0), .in1(andOp_178_in1), .out(andOp_178_out));

	reg [0:0] notOp_179_in0;
	wire [0:0] notOp_179_out;
	notOp #(.WIDTH(1)) notOp_179(.in(notOp_179_in0), .out(notOp_179_out));

	reg [0:0] andOp_180_in0;
	reg [0:0] andOp_180_in1;
	wire [0:0] andOp_180_out;
	andOp #(.WIDTH(1)) andOp_180(.in0(andOp_180_in0), .in1(andOp_180_in1), .out(andOp_180_out));

	reg [31:0] eq_181_in0;
	reg [31:0] eq_181_in1;
	wire [0:0] eq_181_out;
	eq #(.WIDTH(32)) eq_181(.in0(eq_181_in0), .in1(eq_181_in1), .out(eq_181_out));

	reg [0:0] andOp_182_in0;
	reg [0:0] andOp_182_in1;
	wire [0:0] andOp_182_out;
	andOp #(.WIDTH(1)) andOp_182(.in0(andOp_182_in0), .in1(andOp_182_in1), .out(andOp_182_out));

	reg [31:0] eq_183_in0;
	reg [31:0] eq_183_in1;
	wire [0:0] eq_183_out;
	eq #(.WIDTH(32)) eq_183(.in0(eq_183_in0), .in1(eq_183_in1), .out(eq_183_out));

	reg [0:0] andOp_184_in0;
	reg [0:0] andOp_184_in1;
	wire [0:0] andOp_184_out;
	andOp #(.WIDTH(1)) andOp_184(.in0(andOp_184_in0), .in1(andOp_184_in1), .out(andOp_184_out));

	reg [0:0] notOp_185_in0;
	wire [0:0] notOp_185_out;
	notOp #(.WIDTH(1)) notOp_185(.in(notOp_185_in0), .out(notOp_185_out));

	reg [0:0] andOp_186_in0;
	reg [0:0] andOp_186_in1;
	wire [0:0] andOp_186_out;
	andOp #(.WIDTH(1)) andOp_186(.in0(andOp_186_in0), .in1(andOp_186_in1), .out(andOp_186_out));

	reg [31:0] eq_187_in0;
	reg [31:0] eq_187_in1;
	wire [0:0] eq_187_out;
	eq #(.WIDTH(32)) eq_187(.in0(eq_187_in0), .in1(eq_187_in1), .out(eq_187_out));

	reg [0:0] andOp_188_in0;
	reg [0:0] andOp_188_in1;
	wire [0:0] andOp_188_out;
	andOp #(.WIDTH(1)) andOp_188(.in0(andOp_188_in0), .in1(andOp_188_in1), .out(andOp_188_out));

	reg [0:0] notOp_189_in0;
	wire [0:0] notOp_189_out;
	notOp #(.WIDTH(1)) notOp_189(.in(notOp_189_in0), .out(notOp_189_out));

	reg [0:0] andOp_190_in0;
	reg [0:0] andOp_190_in1;
	wire [0:0] andOp_190_out;
	andOp #(.WIDTH(1)) andOp_190(.in0(andOp_190_in0), .in1(andOp_190_in1), .out(andOp_190_out));

	reg [31:0] eq_191_in0;
	reg [31:0] eq_191_in1;
	wire [0:0] eq_191_out;
	eq #(.WIDTH(32)) eq_191(.in0(eq_191_in0), .in1(eq_191_in1), .out(eq_191_out));

	reg [0:0] andOp_192_in0;
	reg [0:0] andOp_192_in1;
	wire [0:0] andOp_192_out;
	andOp #(.WIDTH(1)) andOp_192(.in0(andOp_192_in0), .in1(andOp_192_in1), .out(andOp_192_out));

	reg [31:0] eq_193_in0;
	reg [31:0] eq_193_in1;
	wire [0:0] eq_193_out;
	eq #(.WIDTH(32)) eq_193(.in0(eq_193_in0), .in1(eq_193_in1), .out(eq_193_out));

	reg [0:0] andOp_194_in0;
	reg [0:0] andOp_194_in1;
	wire [0:0] andOp_194_out;
	andOp #(.WIDTH(1)) andOp_194(.in0(andOp_194_in0), .in1(andOp_194_in1), .out(andOp_194_out));

	reg [0:0] notOp_195_in0;
	wire [0:0] notOp_195_out;
	notOp #(.WIDTH(1)) notOp_195(.in(notOp_195_in0), .out(notOp_195_out));

	reg [0:0] andOp_196_in0;
	reg [0:0] andOp_196_in1;
	wire [0:0] andOp_196_out;
	andOp #(.WIDTH(1)) andOp_196(.in0(andOp_196_in0), .in1(andOp_196_in1), .out(andOp_196_out));

	reg [31:0] eq_197_in0;
	reg [31:0] eq_197_in1;
	wire [0:0] eq_197_out;
	eq #(.WIDTH(32)) eq_197(.in0(eq_197_in0), .in1(eq_197_in1), .out(eq_197_out));

	reg [0:0] andOp_198_in0;
	reg [0:0] andOp_198_in1;
	wire [0:0] andOp_198_out;
	andOp #(.WIDTH(1)) andOp_198(.in0(andOp_198_in0), .in1(andOp_198_in1), .out(andOp_198_out));

	reg [31:0] eq_199_in0;
	reg [31:0] eq_199_in1;
	wire [0:0] eq_199_out;
	eq #(.WIDTH(32)) eq_199(.in0(eq_199_in0), .in1(eq_199_in1), .out(eq_199_out));

	reg [0:0] andOp_200_in0;
	reg [0:0] andOp_200_in1;
	wire [0:0] andOp_200_out;
	andOp #(.WIDTH(1)) andOp_200(.in0(andOp_200_in0), .in1(andOp_200_in1), .out(andOp_200_out));

	reg [31:0] eq_201_in0;
	reg [31:0] eq_201_in1;
	wire [0:0] eq_201_out;
	eq #(.WIDTH(32)) eq_201(.in0(eq_201_in0), .in1(eq_201_in1), .out(eq_201_out));

	reg [0:0] andOp_202_in0;
	reg [0:0] andOp_202_in1;
	wire [0:0] andOp_202_out;
	andOp #(.WIDTH(1)) andOp_202(.in0(andOp_202_in0), .in1(andOp_202_in1), .out(andOp_202_out));

	reg [0:0] notOp_203_in0;
	wire [0:0] notOp_203_out;
	notOp #(.WIDTH(1)) notOp_203(.in(notOp_203_in0), .out(notOp_203_out));

	reg [0:0] andOp_204_in0;
	reg [0:0] andOp_204_in1;
	wire [0:0] andOp_204_out;
	andOp #(.WIDTH(1)) andOp_204(.in0(andOp_204_in0), .in1(andOp_204_in1), .out(andOp_204_out));

	reg [31:0] eq_205_in0;
	reg [31:0] eq_205_in1;
	wire [0:0] eq_205_out;
	eq #(.WIDTH(32)) eq_205(.in0(eq_205_in0), .in1(eq_205_in1), .out(eq_205_out));

	reg [0:0] andOp_206_in0;
	reg [0:0] andOp_206_in1;
	wire [0:0] andOp_206_out;
	andOp #(.WIDTH(1)) andOp_206(.in0(andOp_206_in0), .in1(andOp_206_in1), .out(andOp_206_out));

	reg [31:0] eq_207_in0;
	reg [31:0] eq_207_in1;
	wire [0:0] eq_207_out;
	eq #(.WIDTH(32)) eq_207(.in0(eq_207_in0), .in1(eq_207_in1), .out(eq_207_out));

	reg [0:0] andOp_208_in0;
	reg [0:0] andOp_208_in1;
	wire [0:0] andOp_208_out;
	andOp #(.WIDTH(1)) andOp_208(.in0(andOp_208_in0), .in1(andOp_208_in1), .out(andOp_208_out));

	reg [0:0] notOp_209_in0;
	wire [0:0] notOp_209_out;
	notOp #(.WIDTH(1)) notOp_209(.in(notOp_209_in0), .out(notOp_209_out));

	reg [0:0] andOp_210_in0;
	reg [0:0] andOp_210_in1;
	wire [0:0] andOp_210_out;
	andOp #(.WIDTH(1)) andOp_210(.in0(andOp_210_in0), .in1(andOp_210_in1), .out(andOp_210_out));

	reg [31:0] eq_211_in0;
	reg [31:0] eq_211_in1;
	wire [0:0] eq_211_out;
	eq #(.WIDTH(32)) eq_211(.in0(eq_211_in0), .in1(eq_211_in1), .out(eq_211_out));

	reg [0:0] andOp_212_in0;
	reg [0:0] andOp_212_in1;
	wire [0:0] andOp_212_out;
	andOp #(.WIDTH(1)) andOp_212(.in0(andOp_212_in0), .in1(andOp_212_in1), .out(andOp_212_out));

	reg [31:0] eq_213_in0;
	reg [31:0] eq_213_in1;
	wire [0:0] eq_213_out;
	eq #(.WIDTH(32)) eq_213(.in0(eq_213_in0), .in1(eq_213_in1), .out(eq_213_out));

	reg [0:0] andOp_214_in0;
	reg [0:0] andOp_214_in1;
	wire [0:0] andOp_214_out;
	andOp #(.WIDTH(1)) andOp_214(.in0(andOp_214_in0), .in1(andOp_214_in1), .out(andOp_214_out));

	reg [0:0] notOp_215_in0;
	wire [0:0] notOp_215_out;
	notOp #(.WIDTH(1)) notOp_215(.in(notOp_215_in0), .out(notOp_215_out));

	reg [0:0] andOp_216_in0;
	reg [0:0] andOp_216_in1;
	wire [0:0] andOp_216_out;
	andOp #(.WIDTH(1)) andOp_216(.in0(andOp_216_in0), .in1(andOp_216_in1), .out(andOp_216_out));

	reg [31:0] eq_217_in0;
	reg [31:0] eq_217_in1;
	wire [0:0] eq_217_out;
	eq #(.WIDTH(32)) eq_217(.in0(eq_217_in0), .in1(eq_217_in1), .out(eq_217_out));

	reg [0:0] andOp_218_in0;
	reg [0:0] andOp_218_in1;
	wire [0:0] andOp_218_out;
	andOp #(.WIDTH(1)) andOp_218(.in0(andOp_218_in0), .in1(andOp_218_in1), .out(andOp_218_out));

	reg [0:0] andOp_219_in0;
	reg [0:0] andOp_219_in1;
	wire [0:0] andOp_219_out;
	andOp #(.WIDTH(1)) andOp_219(.in0(andOp_219_in0), .in1(andOp_219_in1), .out(andOp_219_out));

	reg [31:0] eq_220_in0;
	reg [31:0] eq_220_in1;
	wire [0:0] eq_220_out;
	eq #(.WIDTH(32)) eq_220(.in0(eq_220_in0), .in1(eq_220_in1), .out(eq_220_out));

	reg [0:0] andOp_221_in0;
	reg [0:0] andOp_221_in1;
	wire [0:0] andOp_221_out;
	andOp #(.WIDTH(1)) andOp_221(.in0(andOp_221_in0), .in1(andOp_221_in1), .out(andOp_221_out));

	reg [0:0] notOp_222_in0;
	wire [0:0] notOp_222_out;
	notOp #(.WIDTH(1)) notOp_222(.in(notOp_222_in0), .out(notOp_222_out));

	reg [31:0] eq_223_in0;
	reg [31:0] eq_223_in1;
	wire [0:0] eq_223_out;
	eq #(.WIDTH(32)) eq_223(.in0(eq_223_in0), .in1(eq_223_in1), .out(eq_223_out));

	reg [0:0] andOp_224_in0;
	reg [0:0] andOp_224_in1;
	wire [0:0] andOp_224_out;
	andOp #(.WIDTH(1)) andOp_224(.in0(andOp_224_in0), .in1(andOp_224_in1), .out(andOp_224_out));

	reg [0:0] andOp_225_in0;
	reg [0:0] andOp_225_in1;
	wire [0:0] andOp_225_out;
	andOp #(.WIDTH(1)) andOp_225(.in0(andOp_225_in0), .in1(andOp_225_in1), .out(andOp_225_out));

	reg [31:0] eq_226_in0;
	reg [31:0] eq_226_in1;
	wire [0:0] eq_226_out;
	eq #(.WIDTH(32)) eq_226(.in0(eq_226_in0), .in1(eq_226_in1), .out(eq_226_out));

	reg [0:0] andOp_227_in0;
	reg [0:0] andOp_227_in1;
	wire [0:0] andOp_227_out;
	andOp #(.WIDTH(1)) andOp_227(.in0(andOp_227_in0), .in1(andOp_227_in1), .out(andOp_227_out));

	reg [31:0] eq_228_in0;
	reg [31:0] eq_228_in1;
	wire [0:0] eq_228_out;
	eq #(.WIDTH(32)) eq_228(.in0(eq_228_in0), .in1(eq_228_in1), .out(eq_228_out));

	reg [0:0] andOp_229_in0;
	reg [0:0] andOp_229_in1;
	wire [0:0] andOp_229_out;
	andOp #(.WIDTH(1)) andOp_229(.in0(andOp_229_in0), .in1(andOp_229_in1), .out(andOp_229_out));

	reg [0:0] andOp_230_in0;
	reg [0:0] andOp_230_in1;
	wire [0:0] andOp_230_out;
	andOp #(.WIDTH(1)) andOp_230(.in0(andOp_230_in0), .in1(andOp_230_in1), .out(andOp_230_out));

	reg [31:0] eq_231_in0;
	reg [31:0] eq_231_in1;
	wire [0:0] eq_231_out;
	eq #(.WIDTH(32)) eq_231(.in0(eq_231_in0), .in1(eq_231_in1), .out(eq_231_out));

	reg [0:0] andOp_232_in0;
	reg [0:0] andOp_232_in1;
	wire [0:0] andOp_232_out;
	andOp #(.WIDTH(1)) andOp_232(.in0(andOp_232_in0), .in1(andOp_232_in1), .out(andOp_232_out));

	reg [31:0] eq_233_in0;
	reg [31:0] eq_233_in1;
	wire [0:0] eq_233_out;
	eq #(.WIDTH(32)) eq_233(.in0(eq_233_in0), .in1(eq_233_in1), .out(eq_233_out));

	reg [0:0] andOp_234_in0;
	reg [0:0] andOp_234_in1;
	wire [0:0] andOp_234_out;
	andOp #(.WIDTH(1)) andOp_234(.in0(andOp_234_in0), .in1(andOp_234_in1), .out(andOp_234_out));

	reg [0:0] andOp_235_in0;
	reg [0:0] andOp_235_in1;
	wire [0:0] andOp_235_out;
	andOp #(.WIDTH(1)) andOp_235(.in0(andOp_235_in0), .in1(andOp_235_in1), .out(andOp_235_out));

	reg [31:0] eq_236_in0;
	reg [31:0] eq_236_in1;
	wire [0:0] eq_236_out;
	eq #(.WIDTH(32)) eq_236(.in0(eq_236_in0), .in1(eq_236_in1), .out(eq_236_out));

	reg [0:0] andOp_237_in0;
	reg [0:0] andOp_237_in1;
	wire [0:0] andOp_237_out;
	andOp #(.WIDTH(1)) andOp_237(.in0(andOp_237_in0), .in1(andOp_237_in1), .out(andOp_237_out));

	reg [31:0] eq_238_in0;
	reg [31:0] eq_238_in1;
	wire [0:0] eq_238_out;
	eq #(.WIDTH(32)) eq_238(.in0(eq_238_in0), .in1(eq_238_in1), .out(eq_238_out));

	reg [0:0] andOp_239_in0;
	reg [0:0] andOp_239_in1;
	wire [0:0] andOp_239_out;
	andOp #(.WIDTH(1)) andOp_239(.in0(andOp_239_in0), .in1(andOp_239_in1), .out(andOp_239_out));

	reg [0:0] andOp_240_in0;
	reg [0:0] andOp_240_in1;
	wire [0:0] andOp_240_out;
	andOp #(.WIDTH(1)) andOp_240(.in0(andOp_240_in0), .in1(andOp_240_in1), .out(andOp_240_out));

	reg [31:0] eq_241_in0;
	reg [31:0] eq_241_in1;
	wire [0:0] eq_241_out;
	eq #(.WIDTH(32)) eq_241(.in0(eq_241_in0), .in1(eq_241_in1), .out(eq_241_out));

	reg [0:0] andOp_242_in0;
	reg [0:0] andOp_242_in1;
	wire [0:0] andOp_242_out;
	andOp #(.WIDTH(1)) andOp_242(.in0(andOp_242_in0), .in1(andOp_242_in1), .out(andOp_242_out));

	reg [0:0] notOp_243_in0;
	wire [0:0] notOp_243_out;
	notOp #(.WIDTH(1)) notOp_243(.in(notOp_243_in0), .out(notOp_243_out));

	reg [31:0] eq_244_in0;
	reg [31:0] eq_244_in1;
	wire [0:0] eq_244_out;
	eq #(.WIDTH(32)) eq_244(.in0(eq_244_in0), .in1(eq_244_in1), .out(eq_244_out));

	reg [0:0] andOp_245_in0;
	reg [0:0] andOp_245_in1;
	wire [0:0] andOp_245_out;
	andOp #(.WIDTH(1)) andOp_245(.in0(andOp_245_in0), .in1(andOp_245_in1), .out(andOp_245_out));

	reg [0:0] andOp_246_in0;
	reg [0:0] andOp_246_in1;
	wire [0:0] andOp_246_out;
	andOp #(.WIDTH(1)) andOp_246(.in0(andOp_246_in0), .in1(andOp_246_in1), .out(andOp_246_out));

	reg [31:0] eq_247_in0;
	reg [31:0] eq_247_in1;
	wire [0:0] eq_247_out;
	eq #(.WIDTH(32)) eq_247(.in0(eq_247_in0), .in1(eq_247_in1), .out(eq_247_out));

	reg [0:0] andOp_248_in0;
	reg [0:0] andOp_248_in1;
	wire [0:0] andOp_248_out;
	andOp #(.WIDTH(1)) andOp_248(.in0(andOp_248_in0), .in1(andOp_248_in1), .out(andOp_248_out));

	reg [0:0] notOp_249_in0;
	wire [0:0] notOp_249_out;
	notOp #(.WIDTH(1)) notOp_249(.in(notOp_249_in0), .out(notOp_249_out));

	reg [31:0] eq_250_in0;
	reg [31:0] eq_250_in1;
	wire [0:0] eq_250_out;
	eq #(.WIDTH(32)) eq_250(.in0(eq_250_in0), .in1(eq_250_in1), .out(eq_250_out));

	reg [0:0] andOp_251_in0;
	reg [0:0] andOp_251_in1;
	wire [0:0] andOp_251_out;
	andOp #(.WIDTH(1)) andOp_251(.in0(andOp_251_in0), .in1(andOp_251_in1), .out(andOp_251_out));

	reg [0:0] andOp_252_in0;
	reg [0:0] andOp_252_in1;
	wire [0:0] andOp_252_out;
	andOp #(.WIDTH(1)) andOp_252(.in0(andOp_252_in0), .in1(andOp_252_in1), .out(andOp_252_out));

	reg [31:0] eq_253_in0;
	reg [31:0] eq_253_in1;
	wire [0:0] eq_253_out;
	eq #(.WIDTH(32)) eq_253(.in0(eq_253_in0), .in1(eq_253_in1), .out(eq_253_out));

	reg [0:0] andOp_254_in0;
	reg [0:0] andOp_254_in1;
	wire [0:0] andOp_254_out;
	andOp #(.WIDTH(1)) andOp_254(.in0(andOp_254_in0), .in1(andOp_254_in1), .out(andOp_254_out));

	reg [31:0] eq_255_in0;
	reg [31:0] eq_255_in1;
	wire [0:0] eq_255_out;
	eq #(.WIDTH(32)) eq_255(.in0(eq_255_in0), .in1(eq_255_in1), .out(eq_255_out));

	reg [0:0] andOp_256_in0;
	reg [0:0] andOp_256_in1;
	wire [0:0] andOp_256_out;
	andOp #(.WIDTH(1)) andOp_256(.in0(andOp_256_in0), .in1(andOp_256_in1), .out(andOp_256_out));

	reg [0:0] andOp_257_in0;
	reg [0:0] andOp_257_in1;
	wire [0:0] andOp_257_out;
	andOp #(.WIDTH(1)) andOp_257(.in0(andOp_257_in0), .in1(andOp_257_in1), .out(andOp_257_out));

	reg [31:0] eq_258_in0;
	reg [31:0] eq_258_in1;
	wire [0:0] eq_258_out;
	eq #(.WIDTH(32)) eq_258(.in0(eq_258_in0), .in1(eq_258_in1), .out(eq_258_out));

	reg [0:0] andOp_259_in0;
	reg [0:0] andOp_259_in1;
	wire [0:0] andOp_259_out;
	andOp #(.WIDTH(1)) andOp_259(.in0(andOp_259_in0), .in1(andOp_259_in1), .out(andOp_259_out));

	reg [31:0] eq_260_in0;
	reg [31:0] eq_260_in1;
	wire [0:0] eq_260_out;
	eq #(.WIDTH(32)) eq_260(.in0(eq_260_in0), .in1(eq_260_in1), .out(eq_260_out));

	reg [0:0] andOp_261_in0;
	reg [0:0] andOp_261_in1;
	wire [0:0] andOp_261_out;
	andOp #(.WIDTH(1)) andOp_261(.in0(andOp_261_in0), .in1(andOp_261_in1), .out(andOp_261_out));

	reg [31:0] eq_262_in0;
	reg [31:0] eq_262_in1;
	wire [0:0] eq_262_out;
	eq #(.WIDTH(32)) eq_262(.in0(eq_262_in0), .in1(eq_262_in1), .out(eq_262_out));

	reg [0:0] andOp_263_in0;
	reg [0:0] andOp_263_in1;
	wire [0:0] andOp_263_out;
	andOp #(.WIDTH(1)) andOp_263(.in0(andOp_263_in0), .in1(andOp_263_in1), .out(andOp_263_out));

	reg [31:0] eq_264_in0;
	reg [31:0] eq_264_in1;
	wire [0:0] eq_264_out;
	eq #(.WIDTH(32)) eq_264(.in0(eq_264_in0), .in1(eq_264_in1), .out(eq_264_out));

	reg [0:0] andOp_265_in0;
	reg [0:0] andOp_265_in1;
	wire [0:0] andOp_265_out;
	andOp #(.WIDTH(1)) andOp_265(.in0(andOp_265_in0), .in1(andOp_265_in1), .out(andOp_265_out));

	reg [31:0] eq_266_in0;
	reg [31:0] eq_266_in1;
	wire [0:0] eq_266_out;
	eq #(.WIDTH(32)) eq_266(.in0(eq_266_in0), .in1(eq_266_in1), .out(eq_266_out));

	reg [0:0] andOp_267_in0;
	reg [0:0] andOp_267_in1;
	wire [0:0] andOp_267_out;
	andOp #(.WIDTH(1)) andOp_267(.in0(andOp_267_in0), .in1(andOp_267_in1), .out(andOp_267_out));

	// End Functional Units

	reg [31:0] add_tmp_4;
	reg [31:0] call_tmp_6;
	reg [31:0] global_next_block;
	reg [31:0] global_state;
	reg [0:0] icmp_tmp_5;
	reg [31:0] last_BB_reg;
	reg [31:0] phi_tmp_0;

	// controller for add_add_12.add_in0_add_12
	// controller for add_add_12.add_in1_add_12
	// Insensitive connections
	always @(*) begin
		add_in0_add_12 = valid ? rdata_ram_0 : rdata_ram_0;
		add_in1_add_12 = valid ? tmp_output_135_out_data : tmp_output_135_out_data;
	end
	// controller for add_add_14.add_in0_add_14
	// controller for add_add_14.add_in1_add_14
	// Insensitive connections
	always @(*) begin
		add_in0_add_14 = valid ? phi_tmp_0 : phi_tmp_0;
		add_in1_add_14 = valid ? 32'd1 : 32'd1;
	end
	// controller for andOp_1.andOp_1_in0
	// controller for andOp_1.andOp_1_in1
	// Insensitive connections
	always @(*) begin
		andOp_1_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_1_in1 = valid ? eq_0_out : eq_0_out;
	end
	// controller for andOp_10.andOp_10_in0
	// controller for andOp_10.andOp_10_in1
	// Insensitive connections
	always @(*) begin
		andOp_10_in0 = valid ? andOp_9_out : andOp_9_out;
		andOp_10_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_101.andOp_101_in0
	// controller for andOp_101.andOp_101_in1
	// Insensitive connections
	always @(*) begin
		andOp_101_in0 = valid ? notOp_100_out : notOp_100_out;
		andOp_101_in1 = valid ? andOp_27_out : andOp_27_out;
	end
	// controller for andOp_104.andOp_104_in0
	// controller for andOp_104.andOp_104_in1
	// Insensitive connections
	always @(*) begin
		andOp_104_in0 = valid ? notOp_103_out : notOp_103_out;
		andOp_104_in1 = valid ? andOp_10_out : andOp_10_out;
	end
	// controller for andOp_107.andOp_107_in0
	// controller for andOp_107.andOp_107_in1
	// Insensitive connections
	always @(*) begin
		andOp_107_in0 = valid ? notOp_106_out : notOp_106_out;
		andOp_107_in1 = valid ? andOp_36_out : andOp_36_out;
	end
	// controller for andOp_110.andOp_110_in0
	// controller for andOp_110.andOp_110_in1
	// Insensitive connections
	always @(*) begin
		andOp_110_in0 = valid ? notOp_109_out : notOp_109_out;
		andOp_110_in1 = valid ? andOp_42_out : andOp_42_out;
	end
	// controller for andOp_112.andOp_112_in0
	// controller for andOp_112.andOp_112_in1
	// Insensitive connections
	always @(*) begin
		andOp_112_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_112_in1 = valid ? eq_111_out : eq_111_out;
	end
	// controller for andOp_114.andOp_114_in0
	// controller for andOp_114.andOp_114_in1
	// Insensitive connections
	always @(*) begin
		andOp_114_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_114_in1 = valid ? eq_113_out : eq_113_out;
	end
	// controller for andOp_116.andOp_116_in0
	// controller for andOp_116.andOp_116_in1
	// Insensitive connections
	always @(*) begin
		andOp_116_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_116_in1 = valid ? eq_115_out : eq_115_out;
	end
	// controller for andOp_118.andOp_118_in0
	// controller for andOp_118.andOp_118_in1
	// Insensitive connections
	always @(*) begin
		andOp_118_in0 = valid ? bb_7_active_out_data : bb_7_active_out_data;
		andOp_118_in1 = valid ? eq_117_out : eq_117_out;
	end
	// controller for andOp_120.andOp_120_in0
	// controller for andOp_120.andOp_120_in1
	// Insensitive connections
	always @(*) begin
		andOp_120_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_120_in1 = valid ? eq_119_out : eq_119_out;
	end
	// controller for andOp_122.andOp_122_in0
	// controller for andOp_122.andOp_122_in1
	// Insensitive connections
	always @(*) begin
		andOp_122_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_122_in1 = valid ? eq_121_out : eq_121_out;
	end
	// controller for andOp_124.andOp_124_in0
	// controller for andOp_124.andOp_124_in1
	// Insensitive connections
	always @(*) begin
		andOp_124_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_124_in1 = valid ? eq_123_out : eq_123_out;
	end
	// controller for andOp_126.andOp_126_in0
	// controller for andOp_126.andOp_126_in1
	// Insensitive connections
	always @(*) begin
		andOp_126_in0 = valid ? bb_3_active_out_data : bb_3_active_out_data;
		andOp_126_in1 = valid ? eq_125_out : eq_125_out;
	end
	// controller for andOp_128.andOp_128_in0
	// controller for andOp_128.andOp_128_in1
	// Insensitive connections
	always @(*) begin
		andOp_128_in0 = valid ? bb_9_active_out_data : bb_9_active_out_data;
		andOp_128_in1 = valid ? eq_127_out : eq_127_out;
	end
	// controller for andOp_13.andOp_13_in0
	// controller for andOp_13.andOp_13_in1
	// Insensitive connections
	always @(*) begin
		andOp_13_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_13_in1 = valid ? eq_12_out : eq_12_out;
	end
	// controller for andOp_130.andOp_130_in0
	// controller for andOp_130.andOp_130_in1
	// Insensitive connections
	always @(*) begin
		andOp_130_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_130_in1 = valid ? eq_129_out : eq_129_out;
	end
	// controller for andOp_132.andOp_132_in0
	// controller for andOp_132.andOp_132_in1
	// Insensitive connections
	always @(*) begin
		andOp_132_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_132_in1 = valid ? eq_131_out : eq_131_out;
	end
	// controller for andOp_134.andOp_134_in0
	// controller for andOp_134.andOp_134_in1
	// Insensitive connections
	always @(*) begin
		andOp_134_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_134_in1 = valid ? eq_133_out : eq_133_out;
	end
	// controller for andOp_138.andOp_138_in0
	// controller for andOp_138.andOp_138_in1
	// Insensitive connections
	always @(*) begin
		andOp_138_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_138_in1 = valid ? eq_137_out : eq_137_out;
	end
	// controller for andOp_14.andOp_14_in0
	// controller for andOp_14.andOp_14_in1
	// Insensitive connections
	always @(*) begin
		andOp_14_in0 = valid ? andOp_13_out : andOp_13_out;
		andOp_14_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_140.andOp_140_in0
	// controller for andOp_140.andOp_140_in1
	// Insensitive connections
	always @(*) begin
		andOp_140_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_140_in1 = valid ? eq_139_out : eq_139_out;
	end
	// controller for andOp_142.andOp_142_in0
	// controller for andOp_142.andOp_142_in1
	// Insensitive connections
	always @(*) begin
		andOp_142_in0 = valid ? bb_2_active_out_data : bb_2_active_out_data;
		andOp_142_in1 = valid ? eq_141_out : eq_141_out;
	end
	// controller for andOp_144.andOp_144_in0
	// controller for andOp_144.andOp_144_in1
	// Insensitive connections
	always @(*) begin
		andOp_144_in0 = valid ? bb_2_active_out_data : bb_2_active_out_data;
		andOp_144_in1 = valid ? eq_143_out : eq_143_out;
	end
	// controller for andOp_146.andOp_146_in0
	// controller for andOp_146.andOp_146_in1
	// Insensitive connections
	always @(*) begin
		andOp_146_in0 = valid ? bb_7_active_out_data : bb_7_active_out_data;
		andOp_146_in1 = valid ? eq_145_out : eq_145_out;
	end
	// controller for andOp_148.andOp_148_in0
	// controller for andOp_148.andOp_148_in1
	// Insensitive connections
	always @(*) begin
		andOp_148_in0 = valid ? bb_7_active_out_data : bb_7_active_out_data;
		andOp_148_in1 = valid ? eq_147_out : eq_147_out;
	end
	// controller for andOp_150.andOp_150_in0
	// controller for andOp_150.andOp_150_in1
	// Insensitive connections
	always @(*) begin
		andOp_150_in0 = valid ? bb_6_active_out_data : bb_6_active_out_data;
		andOp_150_in1 = valid ? eq_149_out : eq_149_out;
	end
	// controller for andOp_152.andOp_152_in0
	// controller for andOp_152.andOp_152_in1
	// Insensitive connections
	always @(*) begin
		andOp_152_in0 = valid ? bb_3_active_out_data : bb_3_active_out_data;
		andOp_152_in1 = valid ? eq_151_out : eq_151_out;
	end
	// controller for andOp_154.andOp_154_in0
	// controller for andOp_154.andOp_154_in1
	// Insensitive connections
	always @(*) begin
		andOp_154_in0 = valid ? bb_8_active_out_data : bb_8_active_out_data;
		andOp_154_in1 = valid ? eq_153_out : eq_153_out;
	end
	// controller for andOp_156.andOp_156_in0
	// controller for andOp_156.andOp_156_in1
	// Insensitive connections
	always @(*) begin
		andOp_156_in0 = valid ? notOp_155_out : notOp_155_out;
		andOp_156_in1 = valid ? andOp_152_out : andOp_152_out;
	end
	// controller for andOp_158.andOp_158_in0
	// controller for andOp_158.andOp_158_in1
	// Insensitive connections
	always @(*) begin
		andOp_158_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_158_in1 = valid ? eq_157_out : eq_157_out;
	end
	// controller for andOp_16.andOp_16_in0
	// controller for andOp_16.andOp_16_in1
	// Insensitive connections
	always @(*) begin
		andOp_16_in0 = valid ? andOp_14_out : andOp_14_out;
		andOp_16_in1 = valid ? icmp_tmp_5 : icmp_tmp_5;
	end
	// controller for andOp_160.andOp_160_in0
	// controller for andOp_160.andOp_160_in1
	// Insensitive connections
	always @(*) begin
		andOp_160_in0 = valid ? bb_3_active_out_data : bb_3_active_out_data;
		andOp_160_in1 = valid ? eq_159_out : eq_159_out;
	end
	// controller for andOp_162.andOp_162_in0
	// controller for andOp_162.andOp_162_in1
	// Insensitive connections
	always @(*) begin
		andOp_162_in0 = valid ? notOp_161_out : notOp_161_out;
		andOp_162_in1 = valid ? andOp_158_out : andOp_158_out;
	end
	// controller for andOp_164.andOp_164_in0
	// controller for andOp_164.andOp_164_in1
	// Insensitive connections
	always @(*) begin
		andOp_164_in0 = valid ? bb_9_active_out_data : bb_9_active_out_data;
		andOp_164_in1 = valid ? eq_163_out : eq_163_out;
	end
	// controller for andOp_166.andOp_166_in0
	// controller for andOp_166.andOp_166_in1
	// Insensitive connections
	always @(*) begin
		andOp_166_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_166_in1 = valid ? eq_165_out : eq_165_out;
	end
	// controller for andOp_168.andOp_168_in0
	// controller for andOp_168.andOp_168_in1
	// Insensitive connections
	always @(*) begin
		andOp_168_in0 = valid ? notOp_167_out : notOp_167_out;
		andOp_168_in1 = valid ? andOp_164_out : andOp_164_out;
	end
	// controller for andOp_170.andOp_170_in0
	// controller for andOp_170.andOp_170_in1
	// Insensitive connections
	always @(*) begin
		andOp_170_in0 = valid ? bb_8_active_out_data : bb_8_active_out_data;
		andOp_170_in1 = valid ? eq_169_out : eq_169_out;
	end
	// controller for andOp_172.andOp_172_in0
	// controller for andOp_172.andOp_172_in1
	// Insensitive connections
	always @(*) begin
		andOp_172_in0 = valid ? bb_9_active_out_data : bb_9_active_out_data;
		andOp_172_in1 = valid ? eq_171_out : eq_171_out;
	end
	// controller for andOp_174.andOp_174_in0
	// controller for andOp_174.andOp_174_in1
	// Insensitive connections
	always @(*) begin
		andOp_174_in0 = valid ? notOp_173_out : notOp_173_out;
		andOp_174_in1 = valid ? andOp_170_out : andOp_170_out;
	end
	// controller for andOp_176.andOp_176_in0
	// controller for andOp_176.andOp_176_in1
	// Insensitive connections
	always @(*) begin
		andOp_176_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_176_in1 = valid ? eq_175_out : eq_175_out;
	end
	// controller for andOp_178.andOp_178_in0
	// controller for andOp_178.andOp_178_in1
	// Insensitive connections
	always @(*) begin
		andOp_178_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_178_in1 = valid ? eq_177_out : eq_177_out;
	end
	// controller for andOp_18.andOp_18_in0
	// controller for andOp_18.andOp_18_in1
	// Insensitive connections
	always @(*) begin
		andOp_18_in0 = valid ? andOp_14_out : andOp_14_out;
		andOp_18_in1 = valid ? notOp_17_out : notOp_17_out;
	end
	// controller for andOp_180.andOp_180_in0
	// controller for andOp_180.andOp_180_in1
	// Insensitive connections
	always @(*) begin
		andOp_180_in0 = valid ? notOp_179_out : notOp_179_out;
		andOp_180_in1 = valid ? andOp_176_out : andOp_176_out;
	end
	// controller for andOp_182.andOp_182_in0
	// controller for andOp_182.andOp_182_in1
	// Insensitive connections
	always @(*) begin
		andOp_182_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_182_in1 = valid ? eq_181_out : eq_181_out;
	end
	// controller for andOp_184.andOp_184_in0
	// controller for andOp_184.andOp_184_in1
	// Insensitive connections
	always @(*) begin
		andOp_184_in0 = valid ? bb_1_active_out_data : bb_1_active_out_data;
		andOp_184_in1 = valid ? eq_183_out : eq_183_out;
	end
	// controller for andOp_186.andOp_186_in0
	// controller for andOp_186.andOp_186_in1
	// Insensitive connections
	always @(*) begin
		andOp_186_in0 = valid ? notOp_185_out : notOp_185_out;
		andOp_186_in1 = valid ? andOp_182_out : andOp_182_out;
	end
	// controller for andOp_188.andOp_188_in0
	// controller for andOp_188.andOp_188_in1
	// Insensitive connections
	always @(*) begin
		andOp_188_in0 = valid ? bb_3_active_out_data : bb_3_active_out_data;
		andOp_188_in1 = valid ? eq_187_out : eq_187_out;
	end
	// controller for andOp_190.andOp_190_in0
	// controller for andOp_190.andOp_190_in1
	// Insensitive connections
	always @(*) begin
		andOp_190_in0 = valid ? notOp_189_out : notOp_189_out;
		andOp_190_in1 = valid ? andOp_186_out : andOp_186_out;
	end
	// controller for andOp_192.andOp_192_in0
	// controller for andOp_192.andOp_192_in1
	// Insensitive connections
	always @(*) begin
		andOp_192_in0 = valid ? bb_1_active_out_data : bb_1_active_out_data;
		andOp_192_in1 = valid ? eq_191_out : eq_191_out;
	end
	// controller for andOp_194.andOp_194_in0
	// controller for andOp_194.andOp_194_in1
	// Insensitive connections
	always @(*) begin
		andOp_194_in0 = valid ? bb_5_active_out_data : bb_5_active_out_data;
		andOp_194_in1 = valid ? eq_193_out : eq_193_out;
	end
	// controller for andOp_196.andOp_196_in0
	// controller for andOp_196.andOp_196_in1
	// Insensitive connections
	always @(*) begin
		andOp_196_in0 = valid ? notOp_195_out : notOp_195_out;
		andOp_196_in1 = valid ? andOp_192_out : andOp_192_out;
	end
	// controller for andOp_198.andOp_198_in0
	// controller for andOp_198.andOp_198_in1
	// Insensitive connections
	always @(*) begin
		andOp_198_in0 = valid ? bb_2_active_out_data : bb_2_active_out_data;
		andOp_198_in1 = valid ? eq_197_out : eq_197_out;
	end
	// controller for andOp_2.andOp_2_in0
	// controller for andOp_2.andOp_2_in1
	// Insensitive connections
	always @(*) begin
		andOp_2_in0 = valid ? andOp_1_out : andOp_1_out;
		andOp_2_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_20.andOp_20_in0
	// controller for andOp_20.andOp_20_in1
	// Insensitive connections
	always @(*) begin
		andOp_20_in0 = valid ? bb_5_active_out_data : bb_5_active_out_data;
		andOp_20_in1 = valid ? eq_19_out : eq_19_out;
	end
	// controller for andOp_200.andOp_200_in0
	// controller for andOp_200.andOp_200_in1
	// Insensitive connections
	always @(*) begin
		andOp_200_in0 = valid ? bb_5_active_out_data : bb_5_active_out_data;
		andOp_200_in1 = valid ? eq_199_out : eq_199_out;
	end
	// controller for andOp_202.andOp_202_in0
	// controller for andOp_202.andOp_202_in1
	// Insensitive connections
	always @(*) begin
		andOp_202_in0 = valid ? bb_6_active_out_data : bb_6_active_out_data;
		andOp_202_in1 = valid ? eq_201_out : eq_201_out;
	end
	// controller for andOp_204.andOp_204_in0
	// controller for andOp_204.andOp_204_in1
	// Insensitive connections
	always @(*) begin
		andOp_204_in0 = valid ? notOp_203_out : notOp_203_out;
		andOp_204_in1 = valid ? andOp_200_out : andOp_200_out;
	end
	// controller for andOp_206.andOp_206_in0
	// controller for andOp_206.andOp_206_in1
	// Insensitive connections
	always @(*) begin
		andOp_206_in0 = valid ? bb_7_active_out_data : bb_7_active_out_data;
		andOp_206_in1 = valid ? eq_205_out : eq_205_out;
	end
	// controller for andOp_208.andOp_208_in0
	// controller for andOp_208.andOp_208_in1
	// Insensitive connections
	always @(*) begin
		andOp_208_in0 = valid ? bb_2_active_out_data : bb_2_active_out_data;
		andOp_208_in1 = valid ? eq_207_out : eq_207_out;
	end
	// controller for andOp_21.andOp_21_in0
	// controller for andOp_21.andOp_21_in1
	// Insensitive connections
	always @(*) begin
		andOp_21_in0 = valid ? andOp_20_out : andOp_20_out;
		andOp_21_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_210.andOp_210_in0
	// controller for andOp_210.andOp_210_in1
	// Insensitive connections
	always @(*) begin
		andOp_210_in0 = valid ? notOp_209_out : notOp_209_out;
		andOp_210_in1 = valid ? andOp_206_out : andOp_206_out;
	end
	// controller for andOp_212.andOp_212_in0
	// controller for andOp_212.andOp_212_in1
	// Insensitive connections
	always @(*) begin
		andOp_212_in0 = valid ? bb_6_active_out_data : bb_6_active_out_data;
		andOp_212_in1 = valid ? eq_211_out : eq_211_out;
	end
	// controller for andOp_214.andOp_214_in0
	// controller for andOp_214.andOp_214_in1
	// Insensitive connections
	always @(*) begin
		andOp_214_in0 = valid ? bb_7_active_out_data : bb_7_active_out_data;
		andOp_214_in1 = valid ? eq_213_out : eq_213_out;
	end
	// controller for andOp_216.andOp_216_in0
	// controller for andOp_216.andOp_216_in1
	// Insensitive connections
	always @(*) begin
		andOp_216_in0 = valid ? notOp_215_out : notOp_215_out;
		andOp_216_in1 = valid ? andOp_212_out : andOp_212_out;
	end
	// controller for andOp_218.andOp_218_in0
	// controller for andOp_218.andOp_218_in1
	// Insensitive connections
	always @(*) begin
		andOp_218_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_218_in1 = valid ? eq_217_out : eq_217_out;
	end
	// controller for andOp_219.andOp_219_in0
	// controller for andOp_219.andOp_219_in1
	// Insensitive connections
	always @(*) begin
		andOp_219_in0 = valid ? andOp_218_out : andOp_218_out;
		andOp_219_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_221.andOp_221_in0
	// controller for andOp_221.andOp_221_in1
	// Insensitive connections
	always @(*) begin
		andOp_221_in0 = valid ? eq_220_out : eq_220_out;
		andOp_221_in1 = valid ? andOp_219_out : andOp_219_out;
	end
	// controller for andOp_224.andOp_224_in0
	// controller for andOp_224.andOp_224_in1
	// Insensitive connections
	always @(*) begin
		andOp_224_in0 = valid ? bb_9_active_out_data : bb_9_active_out_data;
		andOp_224_in1 = valid ? eq_223_out : eq_223_out;
	end
	// controller for andOp_225.andOp_225_in0
	// controller for andOp_225.andOp_225_in1
	// Insensitive connections
	always @(*) begin
		andOp_225_in0 = valid ? andOp_224_out : andOp_224_out;
		andOp_225_in1 = valid ? notOp_222_out : notOp_222_out;
	end
	// controller for andOp_227.andOp_227_in0
	// controller for andOp_227.andOp_227_in1
	// Insensitive connections
	always @(*) begin
		andOp_227_in0 = valid ? eq_226_out : eq_226_out;
		andOp_227_in1 = valid ? andOp_225_out : andOp_225_out;
	end
	// controller for andOp_229.andOp_229_in0
	// controller for andOp_229.andOp_229_in1
	// Insensitive connections
	always @(*) begin
		andOp_229_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_229_in1 = valid ? eq_228_out : eq_228_out;
	end
	// controller for andOp_230.andOp_230_in0
	// controller for andOp_230.andOp_230_in1
	// Insensitive connections
	always @(*) begin
		andOp_230_in0 = valid ? andOp_229_out : andOp_229_out;
		andOp_230_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_232.andOp_232_in0
	// controller for andOp_232.andOp_232_in1
	// Insensitive connections
	always @(*) begin
		andOp_232_in0 = valid ? eq_231_out : eq_231_out;
		andOp_232_in1 = valid ? andOp_230_out : andOp_230_out;
	end
	// controller for andOp_234.andOp_234_in0
	// controller for andOp_234.andOp_234_in1
	// Insensitive connections
	always @(*) begin
		andOp_234_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_234_in1 = valid ? eq_233_out : eq_233_out;
	end
	// controller for andOp_235.andOp_235_in0
	// controller for andOp_235.andOp_235_in1
	// Insensitive connections
	always @(*) begin
		andOp_235_in0 = valid ? andOp_234_out : andOp_234_out;
		andOp_235_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_237.andOp_237_in0
	// controller for andOp_237.andOp_237_in1
	// Insensitive connections
	always @(*) begin
		andOp_237_in0 = valid ? eq_236_out : eq_236_out;
		andOp_237_in1 = valid ? andOp_235_out : andOp_235_out;
	end
	// controller for andOp_239.andOp_239_in0
	// controller for andOp_239.andOp_239_in1
	// Insensitive connections
	always @(*) begin
		andOp_239_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_239_in1 = valid ? eq_238_out : eq_238_out;
	end
	// controller for andOp_24.andOp_24_in0
	// controller for andOp_24.andOp_24_in1
	// Insensitive connections
	always @(*) begin
		andOp_24_in0 = valid ? bb_6_active_out_data : bb_6_active_out_data;
		andOp_24_in1 = valid ? eq_23_out : eq_23_out;
	end
	// controller for andOp_240.andOp_240_in0
	// controller for andOp_240.andOp_240_in1
	// Insensitive connections
	always @(*) begin
		andOp_240_in0 = valid ? andOp_239_out : andOp_239_out;
		andOp_240_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_242.andOp_242_in0
	// controller for andOp_242.andOp_242_in1
	// Insensitive connections
	always @(*) begin
		andOp_242_in0 = valid ? eq_241_out : eq_241_out;
		andOp_242_in1 = valid ? andOp_240_out : andOp_240_out;
	end
	// controller for andOp_245.andOp_245_in0
	// controller for andOp_245.andOp_245_in1
	// Insensitive connections
	always @(*) begin
		andOp_245_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_245_in1 = valid ? eq_244_out : eq_244_out;
	end
	// controller for andOp_246.andOp_246_in0
	// controller for andOp_246.andOp_246_in1
	// Insensitive connections
	always @(*) begin
		andOp_246_in0 = valid ? andOp_245_out : andOp_245_out;
		andOp_246_in1 = valid ? notOp_243_out : notOp_243_out;
	end
	// controller for andOp_248.andOp_248_in0
	// controller for andOp_248.andOp_248_in1
	// Insensitive connections
	always @(*) begin
		andOp_248_in0 = valid ? eq_247_out : eq_247_out;
		andOp_248_in1 = valid ? andOp_246_out : andOp_246_out;
	end
	// controller for andOp_25.andOp_25_in0
	// controller for andOp_25.andOp_25_in1
	// Insensitive connections
	always @(*) begin
		andOp_25_in0 = valid ? andOp_24_out : andOp_24_out;
		andOp_25_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_251.andOp_251_in0
	// controller for andOp_251.andOp_251_in1
	// Insensitive connections
	always @(*) begin
		andOp_251_in0 = valid ? bb_6_active_out_data : bb_6_active_out_data;
		andOp_251_in1 = valid ? eq_250_out : eq_250_out;
	end
	// controller for andOp_252.andOp_252_in0
	// controller for andOp_252.andOp_252_in1
	// Insensitive connections
	always @(*) begin
		andOp_252_in0 = valid ? andOp_251_out : andOp_251_out;
		andOp_252_in1 = valid ? notOp_249_out : notOp_249_out;
	end
	// controller for andOp_254.andOp_254_in0
	// controller for andOp_254.andOp_254_in1
	// Insensitive connections
	always @(*) begin
		andOp_254_in0 = valid ? eq_253_out : eq_253_out;
		andOp_254_in1 = valid ? andOp_252_out : andOp_252_out;
	end
	// controller for andOp_256.andOp_256_in0
	// controller for andOp_256.andOp_256_in1
	// Insensitive connections
	always @(*) begin
		andOp_256_in0 = valid ? bb_2_active_out_data : bb_2_active_out_data;
		andOp_256_in1 = valid ? eq_255_out : eq_255_out;
	end
	// controller for andOp_257.andOp_257_in0
	// controller for andOp_257.andOp_257_in1
	// Insensitive connections
	always @(*) begin
		andOp_257_in0 = valid ? andOp_256_out : andOp_256_out;
		andOp_257_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_259.andOp_259_in0
	// controller for andOp_259.andOp_259_in1
	// Insensitive connections
	always @(*) begin
		andOp_259_in0 = valid ? eq_258_out : eq_258_out;
		andOp_259_in1 = valid ? andOp_257_out : andOp_257_out;
	end
	// controller for andOp_261.andOp_261_in0
	// controller for andOp_261.andOp_261_in1
	// Insensitive connections
	always @(*) begin
		andOp_261_in0 = valid ? bb_3_active_out_data : bb_3_active_out_data;
		andOp_261_in1 = valid ? eq_260_out : eq_260_out;
	end
	// controller for andOp_263.andOp_263_in0
	// controller for andOp_263.andOp_263_in1
	// Insensitive connections
	always @(*) begin
		andOp_263_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_263_in1 = valid ? eq_262_out : eq_262_out;
	end
	// controller for andOp_265.andOp_265_in0
	// controller for andOp_265.andOp_265_in1
	// Insensitive connections
	always @(*) begin
		andOp_265_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_265_in1 = valid ? eq_264_out : eq_264_out;
	end
	// controller for andOp_267.andOp_267_in0
	// controller for andOp_267.andOp_267_in1
	// Insensitive connections
	always @(*) begin
		andOp_267_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_267_in1 = valid ? eq_266_out : eq_266_out;
	end
	// controller for andOp_27.andOp_27_in0
	// controller for andOp_27.andOp_27_in1
	// Insensitive connections
	always @(*) begin
		andOp_27_in0 = valid ? andOp_25_out : andOp_25_out;
		andOp_27_in1 = valid ? out_write_ready : out_write_ready;
	end
	// controller for andOp_29.andOp_29_in0
	// controller for andOp_29.andOp_29_in1
	// Insensitive connections
	always @(*) begin
		andOp_29_in0 = valid ? andOp_25_out : andOp_25_out;
		andOp_29_in1 = valid ? notOp_28_out : notOp_28_out;
	end
	// controller for andOp_31.andOp_31_in0
	// controller for andOp_31.andOp_31_in1
	// Insensitive connections
	always @(*) begin
		andOp_31_in0 = valid ? bb_7_active_out_data : bb_7_active_out_data;
		andOp_31_in1 = valid ? eq_30_out : eq_30_out;
	end
	// controller for andOp_32.andOp_32_in0
	// controller for andOp_32.andOp_32_in1
	// Insensitive connections
	always @(*) begin
		andOp_32_in0 = valid ? andOp_31_out : andOp_31_out;
		andOp_32_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_35.andOp_35_in0
	// controller for andOp_35.andOp_35_in1
	// Insensitive connections
	always @(*) begin
		andOp_35_in0 = valid ? bb_8_active_out_data : bb_8_active_out_data;
		andOp_35_in1 = valid ? eq_34_out : eq_34_out;
	end
	// controller for andOp_36.andOp_36_in0
	// controller for andOp_36.andOp_36_in1
	// Insensitive connections
	always @(*) begin
		andOp_36_in0 = valid ? andOp_35_out : andOp_35_out;
		andOp_36_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_39.andOp_39_in0
	// controller for andOp_39.andOp_39_in1
	// Insensitive connections
	always @(*) begin
		andOp_39_in0 = valid ? bb_9_active_out_data : bb_9_active_out_data;
		andOp_39_in1 = valid ? eq_38_out : eq_38_out;
	end
	// controller for andOp_40.andOp_40_in0
	// controller for andOp_40.andOp_40_in1
	// Insensitive connections
	always @(*) begin
		andOp_40_in0 = valid ? andOp_39_out : andOp_39_out;
		andOp_40_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_42.andOp_42_in0
	// controller for andOp_42.andOp_42_in1
	// Insensitive connections
	always @(*) begin
		andOp_42_in0 = valid ? andOp_40_out : andOp_40_out;
		andOp_42_in1 = valid ? in_read_ready : in_read_ready;
	end
	// controller for andOp_44.andOp_44_in0
	// controller for andOp_44.andOp_44_in1
	// Insensitive connections
	always @(*) begin
		andOp_44_in0 = valid ? andOp_40_out : andOp_40_out;
		andOp_44_in1 = valid ? notOp_43_out : notOp_43_out;
	end
	// controller for andOp_46.andOp_46_in0
	// controller for andOp_46.andOp_46_in1
	// Insensitive connections
	always @(*) begin
		andOp_46_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_46_in1 = valid ? eq_45_out : eq_45_out;
	end
	// controller for andOp_47.andOp_47_in0
	// controller for andOp_47.andOp_47_in1
	// Insensitive connections
	always @(*) begin
		andOp_47_in0 = valid ? andOp_46_out : andOp_46_out;
		andOp_47_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_5.andOp_5_in0
	// controller for andOp_5.andOp_5_in1
	// Insensitive connections
	always @(*) begin
		andOp_5_in0 = valid ? bb_1_active_out_data : bb_1_active_out_data;
		andOp_5_in1 = valid ? eq_4_out : eq_4_out;
	end
	// controller for andOp_6.andOp_6_in0
	// controller for andOp_6.andOp_6_in1
	// Insensitive connections
	always @(*) begin
		andOp_6_in0 = valid ? andOp_5_out : andOp_5_out;
		andOp_6_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_71.andOp_71_in0
	// controller for andOp_71.andOp_71_in1
	// Insensitive connections
	always @(*) begin
		andOp_71_in0 = valid ? bb_0_active_out_data : bb_0_active_out_data;
		andOp_71_in1 = valid ? eq_70_out : eq_70_out;
	end
	// controller for andOp_73.andOp_73_in0
	// controller for andOp_73.andOp_73_in1
	// Insensitive connections
	always @(*) begin
		andOp_73_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_73_in1 = valid ? eq_72_out : eq_72_out;
	end
	// controller for andOp_75.andOp_75_in0
	// controller for andOp_75.andOp_75_in1
	// Insensitive connections
	always @(*) begin
		andOp_75_in0 = valid ? bb_10_active_out_data : bb_10_active_out_data;
		andOp_75_in1 = valid ? eq_74_out : eq_74_out;
	end
	// controller for andOp_77.andOp_77_in0
	// controller for andOp_77.andOp_77_in1
	// Insensitive connections
	always @(*) begin
		andOp_77_in0 = valid ? bb_4_active_out_data : bb_4_active_out_data;
		andOp_77_in1 = valid ? eq_76_out : eq_76_out;
	end
	// controller for andOp_79.andOp_79_in0
	// controller for andOp_79.andOp_79_in1
	// Insensitive connections
	always @(*) begin
		andOp_79_in0 = valid ? bb_2_active_out_data : bb_2_active_out_data;
		andOp_79_in1 = valid ? eq_78_out : eq_78_out;
	end
	// controller for andOp_83.andOp_83_in0
	// controller for andOp_83.andOp_83_in1
	// Insensitive connections
	always @(*) begin
		andOp_83_in0 = valid ? notOp_82_out : notOp_82_out;
		andOp_83_in1 = valid ? andOp_16_out : andOp_16_out;
	end
	// controller for andOp_86.andOp_86_in0
	// controller for andOp_86.andOp_86_in1
	// Insensitive connections
	always @(*) begin
		andOp_86_in0 = valid ? notOp_85_out : notOp_85_out;
		andOp_86_in1 = valid ? andOp_32_out : andOp_32_out;
	end
	// controller for andOp_89.andOp_89_in0
	// controller for andOp_89.andOp_89_in1
	// Insensitive connections
	always @(*) begin
		andOp_89_in0 = valid ? notOp_88_out : notOp_88_out;
		andOp_89_in1 = valid ? andOp_2_out : andOp_2_out;
	end
	// controller for andOp_9.andOp_9_in0
	// controller for andOp_9.andOp_9_in1
	// Insensitive connections
	always @(*) begin
		andOp_9_in0 = valid ? bb_3_active_out_data : bb_3_active_out_data;
		andOp_9_in1 = valid ? eq_8_out : eq_8_out;
	end
	// controller for andOp_92.andOp_92_in0
	// controller for andOp_92.andOp_92_in1
	// Insensitive connections
	always @(*) begin
		andOp_92_in0 = valid ? notOp_91_out : notOp_91_out;
		andOp_92_in1 = valid ? andOp_47_out : andOp_47_out;
	end
	// controller for andOp_95.andOp_95_in0
	// controller for andOp_95.andOp_95_in1
	// Insensitive connections
	always @(*) begin
		andOp_95_in0 = valid ? notOp_94_out : notOp_94_out;
		andOp_95_in1 = valid ? andOp_6_out : andOp_6_out;
	end
	// controller for andOp_98.andOp_98_in0
	// controller for andOp_98.andOp_98_in1
	// Insensitive connections
	always @(*) begin
		andOp_98_in0 = valid ? notOp_97_out : notOp_97_out;
		andOp_98_in1 = valid ? andOp_21_out : andOp_21_out;
	end
	// controller for bb_0_active.bb_0_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_data = eq_49_out;
		end else begin
			bb_0_active_in_data = 0;
		end
	end
	// controller for bb_0_predecessor.bb_0_predecessor_in_data
	always @(*) begin
		if (eq_80_out) begin 
			bb_0_predecessor_in_data = last_BB_reg;
		end else begin
			bb_0_predecessor_in_data = 0;
		end
	end
	// controller for bb_10_active.bb_10_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_data = orOp_69_out;
		end else begin
			bb_10_active_in_data = 0;
		end
	end
	// controller for bb_10_predecessor.bb_10_predecessor_in_data
	always @(*) begin
		if (andOp_110_out) begin 
			bb_10_predecessor_in_data = 32'd9;
		end else if (eq_108_out) begin 
			bb_10_predecessor_in_data = last_BB_reg;
		end else begin
			bb_10_predecessor_in_data = 0;
		end
	end
	// controller for bb_1_active.bb_1_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_data = orOp_51_out;
		end else begin
			bb_1_active_in_data = 0;
		end
	end
	// controller for bb_1_predecessor.bb_1_predecessor_in_data
	always @(*) begin
		if (andOp_83_out) begin 
			bb_1_predecessor_in_data = 32'd4;
		end else if (eq_81_out) begin 
			bb_1_predecessor_in_data = last_BB_reg;
		end else begin
			bb_1_predecessor_in_data = 0;
		end
	end
	// controller for bb_2_active.bb_2_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_data = orOp_53_out;
		end else begin
			bb_2_active_in_data = 0;
		end
	end
	// controller for bb_2_predecessor.bb_2_predecessor_in_data
	always @(*) begin
		if (andOp_86_out) begin 
			bb_2_predecessor_in_data = 32'd7;
		end else if (eq_84_out) begin 
			bb_2_predecessor_in_data = last_BB_reg;
		end else begin
			bb_2_predecessor_in_data = 0;
		end
	end
	// controller for bb_3_active.bb_3_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_data = orOp_55_out;
		end else begin
			bb_3_active_in_data = 0;
		end
	end
	// controller for bb_3_predecessor.bb_3_predecessor_in_data
	always @(*) begin
		if (andOp_89_out) begin 
			bb_3_predecessor_in_data = 32'd0;
		end else if (eq_87_out) begin 
			bb_3_predecessor_in_data = last_BB_reg;
		end else begin
			bb_3_predecessor_in_data = 0;
		end
	end
	// controller for bb_4_active.bb_4_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_data = orOp_57_out;
		end else begin
			bb_4_active_in_data = 0;
		end
	end
	// controller for bb_4_predecessor.bb_4_predecessor_in_data
	always @(*) begin
		if (andOp_92_out) begin 
			bb_4_predecessor_in_data = 32'd10;
		end else if (eq_90_out) begin 
			bb_4_predecessor_in_data = last_BB_reg;
		end else begin
			bb_4_predecessor_in_data = 0;
		end
	end
	// controller for bb_5_active.bb_5_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_5_active_in_data = orOp_59_out;
		end else begin
			bb_5_active_in_data = 0;
		end
	end
	// controller for bb_5_predecessor.bb_5_predecessor_in_data
	always @(*) begin
		if (andOp_95_out) begin 
			bb_5_predecessor_in_data = 32'd1;
		end else if (eq_93_out) begin 
			bb_5_predecessor_in_data = last_BB_reg;
		end else begin
			bb_5_predecessor_in_data = 0;
		end
	end
	// controller for bb_6_active.bb_6_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_6_active_in_data = orOp_61_out;
		end else begin
			bb_6_active_in_data = 0;
		end
	end
	// controller for bb_6_predecessor.bb_6_predecessor_in_data
	always @(*) begin
		if (andOp_98_out) begin 
			bb_6_predecessor_in_data = 32'd5;
		end else if (eq_96_out) begin 
			bb_6_predecessor_in_data = last_BB_reg;
		end else begin
			bb_6_predecessor_in_data = 0;
		end
	end
	// controller for bb_7_active.bb_7_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_7_active_in_data = orOp_63_out;
		end else begin
			bb_7_active_in_data = 0;
		end
	end
	// controller for bb_7_predecessor.bb_7_predecessor_in_data
	always @(*) begin
		if (andOp_101_out) begin 
			bb_7_predecessor_in_data = 32'd6;
		end else if (eq_99_out) begin 
			bb_7_predecessor_in_data = last_BB_reg;
		end else begin
			bb_7_predecessor_in_data = 0;
		end
	end
	// controller for bb_8_active.bb_8_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_data = orOp_65_out;
		end else begin
			bb_8_active_in_data = 0;
		end
	end
	// controller for bb_8_predecessor.bb_8_predecessor_in_data
	always @(*) begin
		if (andOp_104_out) begin 
			bb_8_predecessor_in_data = 32'd3;
		end else if (eq_102_out) begin 
			bb_8_predecessor_in_data = last_BB_reg;
		end else begin
			bb_8_predecessor_in_data = 0;
		end
	end
	// controller for bb_9_active.bb_9_active_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_9_active_in_data = orOp_67_out;
		end else begin
			bb_9_active_in_data = 0;
		end
	end
	// controller for bb_9_predecessor.bb_9_predecessor_in_data
	always @(*) begin
		if (andOp_107_out) begin 
			bb_9_predecessor_in_data = 32'd8;
		end else if (eq_105_out) begin 
			bb_9_predecessor_in_data = last_BB_reg;
		end else begin
			bb_9_predecessor_in_data = 0;
		end
	end
	// controller for br_0_happened.br_0_happened_in_data
	always @(*) begin
		if (andOp_2_out) begin 
			br_0_happened_in_data = 1'd1;
		end else if (notOp_3_out) begin 
			br_0_happened_in_data = 1'd0;
		end else begin
			br_0_happened_in_data = 0;
		end
	end
	// controller for br_10_happened.br_10_happened_in_data
	always @(*) begin
		if (andOp_47_out) begin 
			br_10_happened_in_data = 1'd1;
		end else if (notOp_48_out) begin 
			br_10_happened_in_data = 1'd0;
		end else begin
			br_10_happened_in_data = 0;
		end
	end
	// controller for br_1_happened.br_1_happened_in_data
	always @(*) begin
		if (andOp_6_out) begin 
			br_1_happened_in_data = 1'd1;
		end else if (notOp_7_out) begin 
			br_1_happened_in_data = 1'd0;
		end else begin
			br_1_happened_in_data = 0;
		end
	end
	// controller for br_3_happened.br_3_happened_in_data
	always @(*) begin
		if (andOp_10_out) begin 
			br_3_happened_in_data = 1'd1;
		end else if (notOp_11_out) begin 
			br_3_happened_in_data = 1'd0;
		end else begin
			br_3_happened_in_data = 0;
		end
	end
	// controller for br_4_happened.br_4_happened_in_data
	always @(*) begin
		if (andOp_14_out) begin 
			br_4_happened_in_data = 1'd1;
		end else if (notOp_15_out) begin 
			br_4_happened_in_data = 1'd0;
		end else begin
			br_4_happened_in_data = 0;
		end
	end
	// controller for br_5_happened.br_5_happened_in_data
	always @(*) begin
		if (andOp_21_out) begin 
			br_5_happened_in_data = 1'd1;
		end else if (notOp_22_out) begin 
			br_5_happened_in_data = 1'd0;
		end else begin
			br_5_happened_in_data = 0;
		end
	end
	// controller for br_6_happened.br_6_happened_in_data
	always @(*) begin
		if (andOp_25_out) begin 
			br_6_happened_in_data = 1'd1;
		end else if (notOp_26_out) begin 
			br_6_happened_in_data = 1'd0;
		end else begin
			br_6_happened_in_data = 0;
		end
	end
	// controller for br_7_happened.br_7_happened_in_data
	always @(*) begin
		if (andOp_32_out) begin 
			br_7_happened_in_data = 1'd1;
		end else if (notOp_33_out) begin 
			br_7_happened_in_data = 1'd0;
		end else begin
			br_7_happened_in_data = 0;
		end
	end
	// controller for br_8_happened.br_8_happened_in_data
	always @(*) begin
		if (andOp_36_out) begin 
			br_8_happened_in_data = 1'd1;
		end else if (notOp_37_out) begin 
			br_8_happened_in_data = 1'd0;
		end else begin
			br_8_happened_in_data = 0;
		end
	end
	// controller for br_9_happened.br_9_happened_in_data
	always @(*) begin
		if (andOp_40_out) begin 
			br_9_happened_in_data = 1'd1;
		end else if (notOp_41_out) begin 
			br_9_happened_in_data = 1'd0;
		end else begin
			br_9_happened_in_data = 0;
		end
	end
	// controller for eq_0.eq_0_in0
	// controller for eq_0.eq_0_in1
	// Insensitive connections
	always @(*) begin
		eq_0_in0 = valid ? 32'd1 : 32'd1;
		eq_0_in1 = valid ? global_state : global_state;
	end
	// controller for eq_102.eq_102_in0
	// controller for eq_102.eq_102_in1
	// Insensitive connections
	always @(*) begin
		eq_102_in0 = valid ? 32'd8 : 32'd8;
		eq_102_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_105.eq_105_in0
	// controller for eq_105.eq_105_in1
	// Insensitive connections
	always @(*) begin
		eq_105_in0 = valid ? 32'd9 : 32'd9;
		eq_105_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_108.eq_108_in0
	// controller for eq_108.eq_108_in1
	// Insensitive connections
	always @(*) begin
		eq_108_in0 = valid ? 32'd10 : 32'd10;
		eq_108_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_111.eq_111_in0
	// controller for eq_111.eq_111_in1
	// Insensitive connections
	always @(*) begin
		eq_111_in0 = valid ? 32'd0 : 32'd0;
		eq_111_in1 = valid ? global_state : global_state;
	end
	// controller for eq_113.eq_113_in0
	// controller for eq_113.eq_113_in1
	// Insensitive connections
	always @(*) begin
		eq_113_in0 = valid ? 32'd3 : 32'd3;
		eq_113_in1 = valid ? global_state : global_state;
	end
	// controller for eq_115.eq_115_in0
	// controller for eq_115.eq_115_in1
	// Insensitive connections
	always @(*) begin
		eq_115_in0 = valid ? 32'd3 : 32'd3;
		eq_115_in1 = valid ? global_state : global_state;
	end
	// controller for eq_117.eq_117_in0
	// controller for eq_117.eq_117_in1
	// Insensitive connections
	always @(*) begin
		eq_117_in0 = valid ? 32'd4 : 32'd4;
		eq_117_in1 = valid ? global_state : global_state;
	end
	// controller for eq_119.eq_119_in0
	// controller for eq_119.eq_119_in1
	// Insensitive connections
	always @(*) begin
		eq_119_in0 = valid ? 32'd0 : 32'd0;
		eq_119_in1 = valid ? global_state : global_state;
	end
	// controller for eq_12.eq_12_in0
	// controller for eq_12.eq_12_in1
	// Insensitive connections
	always @(*) begin
		eq_12_in0 = valid ? 32'd4 : 32'd4;
		eq_12_in1 = valid ? global_state : global_state;
	end
	// controller for eq_121.eq_121_in0
	// controller for eq_121.eq_121_in1
	// Insensitive connections
	always @(*) begin
		eq_121_in0 = valid ? 32'd0 : 32'd0;
		eq_121_in1 = valid ? global_state : global_state;
	end
	// controller for eq_123.eq_123_in0
	// controller for eq_123.eq_123_in1
	// Insensitive connections
	always @(*) begin
		eq_123_in0 = valid ? 32'd0 : 32'd0;
		eq_123_in1 = valid ? global_state : global_state;
	end
	// controller for eq_125.eq_125_in0
	// controller for eq_125.eq_125_in1
	// Insensitive connections
	always @(*) begin
		eq_125_in0 = valid ? 32'd1 : 32'd1;
		eq_125_in1 = valid ? global_state : global_state;
	end
	// controller for eq_127.eq_127_in0
	// controller for eq_127.eq_127_in1
	// Insensitive connections
	always @(*) begin
		eq_127_in0 = valid ? 32'd1 : 32'd1;
		eq_127_in1 = valid ? global_state : global_state;
	end
	// controller for eq_129.eq_129_in0
	// controller for eq_129.eq_129_in1
	// Insensitive connections
	always @(*) begin
		eq_129_in0 = valid ? 32'd2 : 32'd2;
		eq_129_in1 = valid ? global_state : global_state;
	end
	// controller for eq_131.eq_131_in0
	// controller for eq_131.eq_131_in1
	// Insensitive connections
	always @(*) begin
		eq_131_in0 = valid ? 32'd3 : 32'd3;
		eq_131_in1 = valid ? global_state : global_state;
	end
	// controller for eq_133.eq_133_in0
	// controller for eq_133.eq_133_in1
	// Insensitive connections
	always @(*) begin
		eq_133_in0 = valid ? 32'd3 : 32'd3;
		eq_133_in1 = valid ? global_state : global_state;
	end
	// controller for eq_136.eq_136_in0
	// controller for eq_136.eq_136_in1
	// Insensitive connections
	always @(*) begin
		eq_136_in0 = valid ? 32'd10 : 32'd10;
		eq_136_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_137.eq_137_in0
	// controller for eq_137.eq_137_in1
	// Insensitive connections
	always @(*) begin
		eq_137_in0 = valid ? 32'd3 : 32'd3;
		eq_137_in1 = valid ? global_state : global_state;
	end
	// controller for eq_139.eq_139_in0
	// controller for eq_139.eq_139_in1
	// Insensitive connections
	always @(*) begin
		eq_139_in0 = valid ? 32'd3 : 32'd3;
		eq_139_in1 = valid ? global_state : global_state;
	end
	// controller for eq_141.eq_141_in0
	// controller for eq_141.eq_141_in1
	// Insensitive connections
	always @(*) begin
		eq_141_in0 = valid ? 32'd4 : 32'd4;
		eq_141_in1 = valid ? global_state : global_state;
	end
	// controller for eq_143.eq_143_in0
	// controller for eq_143.eq_143_in1
	// Insensitive connections
	always @(*) begin
		eq_143_in0 = valid ? 32'd4 : 32'd4;
		eq_143_in1 = valid ? global_state : global_state;
	end
	// controller for eq_145.eq_145_in0
	// controller for eq_145.eq_145_in1
	// Insensitive connections
	always @(*) begin
		eq_145_in0 = valid ? 32'd4 : 32'd4;
		eq_145_in1 = valid ? global_state : global_state;
	end
	// controller for eq_147.eq_147_in0
	// controller for eq_147.eq_147_in1
	// Insensitive connections
	always @(*) begin
		eq_147_in0 = valid ? 32'd4 : 32'd4;
		eq_147_in1 = valid ? global_state : global_state;
	end
	// controller for eq_149.eq_149_in0
	// controller for eq_149.eq_149_in1
	// Insensitive connections
	always @(*) begin
		eq_149_in0 = valid ? 32'd4 : 32'd4;
		eq_149_in1 = valid ? global_state : global_state;
	end
	// controller for eq_151.eq_151_in0
	// controller for eq_151.eq_151_in1
	// Insensitive connections
	always @(*) begin
		eq_151_in0 = valid ? 32'd1 : 32'd1;
		eq_151_in1 = valid ? global_state : global_state;
	end
	// controller for eq_153.eq_153_in0
	// controller for eq_153.eq_153_in1
	// Insensitive connections
	always @(*) begin
		eq_153_in0 = valid ? 32'd1 : 32'd1;
		eq_153_in1 = valid ? global_state : global_state;
	end
	// controller for eq_157.eq_157_in0
	// controller for eq_157.eq_157_in1
	// Insensitive connections
	always @(*) begin
		eq_157_in0 = valid ? 32'd1 : 32'd1;
		eq_157_in1 = valid ? global_state : global_state;
	end
	// controller for eq_159.eq_159_in0
	// controller for eq_159.eq_159_in1
	// Insensitive connections
	always @(*) begin
		eq_159_in0 = valid ? 32'd1 : 32'd1;
		eq_159_in1 = valid ? global_state : global_state;
	end
	// controller for eq_163.eq_163_in0
	// controller for eq_163.eq_163_in1
	// Insensitive connections
	always @(*) begin
		eq_163_in0 = valid ? 32'd1 : 32'd1;
		eq_163_in1 = valid ? global_state : global_state;
	end
	// controller for eq_165.eq_165_in0
	// controller for eq_165.eq_165_in1
	// Insensitive connections
	always @(*) begin
		eq_165_in0 = valid ? 32'd1 : 32'd1;
		eq_165_in1 = valid ? global_state : global_state;
	end
	// controller for eq_169.eq_169_in0
	// controller for eq_169.eq_169_in1
	// Insensitive connections
	always @(*) begin
		eq_169_in0 = valid ? 32'd1 : 32'd1;
		eq_169_in1 = valid ? global_state : global_state;
	end
	// controller for eq_171.eq_171_in0
	// controller for eq_171.eq_171_in1
	// Insensitive connections
	always @(*) begin
		eq_171_in0 = valid ? 32'd1 : 32'd1;
		eq_171_in1 = valid ? global_state : global_state;
	end
	// controller for eq_175.eq_175_in0
	// controller for eq_175.eq_175_in1
	// Insensitive connections
	always @(*) begin
		eq_175_in0 = valid ? 32'd3 : 32'd3;
		eq_175_in1 = valid ? global_state : global_state;
	end
	// controller for eq_177.eq_177_in0
	// controller for eq_177.eq_177_in1
	// Insensitive connections
	always @(*) begin
		eq_177_in0 = valid ? 32'd3 : 32'd3;
		eq_177_in1 = valid ? global_state : global_state;
	end
	// controller for eq_181.eq_181_in0
	// controller for eq_181.eq_181_in1
	// Insensitive connections
	always @(*) begin
		eq_181_in0 = valid ? 32'd4 : 32'd4;
		eq_181_in1 = valid ? global_state : global_state;
	end
	// controller for eq_183.eq_183_in0
	// controller for eq_183.eq_183_in1
	// Insensitive connections
	always @(*) begin
		eq_183_in0 = valid ? 32'd4 : 32'd4;
		eq_183_in1 = valid ? global_state : global_state;
	end
	// controller for eq_187.eq_187_in0
	// controller for eq_187.eq_187_in1
	// Insensitive connections
	always @(*) begin
		eq_187_in0 = valid ? 32'd4 : 32'd4;
		eq_187_in1 = valid ? global_state : global_state;
	end
	// controller for eq_19.eq_19_in0
	// controller for eq_19.eq_19_in1
	// Insensitive connections
	always @(*) begin
		eq_19_in0 = valid ? 32'd4 : 32'd4;
		eq_19_in1 = valid ? global_state : global_state;
	end
	// controller for eq_191.eq_191_in0
	// controller for eq_191.eq_191_in1
	// Insensitive connections
	always @(*) begin
		eq_191_in0 = valid ? 32'd4 : 32'd4;
		eq_191_in1 = valid ? global_state : global_state;
	end
	// controller for eq_193.eq_193_in0
	// controller for eq_193.eq_193_in1
	// Insensitive connections
	always @(*) begin
		eq_193_in0 = valid ? 32'd4 : 32'd4;
		eq_193_in1 = valid ? global_state : global_state;
	end
	// controller for eq_197.eq_197_in0
	// controller for eq_197.eq_197_in1
	// Insensitive connections
	always @(*) begin
		eq_197_in0 = valid ? 32'd4 : 32'd4;
		eq_197_in1 = valid ? global_state : global_state;
	end
	// controller for eq_199.eq_199_in0
	// controller for eq_199.eq_199_in1
	// Insensitive connections
	always @(*) begin
		eq_199_in0 = valid ? 32'd4 : 32'd4;
		eq_199_in1 = valid ? global_state : global_state;
	end
	// controller for eq_201.eq_201_in0
	// controller for eq_201.eq_201_in1
	// Insensitive connections
	always @(*) begin
		eq_201_in0 = valid ? 32'd4 : 32'd4;
		eq_201_in1 = valid ? global_state : global_state;
	end
	// controller for eq_205.eq_205_in0
	// controller for eq_205.eq_205_in1
	// Insensitive connections
	always @(*) begin
		eq_205_in0 = valid ? 32'd4 : 32'd4;
		eq_205_in1 = valid ? global_state : global_state;
	end
	// controller for eq_207.eq_207_in0
	// controller for eq_207.eq_207_in1
	// Insensitive connections
	always @(*) begin
		eq_207_in0 = valid ? 32'd4 : 32'd4;
		eq_207_in1 = valid ? global_state : global_state;
	end
	// controller for eq_211.eq_211_in0
	// controller for eq_211.eq_211_in1
	// Insensitive connections
	always @(*) begin
		eq_211_in0 = valid ? 32'd4 : 32'd4;
		eq_211_in1 = valid ? global_state : global_state;
	end
	// controller for eq_213.eq_213_in0
	// controller for eq_213.eq_213_in1
	// Insensitive connections
	always @(*) begin
		eq_213_in0 = valid ? 32'd4 : 32'd4;
		eq_213_in1 = valid ? global_state : global_state;
	end
	// controller for eq_217.eq_217_in0
	// controller for eq_217.eq_217_in1
	// Insensitive connections
	always @(*) begin
		eq_217_in0 = valid ? 32'd0 : 32'd0;
		eq_217_in1 = valid ? global_state : global_state;
	end
	// controller for eq_220.eq_220_in0
	// controller for eq_220.eq_220_in1
	// Insensitive connections
	always @(*) begin
		eq_220_in0 = valid ? 32'd0 : 32'd0;
		eq_220_in1 = valid ? global_state : global_state;
	end
	// controller for eq_223.eq_223_in0
	// controller for eq_223.eq_223_in1
	// Insensitive connections
	always @(*) begin
		eq_223_in0 = valid ? 32'd1 : 32'd1;
		eq_223_in1 = valid ? global_state : global_state;
	end
	// controller for eq_226.eq_226_in0
	// controller for eq_226.eq_226_in1
	// Insensitive connections
	always @(*) begin
		eq_226_in0 = valid ? 32'd1 : 32'd1;
		eq_226_in1 = valid ? global_state : global_state;
	end
	// controller for eq_228.eq_228_in0
	// controller for eq_228.eq_228_in1
	// Insensitive connections
	always @(*) begin
		eq_228_in0 = valid ? 32'd1 : 32'd1;
		eq_228_in1 = valid ? global_state : global_state;
	end
	// controller for eq_23.eq_23_in0
	// controller for eq_23.eq_23_in1
	// Insensitive connections
	always @(*) begin
		eq_23_in0 = valid ? 32'd4 : 32'd4;
		eq_23_in1 = valid ? global_state : global_state;
	end
	// controller for eq_231.eq_231_in0
	// controller for eq_231.eq_231_in1
	// Insensitive connections
	always @(*) begin
		eq_231_in0 = valid ? 32'd1 : 32'd1;
		eq_231_in1 = valid ? global_state : global_state;
	end
	// controller for eq_233.eq_233_in0
	// controller for eq_233.eq_233_in1
	// Insensitive connections
	always @(*) begin
		eq_233_in0 = valid ? 32'd2 : 32'd2;
		eq_233_in1 = valid ? global_state : global_state;
	end
	// controller for eq_236.eq_236_in0
	// controller for eq_236.eq_236_in1
	// Insensitive connections
	always @(*) begin
		eq_236_in0 = valid ? 32'd2 : 32'd2;
		eq_236_in1 = valid ? global_state : global_state;
	end
	// controller for eq_238.eq_238_in0
	// controller for eq_238.eq_238_in1
	// Insensitive connections
	always @(*) begin
		eq_238_in0 = valid ? 32'd3 : 32'd3;
		eq_238_in1 = valid ? global_state : global_state;
	end
	// controller for eq_241.eq_241_in0
	// controller for eq_241.eq_241_in1
	// Insensitive connections
	always @(*) begin
		eq_241_in0 = valid ? 32'd3 : 32'd3;
		eq_241_in1 = valid ? global_state : global_state;
	end
	// controller for eq_244.eq_244_in0
	// controller for eq_244.eq_244_in1
	// Insensitive connections
	always @(*) begin
		eq_244_in0 = valid ? 32'd4 : 32'd4;
		eq_244_in1 = valid ? global_state : global_state;
	end
	// controller for eq_247.eq_247_in0
	// controller for eq_247.eq_247_in1
	// Insensitive connections
	always @(*) begin
		eq_247_in0 = valid ? 32'd4 : 32'd4;
		eq_247_in1 = valid ? global_state : global_state;
	end
	// controller for eq_250.eq_250_in0
	// controller for eq_250.eq_250_in1
	// Insensitive connections
	always @(*) begin
		eq_250_in0 = valid ? 32'd4 : 32'd4;
		eq_250_in1 = valid ? global_state : global_state;
	end
	// controller for eq_253.eq_253_in0
	// controller for eq_253.eq_253_in1
	// Insensitive connections
	always @(*) begin
		eq_253_in0 = valid ? 32'd4 : 32'd4;
		eq_253_in1 = valid ? global_state : global_state;
	end
	// controller for eq_255.eq_255_in0
	// controller for eq_255.eq_255_in1
	// Insensitive connections
	always @(*) begin
		eq_255_in0 = valid ? 32'd4 : 32'd4;
		eq_255_in1 = valid ? global_state : global_state;
	end
	// controller for eq_258.eq_258_in0
	// controller for eq_258.eq_258_in1
	// Insensitive connections
	always @(*) begin
		eq_258_in0 = valid ? 32'd4 : 32'd4;
		eq_258_in1 = valid ? global_state : global_state;
	end
	// controller for eq_260.eq_260_in0
	// controller for eq_260.eq_260_in1
	// Insensitive connections
	always @(*) begin
		eq_260_in0 = valid ? 32'd1 : 32'd1;
		eq_260_in1 = valid ? global_state : global_state;
	end
	// controller for eq_262.eq_262_in0
	// controller for eq_262.eq_262_in1
	// Insensitive connections
	always @(*) begin
		eq_262_in0 = valid ? 32'd3 : 32'd3;
		eq_262_in1 = valid ? global_state : global_state;
	end
	// controller for eq_264.eq_264_in0
	// controller for eq_264.eq_264_in1
	// Insensitive connections
	always @(*) begin
		eq_264_in0 = valid ? 32'd3 : 32'd3;
		eq_264_in1 = valid ? global_state : global_state;
	end
	// controller for eq_266.eq_266_in0
	// controller for eq_266.eq_266_in1
	// Insensitive connections
	always @(*) begin
		eq_266_in0 = valid ? 32'd3 : 32'd3;
		eq_266_in1 = valid ? global_state : global_state;
	end
	// controller for eq_30.eq_30_in0
	// controller for eq_30.eq_30_in1
	// Insensitive connections
	always @(*) begin
		eq_30_in0 = valid ? 32'd4 : 32'd4;
		eq_30_in1 = valid ? global_state : global_state;
	end
	// controller for eq_34.eq_34_in0
	// controller for eq_34.eq_34_in1
	// Insensitive connections
	always @(*) begin
		eq_34_in0 = valid ? 32'd1 : 32'd1;
		eq_34_in1 = valid ? global_state : global_state;
	end
	// controller for eq_38.eq_38_in0
	// controller for eq_38.eq_38_in1
	// Insensitive connections
	always @(*) begin
		eq_38_in0 = valid ? 32'd1 : 32'd1;
		eq_38_in1 = valid ? global_state : global_state;
	end
	// controller for eq_4.eq_4_in0
	// controller for eq_4.eq_4_in1
	// Insensitive connections
	always @(*) begin
		eq_4_in0 = valid ? 32'd4 : 32'd4;
		eq_4_in1 = valid ? global_state : global_state;
	end
	// controller for eq_45.eq_45_in0
	// controller for eq_45.eq_45_in1
	// Insensitive connections
	always @(*) begin
		eq_45_in0 = valid ? 32'd3 : 32'd3;
		eq_45_in1 = valid ? global_state : global_state;
	end
	// controller for eq_49.eq_49_in0
	// controller for eq_49.eq_49_in1
	// Insensitive connections
	always @(*) begin
		eq_49_in0 = valid ? 32'd0 : 32'd0;
		eq_49_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_50.eq_50_in0
	// controller for eq_50.eq_50_in1
	// Insensitive connections
	always @(*) begin
		eq_50_in0 = valid ? 32'd1 : 32'd1;
		eq_50_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_52.eq_52_in0
	// controller for eq_52.eq_52_in1
	// Insensitive connections
	always @(*) begin
		eq_52_in0 = valid ? 32'd2 : 32'd2;
		eq_52_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_54.eq_54_in0
	// controller for eq_54.eq_54_in1
	// Insensitive connections
	always @(*) begin
		eq_54_in0 = valid ? 32'd3 : 32'd3;
		eq_54_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_56.eq_56_in0
	// controller for eq_56.eq_56_in1
	// Insensitive connections
	always @(*) begin
		eq_56_in0 = valid ? 32'd4 : 32'd4;
		eq_56_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_58.eq_58_in0
	// controller for eq_58.eq_58_in1
	// Insensitive connections
	always @(*) begin
		eq_58_in0 = valid ? 32'd5 : 32'd5;
		eq_58_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_60.eq_60_in0
	// controller for eq_60.eq_60_in1
	// Insensitive connections
	always @(*) begin
		eq_60_in0 = valid ? 32'd6 : 32'd6;
		eq_60_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_62.eq_62_in0
	// controller for eq_62.eq_62_in1
	// Insensitive connections
	always @(*) begin
		eq_62_in0 = valid ? 32'd7 : 32'd7;
		eq_62_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_64.eq_64_in0
	// controller for eq_64.eq_64_in1
	// Insensitive connections
	always @(*) begin
		eq_64_in0 = valid ? 32'd8 : 32'd8;
		eq_64_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_66.eq_66_in0
	// controller for eq_66.eq_66_in1
	// Insensitive connections
	always @(*) begin
		eq_66_in0 = valid ? 32'd9 : 32'd9;
		eq_66_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_68.eq_68_in0
	// controller for eq_68.eq_68_in1
	// Insensitive connections
	always @(*) begin
		eq_68_in0 = valid ? 32'd10 : 32'd10;
		eq_68_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_70.eq_70_in0
	// controller for eq_70.eq_70_in1
	// Insensitive connections
	always @(*) begin
		eq_70_in0 = valid ? 32'd0 : 32'd0;
		eq_70_in1 = valid ? global_state : global_state;
	end
	// controller for eq_72.eq_72_in0
	// controller for eq_72.eq_72_in1
	// Insensitive connections
	always @(*) begin
		eq_72_in0 = valid ? 32'd1 : 32'd1;
		eq_72_in1 = valid ? global_state : global_state;
	end
	// controller for eq_74.eq_74_in0
	// controller for eq_74.eq_74_in1
	// Insensitive connections
	always @(*) begin
		eq_74_in0 = valid ? 32'd2 : 32'd2;
		eq_74_in1 = valid ? global_state : global_state;
	end
	// controller for eq_76.eq_76_in0
	// controller for eq_76.eq_76_in1
	// Insensitive connections
	always @(*) begin
		eq_76_in0 = valid ? 32'd3 : 32'd3;
		eq_76_in1 = valid ? global_state : global_state;
	end
	// controller for eq_78.eq_78_in0
	// controller for eq_78.eq_78_in1
	// Insensitive connections
	always @(*) begin
		eq_78_in0 = valid ? 32'd4 : 32'd4;
		eq_78_in1 = valid ? global_state : global_state;
	end
	// controller for eq_8.eq_8_in0
	// controller for eq_8.eq_8_in1
	// Insensitive connections
	always @(*) begin
		eq_8_in0 = valid ? 32'd1 : 32'd1;
		eq_8_in1 = valid ? global_state : global_state;
	end
	// controller for eq_80.eq_80_in0
	// controller for eq_80.eq_80_in1
	// Insensitive connections
	always @(*) begin
		eq_80_in0 = valid ? 32'd0 : 32'd0;
		eq_80_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_81.eq_81_in0
	// controller for eq_81.eq_81_in1
	// Insensitive connections
	always @(*) begin
		eq_81_in0 = valid ? 32'd1 : 32'd1;
		eq_81_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_84.eq_84_in0
	// controller for eq_84.eq_84_in1
	// Insensitive connections
	always @(*) begin
		eq_84_in0 = valid ? 32'd2 : 32'd2;
		eq_84_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_87.eq_87_in0
	// controller for eq_87.eq_87_in1
	// Insensitive connections
	always @(*) begin
		eq_87_in0 = valid ? 32'd3 : 32'd3;
		eq_87_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_90.eq_90_in0
	// controller for eq_90.eq_90_in1
	// Insensitive connections
	always @(*) begin
		eq_90_in0 = valid ? 32'd4 : 32'd4;
		eq_90_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_93.eq_93_in0
	// controller for eq_93.eq_93_in1
	// Insensitive connections
	always @(*) begin
		eq_93_in0 = valid ? 32'd5 : 32'd5;
		eq_93_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_96.eq_96_in0
	// controller for eq_96.eq_96_in1
	// Insensitive connections
	always @(*) begin
		eq_96_in0 = valid ? 32'd6 : 32'd6;
		eq_96_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for eq_99.eq_99_in0
	// controller for eq_99.eq_99_in1
	// Insensitive connections
	always @(*) begin
		eq_99_in0 = valid ? 32'd7 : 32'd7;
		eq_99_in1 = valid ? global_next_block : global_next_block;
	end
	// controller for icmp_15.cmp_in0_icmp_15
	// controller for icmp_15.cmp_in1_icmp_15
	// Insensitive connections
	always @(*) begin
		cmp_in0_icmp_15 = valid ? add_out_add_14 : add_out_add_14;
		cmp_in1_icmp_15 = valid ? 32'd4 : 32'd4;
	end
	// controller for in.in_read_valid_reg
	always @(*) begin
		if (andOp_130_out) begin 
			in_read_valid_reg = -(1'd1);
		end else begin
			in_read_valid_reg = 0;
		end
	end
	// controller for notOp_100.notOp_100_in0
	// Insensitive connections
	always @(*) begin
		notOp_100_in0 = valid ? eq_99_out : eq_99_out;
	end
	// controller for notOp_103.notOp_103_in0
	// Insensitive connections
	always @(*) begin
		notOp_103_in0 = valid ? eq_102_out : eq_102_out;
	end
	// controller for notOp_106.notOp_106_in0
	// Insensitive connections
	always @(*) begin
		notOp_106_in0 = valid ? eq_105_out : eq_105_out;
	end
	// controller for notOp_109.notOp_109_in0
	// Insensitive connections
	always @(*) begin
		notOp_109_in0 = valid ? eq_108_out : eq_108_out;
	end
	// controller for notOp_11.notOp_11_in0
	// Insensitive connections
	always @(*) begin
		notOp_11_in0 = valid ? andOp_10_out : andOp_10_out;
	end
	// controller for notOp_15.notOp_15_in0
	// Insensitive connections
	always @(*) begin
		notOp_15_in0 = valid ? andOp_14_out : andOp_14_out;
	end
	// controller for notOp_155.notOp_155_in0
	// Insensitive connections
	always @(*) begin
		notOp_155_in0 = valid ? andOp_154_out : andOp_154_out;
	end
	// controller for notOp_161.notOp_161_in0
	// Insensitive connections
	always @(*) begin
		notOp_161_in0 = valid ? andOp_160_out : andOp_160_out;
	end
	// controller for notOp_167.notOp_167_in0
	// Insensitive connections
	always @(*) begin
		notOp_167_in0 = valid ? andOp_166_out : andOp_166_out;
	end
	// controller for notOp_17.notOp_17_in0
	// Insensitive connections
	always @(*) begin
		notOp_17_in0 = valid ? icmp_tmp_5 : icmp_tmp_5;
	end
	// controller for notOp_173.notOp_173_in0
	// Insensitive connections
	always @(*) begin
		notOp_173_in0 = valid ? andOp_172_out : andOp_172_out;
	end
	// controller for notOp_179.notOp_179_in0
	// Insensitive connections
	always @(*) begin
		notOp_179_in0 = valid ? andOp_178_out : andOp_178_out;
	end
	// controller for notOp_185.notOp_185_in0
	// Insensitive connections
	always @(*) begin
		notOp_185_in0 = valid ? andOp_184_out : andOp_184_out;
	end
	// controller for notOp_189.notOp_189_in0
	// Insensitive connections
	always @(*) begin
		notOp_189_in0 = valid ? andOp_188_out : andOp_188_out;
	end
	// controller for notOp_195.notOp_195_in0
	// Insensitive connections
	always @(*) begin
		notOp_195_in0 = valid ? andOp_194_out : andOp_194_out;
	end
	// controller for notOp_203.notOp_203_in0
	// Insensitive connections
	always @(*) begin
		notOp_203_in0 = valid ? andOp_202_out : andOp_202_out;
	end
	// controller for notOp_209.notOp_209_in0
	// Insensitive connections
	always @(*) begin
		notOp_209_in0 = valid ? andOp_208_out : andOp_208_out;
	end
	// controller for notOp_215.notOp_215_in0
	// Insensitive connections
	always @(*) begin
		notOp_215_in0 = valid ? andOp_214_out : andOp_214_out;
	end
	// controller for notOp_22.notOp_22_in0
	// Insensitive connections
	always @(*) begin
		notOp_22_in0 = valid ? andOp_21_out : andOp_21_out;
	end
	// controller for notOp_222.notOp_222_in0
	// Insensitive connections
	always @(*) begin
		notOp_222_in0 = valid ? in_read_ready : in_read_ready;
	end
	// controller for notOp_243.notOp_243_in0
	// Insensitive connections
	always @(*) begin
		notOp_243_in0 = valid ? icmp_tmp_5 : icmp_tmp_5;
	end
	// controller for notOp_249.notOp_249_in0
	// Insensitive connections
	always @(*) begin
		notOp_249_in0 = valid ? out_write_ready : out_write_ready;
	end
	// controller for notOp_26.notOp_26_in0
	// Insensitive connections
	always @(*) begin
		notOp_26_in0 = valid ? andOp_25_out : andOp_25_out;
	end
	// controller for notOp_28.notOp_28_in0
	// Insensitive connections
	always @(*) begin
		notOp_28_in0 = valid ? out_write_ready : out_write_ready;
	end
	// controller for notOp_3.notOp_3_in0
	// Insensitive connections
	always @(*) begin
		notOp_3_in0 = valid ? andOp_2_out : andOp_2_out;
	end
	// controller for notOp_33.notOp_33_in0
	// Insensitive connections
	always @(*) begin
		notOp_33_in0 = valid ? andOp_32_out : andOp_32_out;
	end
	// controller for notOp_37.notOp_37_in0
	// Insensitive connections
	always @(*) begin
		notOp_37_in0 = valid ? andOp_36_out : andOp_36_out;
	end
	// controller for notOp_41.notOp_41_in0
	// Insensitive connections
	always @(*) begin
		notOp_41_in0 = valid ? andOp_40_out : andOp_40_out;
	end
	// controller for notOp_43.notOp_43_in0
	// Insensitive connections
	always @(*) begin
		notOp_43_in0 = valid ? in_read_ready : in_read_ready;
	end
	// controller for notOp_48.notOp_48_in0
	// Insensitive connections
	always @(*) begin
		notOp_48_in0 = valid ? andOp_47_out : andOp_47_out;
	end
	// controller for notOp_7.notOp_7_in0
	// Insensitive connections
	always @(*) begin
		notOp_7_in0 = valid ? andOp_6_out : andOp_6_out;
	end
	// controller for notOp_82.notOp_82_in0
	// Insensitive connections
	always @(*) begin
		notOp_82_in0 = valid ? eq_81_out : eq_81_out;
	end
	// controller for notOp_85.notOp_85_in0
	// Insensitive connections
	always @(*) begin
		notOp_85_in0 = valid ? eq_84_out : eq_84_out;
	end
	// controller for notOp_88.notOp_88_in0
	// Insensitive connections
	always @(*) begin
		notOp_88_in0 = valid ? eq_87_out : eq_87_out;
	end
	// controller for notOp_91.notOp_91_in0
	// Insensitive connections
	always @(*) begin
		notOp_91_in0 = valid ? eq_90_out : eq_90_out;
	end
	// controller for notOp_94.notOp_94_in0
	// Insensitive connections
	always @(*) begin
		notOp_94_in0 = valid ? eq_93_out : eq_93_out;
	end
	// controller for notOp_97.notOp_97_in0
	// Insensitive connections
	always @(*) begin
		notOp_97_in0 = valid ? eq_96_out : eq_96_out;
	end
	// controller for orOp_51.orOp_51_in0
	// controller for orOp_51.orOp_51_in1
	// Insensitive connections
	always @(*) begin
		orOp_51_in0 = valid ? eq_50_out : eq_50_out;
		orOp_51_in1 = valid ? andOp_16_out : andOp_16_out;
	end
	// controller for orOp_53.orOp_53_in0
	// controller for orOp_53.orOp_53_in1
	// Insensitive connections
	always @(*) begin
		orOp_53_in0 = valid ? eq_52_out : eq_52_out;
		orOp_53_in1 = valid ? andOp_32_out : andOp_32_out;
	end
	// controller for orOp_55.orOp_55_in0
	// controller for orOp_55.orOp_55_in1
	// Insensitive connections
	always @(*) begin
		orOp_55_in0 = valid ? eq_54_out : eq_54_out;
		orOp_55_in1 = valid ? andOp_2_out : andOp_2_out;
	end
	// controller for orOp_57.orOp_57_in0
	// controller for orOp_57.orOp_57_in1
	// Insensitive connections
	always @(*) begin
		orOp_57_in0 = valid ? eq_56_out : eq_56_out;
		orOp_57_in1 = valid ? andOp_47_out : andOp_47_out;
	end
	// controller for orOp_59.orOp_59_in0
	// controller for orOp_59.orOp_59_in1
	// Insensitive connections
	always @(*) begin
		orOp_59_in0 = valid ? eq_58_out : eq_58_out;
		orOp_59_in1 = valid ? andOp_6_out : andOp_6_out;
	end
	// controller for orOp_61.orOp_61_in0
	// controller for orOp_61.orOp_61_in1
	// Insensitive connections
	always @(*) begin
		orOp_61_in0 = valid ? eq_60_out : eq_60_out;
		orOp_61_in1 = valid ? andOp_21_out : andOp_21_out;
	end
	// controller for orOp_63.orOp_63_in0
	// controller for orOp_63.orOp_63_in1
	// Insensitive connections
	always @(*) begin
		orOp_63_in0 = valid ? eq_62_out : eq_62_out;
		orOp_63_in1 = valid ? andOp_27_out : andOp_27_out;
	end
	// controller for orOp_65.orOp_65_in0
	// controller for orOp_65.orOp_65_in1
	// Insensitive connections
	always @(*) begin
		orOp_65_in0 = valid ? eq_64_out : eq_64_out;
		orOp_65_in1 = valid ? andOp_10_out : andOp_10_out;
	end
	// controller for orOp_67.orOp_67_in0
	// controller for orOp_67.orOp_67_in1
	// Insensitive connections
	always @(*) begin
		orOp_67_in0 = valid ? eq_66_out : eq_66_out;
		orOp_67_in1 = valid ? andOp_36_out : andOp_36_out;
	end
	// controller for orOp_69.orOp_69_in0
	// controller for orOp_69.orOp_69_in1
	// Insensitive connections
	always @(*) begin
		orOp_69_in0 = valid ? eq_68_out : eq_68_out;
		orOp_69_in1 = valid ? andOp_42_out : andOp_42_out;
	end
	// controller for out.out_in_data_reg
	always @(*) begin
		if (andOp_148_out) begin 
			out_in_data_reg = rdata_ram_0;
		end else begin
			out_in_data_reg = 0;
		end
	end
	// controller for out.out_write_valid_reg
	always @(*) begin
		if (andOp_146_out) begin 
			out_write_valid_reg = -(1'd1);
		end else begin
			out_write_valid_reg = 0;
		end
	end
	// controller for phi_6.phi_in_phi_6
	// controller for phi_6.phi_last_block_phi_6
	// controller for phi_6.phi_s_phi_6
	// Insensitive connections
	always @(*) begin
		phi_in_phi_6 = valid ? {32'd0, add_tmp_4} : {32'd0, add_tmp_4};
		phi_last_block_phi_6 = valid ? bb_3_predecessor_out_data : bb_3_predecessor_out_data;
		phi_s_phi_6 = valid ? {32'd0, 32'd4} : {32'd0, 32'd4};
	end
	// controller for ram_0.raddr_ram_0_reg
	always @(*) begin
		if (andOp_114_out) begin 
			raddr_ram_0_reg = 0;
		end else if (andOp_118_out) begin 
			raddr_ram_0_reg = 0;
		end else begin
			raddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.waddr_ram_0_reg
	always @(*) begin
		if (andOp_112_out) begin 
			waddr_ram_0_reg = 0;
		end else if (andOp_116_out) begin 
			waddr_ram_0_reg = 0;
		end else begin
			waddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wdata_ram_0_reg
	always @(*) begin
		if (andOp_112_out) begin 
			wdata_ram_0_reg = 32'd0;
		end else if (andOp_116_out) begin 
			wdata_ram_0_reg = add_out_add_12;
		end else begin
			wdata_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wen_ram_0_reg
	always @(*) begin
		if (andOp_112_out) begin 
			wen_ram_0_reg = 1;
		end else if (andOp_116_out) begin 
			wen_ram_0_reg = 1;
		end else begin
			wen_ram_0_reg = 0;
		end
	end
	// controller for ret_21.valid_reg
	always @(*) begin
		if (andOp_144_out) begin 
			valid_reg = 1;
		end else begin
			valid_reg = 0;
		end
	end
	// controller for tmp_output_135.tmp_output_135_in_data
	always @(*) begin
		if (eq_136_out) begin 
			tmp_output_135_in_data = in_out_data;
		end else begin
			tmp_output_135_in_data = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			add_tmp_4 <= 0;
		end else begin
			if (andOp_263_out) begin
				add_tmp_4 <= add_out_add_14;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			call_tmp_6 <= 0;
		end else begin
			if (andOp_267_out) begin
				call_tmp_6 <= in_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_next_block <= 0;
		end else begin
			if (andOp_18_out) begin
				global_next_block <= 32'd3;
			end
			if (andOp_29_out) begin
				global_next_block <= 32'd6;
			end
			if (andOp_44_out) begin
				global_next_block <= 32'd9;
			end
			if (andOp_71_out) begin
				global_next_block <= 32'd0;
			end
			if (andOp_73_out) begin
				global_next_block <= 32'd10;
			end
			if (andOp_75_out) begin
				global_next_block <= 32'd10;
			end
			if (andOp_77_out) begin
				global_next_block <= 32'd4;
			end
			if (andOp_79_out) begin
				global_next_block <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_221_out) begin
				global_state <= 32'd1;
			end
			if (andOp_227_out) begin
				global_state <= 32'd1;
			end
			if (andOp_232_out) begin
				global_state <= 32'd2;
			end
			if (andOp_237_out) begin
				global_state <= 32'd3;
			end
			if (andOp_242_out) begin
				global_state <= 32'd4;
			end
			if (andOp_248_out) begin
				global_state <= 32'd1;
			end
			if (andOp_254_out) begin
				global_state <= 32'd4;
			end
			if (andOp_259_out) begin
				global_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			icmp_tmp_5 <= 0;
		end else begin
			if (andOp_265_out) begin
				icmp_tmp_5 <= cmp_out_icmp_15;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			last_BB_reg <= 0;
		end else begin
			if (andOp_156_out) begin
				last_BB_reg <= 32'd3;
			end
			if (andOp_162_out) begin
				last_BB_reg <= 32'd0;
			end
			if (andOp_168_out) begin
				last_BB_reg <= 32'd9;
			end
			if (andOp_174_out) begin
				last_BB_reg <= 32'd8;
			end
			if (andOp_180_out) begin
				last_BB_reg <= 32'd10;
			end
			if (andOp_190_out) begin
				last_BB_reg <= 32'd4;
			end
			if (andOp_196_out) begin
				last_BB_reg <= 32'd1;
			end
			if (andOp_198_out) begin
				last_BB_reg <= 32'd2;
			end
			if (andOp_204_out) begin
				last_BB_reg <= 32'd5;
			end
			if (andOp_210_out) begin
				last_BB_reg <= 32'd7;
			end
			if (andOp_216_out) begin
				last_BB_reg <= 32'd6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			phi_tmp_0 <= 0;
		end else begin
			if (andOp_261_out) begin
				phi_tmp_0 <= phi_out_phi_6;
			end
		end
	end

endmodule

