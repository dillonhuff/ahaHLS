module channel_reduce_4(input [0:0] clk, input [0:0] rst, output [31:0] in_in_data, output [0:0] in_read_valid, output [0:0] in_rst, output [0:0] in_write_valid, input [31:0] in_out_data, input [0:0] in_read_ready, input [0:0] in_write_ready, output [31:0] out_in_data, output [0:0] out_read_valid, output [0:0] out_rst, output [0:0] out_write_valid, input [31:0] out_out_data, input [0:0] out_read_ready, input [0:0] out_write_ready, output [0:0] valid);

	reg [31:0] in_in_data_reg;
	reg [0:0] in_read_valid_reg;
	reg [0:0] in_rst_reg;
	reg [0:0] in_write_valid_reg;
	reg [31:0] out_in_data_reg;
	reg [0:0] out_read_valid_reg;
	reg [0:0] out_rst_reg;
	reg [0:0] out_write_valid_reg;
	reg [0:0] valid_reg;

	assign in_in_data = in_in_data_reg;
	assign in_read_valid = in_read_valid_reg;
	assign in_rst = in_rst_reg;
	assign in_write_valid = in_write_valid_reg;
	assign out_in_data = out_in_data_reg;
	assign out_read_valid = out_read_valid_reg;
	assign out_rst = out_rst_reg;
	assign out_write_valid = out_write_valid_reg;
	assign valid = valid_reg;

	// Start debug wires and ports

	initial begin
	end





	// End debug wires and ports

	// Start Functional Units
	br_dummy br_unit();

	add alloca_0();

	add bitcast_1();

	add call_2();

	reg [31:0] raddr_ram_0_reg;
	reg [31:0] waddr_ram_0_reg;
	reg [31:0] wdata_ram_0_reg;
	reg [0:0] wen_ram_0_reg;
	wire [31:0] rdata_ram_0;
	register #(.WIDTH(32)) ram_0(.clk(clk), .raddr(raddr_ram_0_reg), .rdata(rdata_ram_0), .rst(rst), .waddr(waddr_ram_0_reg), .wdata(wdata_ram_0_reg), .wen(wen_ram_0_reg));

	add call_22();

	reg [63:0] phi_in_phi_7;
	reg [31:0] phi_last_block_phi_7;
	reg [63:0] phi_s_phi_7;
	wire [31:0] phi_out_phi_7;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_7(.in(phi_in_phi_7), .last_block(phi_last_block_phi_7), .out(phi_out_phi_7), .s(phi_s_phi_7));

	reg [31:0] add_in0_add_14;
	reg [31:0] add_in1_add_14;
	wire [31:0] add_out_add_14;
	add #(.WIDTH(32)) add_add_14(.in0(add_in0_add_14), .in1(add_in1_add_14), .out(add_out_add_14));

	reg [31:0] add_in0_add_16;
	reg [31:0] add_in1_add_16;
	wire [31:0] add_out_add_16;
	add #(.WIDTH(32)) add_add_16(.in0(add_in0_add_16), .in1(add_in1_add_16), .out(add_out_add_16));

	reg [31:0] cmp_in0_icmp_17;
	reg [31:0] cmp_in1_icmp_17;
	wire [0:0] cmp_out_icmp_17;
	eq #(.WIDTH(32)) icmp_17(.in0(cmp_in0_icmp_17), .in1(cmp_in1_icmp_17), .out(cmp_out_icmp_17));

	reg [0:0] data_in_0_1_in_data;
	wire [0:0] data_in_0_1_out_data;
	hls_wire #(.WIDTH(1)) data_in_0_1(.in_data(data_in_0_1_in_data), .out_data(data_in_0_1_out_data));

	reg [31:0] data_in_0_3_in_data;
	wire [31:0] data_in_0_3_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_3(.in_data(data_in_0_3_in_data), .out_data(data_in_0_3_out_data));

	reg [31:0] data_in_0_5_in_data;
	wire [31:0] data_in_0_5_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_5(.in_data(data_in_0_5_in_data), .out_data(data_in_0_5_out_data));

	reg [31:0] data_in_0_7_in_data;
	wire [31:0] data_in_0_7_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_7(.in_data(data_in_0_7_in_data), .out_data(data_in_0_7_out_data));

	reg [31:0] data_in_0_9_in_data;
	wire [31:0] data_in_0_9_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_9(.in_data(data_in_0_9_in_data), .out_data(data_in_0_9_out_data));

	reg [31:0] data_in_0_11_in_data;
	wire [31:0] data_in_0_11_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_11(.in_data(data_in_0_11_in_data), .out_data(data_in_0_11_out_data));

	reg [0:0] data_in_0_13_in_data;
	wire [0:0] data_in_0_13_out_data;
	hls_wire #(.WIDTH(1)) data_in_0_13(.in_data(data_in_0_13_in_data), .out_data(data_in_0_13_out_data));

	reg [31:0] data_in_0_15_in_data;
	wire [31:0] data_in_0_15_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_15(.in_data(data_in_0_15_in_data), .out_data(data_in_0_15_out_data));

	reg [0:0] data_in_0_17_in_data;
	wire [0:0] data_in_0_17_out_data;
	hls_wire #(.WIDTH(1)) data_in_0_17(.in_data(data_in_0_17_in_data), .out_data(data_in_0_17_out_data));

	reg [0:0] data_in_1_19_in_data;
	wire [0:0] data_in_1_19_out_data;
	hls_wire #(.WIDTH(1)) data_in_1_19(.in_data(data_in_1_19_in_data), .out_data(data_in_1_19_out_data));

	reg [31:0] data_in_1_21_in_data;
	wire [31:0] data_in_1_21_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_21(.in_data(data_in_1_21_in_data), .out_data(data_in_1_21_out_data));

	reg [31:0] data_in_1_23_in_data;
	wire [31:0] data_in_1_23_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_23(.in_data(data_in_1_23_in_data), .out_data(data_in_1_23_out_data));

	reg [31:0] data_in_1_25_in_data;
	wire [31:0] data_in_1_25_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_25(.in_data(data_in_1_25_in_data), .out_data(data_in_1_25_out_data));

	reg [31:0] data_in_1_27_in_data;
	wire [31:0] data_in_1_27_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_27(.in_data(data_in_1_27_in_data), .out_data(data_in_1_27_out_data));

	reg [31:0] data_in_1_29_in_data;
	wire [31:0] data_in_1_29_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_29(.in_data(data_in_1_29_in_data), .out_data(data_in_1_29_out_data));

	reg [0:0] data_in_1_31_in_data;
	wire [0:0] data_in_1_31_out_data;
	hls_wire #(.WIDTH(1)) data_in_1_31(.in_data(data_in_1_31_in_data), .out_data(data_in_1_31_out_data));

	reg [31:0] data_in_1_33_in_data;
	wire [31:0] data_in_1_33_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_33(.in_data(data_in_1_33_in_data), .out_data(data_in_1_33_out_data));

	reg [0:0] data_in_1_35_in_data;
	wire [0:0] data_in_1_35_out_data;
	hls_wire #(.WIDTH(1)) data_in_1_35(.in_data(data_in_1_35_in_data), .out_data(data_in_1_35_out_data));

	reg [0:0] data_in_2_37_in_data;
	wire [0:0] data_in_2_37_out_data;
	hls_wire #(.WIDTH(1)) data_in_2_37(.in_data(data_in_2_37_in_data), .out_data(data_in_2_37_out_data));

	reg [31:0] data_in_2_39_in_data;
	wire [31:0] data_in_2_39_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_39(.in_data(data_in_2_39_in_data), .out_data(data_in_2_39_out_data));

	reg [31:0] data_in_2_41_in_data;
	wire [31:0] data_in_2_41_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_41(.in_data(data_in_2_41_in_data), .out_data(data_in_2_41_out_data));

	reg [31:0] data_in_2_43_in_data;
	wire [31:0] data_in_2_43_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_43(.in_data(data_in_2_43_in_data), .out_data(data_in_2_43_out_data));

	reg [31:0] data_in_2_45_in_data;
	wire [31:0] data_in_2_45_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_45(.in_data(data_in_2_45_in_data), .out_data(data_in_2_45_out_data));

	reg [31:0] data_in_2_47_in_data;
	wire [31:0] data_in_2_47_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_47(.in_data(data_in_2_47_in_data), .out_data(data_in_2_47_out_data));

	reg [0:0] data_in_2_49_in_data;
	wire [0:0] data_in_2_49_out_data;
	hls_wire #(.WIDTH(1)) data_in_2_49(.in_data(data_in_2_49_in_data), .out_data(data_in_2_49_out_data));

	reg [31:0] data_in_2_51_in_data;
	wire [31:0] data_in_2_51_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_51(.in_data(data_in_2_51_in_data), .out_data(data_in_2_51_out_data));

	reg [0:0] data_in_2_53_in_data;
	wire [0:0] data_in_2_53_out_data;
	hls_wire #(.WIDTH(1)) data_in_2_53(.in_data(data_in_2_53_in_data), .out_data(data_in_2_53_out_data));

	reg [0:0] data_in_3_55_in_data;
	wire [0:0] data_in_3_55_out_data;
	hls_wire #(.WIDTH(1)) data_in_3_55(.in_data(data_in_3_55_in_data), .out_data(data_in_3_55_out_data));

	reg [31:0] data_in_3_57_in_data;
	wire [31:0] data_in_3_57_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_57(.in_data(data_in_3_57_in_data), .out_data(data_in_3_57_out_data));

	reg [31:0] data_in_3_59_in_data;
	wire [31:0] data_in_3_59_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_59(.in_data(data_in_3_59_in_data), .out_data(data_in_3_59_out_data));

	reg [31:0] data_in_3_61_in_data;
	wire [31:0] data_in_3_61_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_61(.in_data(data_in_3_61_in_data), .out_data(data_in_3_61_out_data));

	reg [31:0] data_in_3_63_in_data;
	wire [31:0] data_in_3_63_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_63(.in_data(data_in_3_63_in_data), .out_data(data_in_3_63_out_data));

	reg [31:0] data_in_3_65_in_data;
	wire [31:0] data_in_3_65_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_65(.in_data(data_in_3_65_in_data), .out_data(data_in_3_65_out_data));

	reg [0:0] data_in_3_67_in_data;
	wire [0:0] data_in_3_67_out_data;
	hls_wire #(.WIDTH(1)) data_in_3_67(.in_data(data_in_3_67_in_data), .out_data(data_in_3_67_out_data));

	reg [31:0] data_in_3_69_in_data;
	wire [31:0] data_in_3_69_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_69(.in_data(data_in_3_69_in_data), .out_data(data_in_3_69_out_data));

	reg [0:0] data_in_3_71_in_data;
	wire [0:0] data_in_3_71_out_data;
	hls_wire #(.WIDTH(1)) data_in_3_71(.in_data(data_in_3_71_in_data), .out_data(data_in_3_71_out_data));

	reg [0:0] data_in_4_73_in_data;
	wire [0:0] data_in_4_73_out_data;
	hls_wire #(.WIDTH(1)) data_in_4_73(.in_data(data_in_4_73_in_data), .out_data(data_in_4_73_out_data));

	reg [31:0] data_in_4_75_in_data;
	wire [31:0] data_in_4_75_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_75(.in_data(data_in_4_75_in_data), .out_data(data_in_4_75_out_data));

	reg [31:0] data_in_4_77_in_data;
	wire [31:0] data_in_4_77_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_77(.in_data(data_in_4_77_in_data), .out_data(data_in_4_77_out_data));

	reg [31:0] data_in_4_79_in_data;
	wire [31:0] data_in_4_79_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_79(.in_data(data_in_4_79_in_data), .out_data(data_in_4_79_out_data));

	reg [31:0] data_in_4_81_in_data;
	wire [31:0] data_in_4_81_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_81(.in_data(data_in_4_81_in_data), .out_data(data_in_4_81_out_data));

	reg [31:0] data_in_4_83_in_data;
	wire [31:0] data_in_4_83_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_83(.in_data(data_in_4_83_in_data), .out_data(data_in_4_83_out_data));

	reg [0:0] data_in_4_85_in_data;
	wire [0:0] data_in_4_85_out_data;
	hls_wire #(.WIDTH(1)) data_in_4_85(.in_data(data_in_4_85_in_data), .out_data(data_in_4_85_out_data));

	reg [31:0] data_in_4_87_in_data;
	wire [31:0] data_in_4_87_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_87(.in_data(data_in_4_87_in_data), .out_data(data_in_4_87_out_data));

	reg [0:0] data_in_4_89_in_data;
	wire [0:0] data_in_4_89_out_data;
	hls_wire #(.WIDTH(1)) data_in_4_89(.in_data(data_in_4_89_in_data), .out_data(data_in_4_89_out_data));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] bb_8_active_in_state_1_in_data;
	wire [0:0] bb_8_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active_in_state_1(.in_data(bb_8_active_in_state_1_in_data), .out_data(bb_8_active_in_state_1_out_data));

	reg [31:0] bb_8_predecessor_in_state_1_in_data;
	wire [31:0] bb_8_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor_in_state_1(.in_data(bb_8_predecessor_in_state_1_in_data), .out_data(bb_8_predecessor_in_state_1_out_data));

	reg [0:0] bb_0_active_in_state_1_in_data;
	wire [0:0] bb_0_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_1(.in_data(bb_0_active_in_state_1_in_data), .out_data(bb_0_active_in_state_1_out_data));

	reg [31:0] bb_0_predecessor_in_state_1_in_data;
	wire [31:0] bb_0_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_1(.in_data(bb_0_predecessor_in_state_1_in_data), .out_data(bb_0_predecessor_in_state_1_out_data));

	reg [0:0] bb_3_active_in_state_1_in_data;
	wire [0:0] bb_3_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_1(.in_data(bb_3_active_in_state_1_in_data), .out_data(bb_3_active_in_state_1_out_data));

	reg [31:0] bb_3_predecessor_in_state_1_in_data;
	wire [31:0] bb_3_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_1(.in_data(bb_3_predecessor_in_state_1_in_data), .out_data(bb_3_predecessor_in_state_1_out_data));

	reg [0:0] bb_9_active_in_state_1_in_data;
	wire [0:0] bb_9_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_9_active_in_state_1(.in_data(bb_9_active_in_state_1_in_data), .out_data(bb_9_active_in_state_1_out_data));

	reg [31:0] bb_9_predecessor_in_state_1_in_data;
	wire [31:0] bb_9_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_9_predecessor_in_state_1(.in_data(bb_9_predecessor_in_state_1_in_data), .out_data(bb_9_predecessor_in_state_1_out_data));

	reg [0:0] bb_10_active_in_state_2_in_data;
	wire [0:0] bb_10_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_2(.in_data(bb_10_active_in_state_2_in_data), .out_data(bb_10_active_in_state_2_out_data));

	reg [31:0] bb_10_predecessor_in_state_2_in_data;
	wire [31:0] bb_10_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_2(.in_data(bb_10_predecessor_in_state_2_in_data), .out_data(bb_10_predecessor_in_state_2_out_data));

	reg [0:0] bb_4_active_in_state_3_in_data;
	wire [0:0] bb_4_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_3(.in_data(bb_4_active_in_state_3_in_data), .out_data(bb_4_active_in_state_3_out_data));

	reg [31:0] bb_4_predecessor_in_state_3_in_data;
	wire [31:0] bb_4_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_3(.in_data(bb_4_predecessor_in_state_3_in_data), .out_data(bb_4_predecessor_in_state_3_out_data));

	reg [0:0] bb_10_active_in_state_3_in_data;
	wire [0:0] bb_10_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_3(.in_data(bb_10_active_in_state_3_in_data), .out_data(bb_10_active_in_state_3_out_data));

	reg [31:0] bb_10_predecessor_in_state_3_in_data;
	wire [31:0] bb_10_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_3(.in_data(bb_10_predecessor_in_state_3_in_data), .out_data(bb_10_predecessor_in_state_3_out_data));

	reg [0:0] bb_5_active_in_state_4_in_data;
	wire [0:0] bb_5_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_5_active_in_state_4(.in_data(bb_5_active_in_state_4_in_data), .out_data(bb_5_active_in_state_4_out_data));

	reg [31:0] bb_5_predecessor_in_state_4_in_data;
	wire [31:0] bb_5_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_5_predecessor_in_state_4(.in_data(bb_5_predecessor_in_state_4_in_data), .out_data(bb_5_predecessor_in_state_4_out_data));

	reg [0:0] bb_6_active_in_state_4_in_data;
	wire [0:0] bb_6_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_6_active_in_state_4(.in_data(bb_6_active_in_state_4_in_data), .out_data(bb_6_active_in_state_4_out_data));

	reg [31:0] bb_6_predecessor_in_state_4_in_data;
	wire [31:0] bb_6_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_6_predecessor_in_state_4(.in_data(bb_6_predecessor_in_state_4_in_data), .out_data(bb_6_predecessor_in_state_4_out_data));

	reg [0:0] bb_7_active_in_state_4_in_data;
	wire [0:0] bb_7_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_7_active_in_state_4(.in_data(bb_7_active_in_state_4_in_data), .out_data(bb_7_active_in_state_4_out_data));

	reg [31:0] bb_7_predecessor_in_state_4_in_data;
	wire [31:0] bb_7_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_7_predecessor_in_state_4(.in_data(bb_7_predecessor_in_state_4_in_data), .out_data(bb_7_predecessor_in_state_4_out_data));

	reg [0:0] bb_4_active_in_state_4_in_data;
	wire [0:0] bb_4_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_4(.in_data(bb_4_active_in_state_4_in_data), .out_data(bb_4_active_in_state_4_out_data));

	reg [31:0] bb_4_predecessor_in_state_4_in_data;
	wire [31:0] bb_4_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_4(.in_data(bb_4_predecessor_in_state_4_in_data), .out_data(bb_4_predecessor_in_state_4_out_data));

	reg [0:0] bb_2_active_in_state_4_in_data;
	wire [0:0] bb_2_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_4(.in_data(bb_2_active_in_state_4_in_data), .out_data(bb_2_active_in_state_4_out_data));

	reg [31:0] bb_2_predecessor_in_state_4_in_data;
	wire [31:0] bb_2_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_4(.in_data(bb_2_predecessor_in_state_4_in_data), .out_data(bb_2_predecessor_in_state_4_out_data));

	reg [0:0] bb_1_active_in_state_4_in_data;
	wire [0:0] bb_1_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_4(.in_data(bb_1_active_in_state_4_in_data), .out_data(bb_1_active_in_state_4_out_data));

	reg [31:0] bb_1_predecessor_in_state_4_in_data;
	wire [31:0] bb_1_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_4(.in_data(bb_1_predecessor_in_state_4_in_data), .out_data(bb_1_predecessor_in_state_4_out_data));

	reg [0:0] andOp_90_in0;
	reg [0:0] andOp_90_in1;
	wire [0:0] andOp_90_out;
	andOp #(.WIDTH(1)) andOp_90(.in0(andOp_90_in0), .in1(andOp_90_in1), .out(andOp_90_out));

	reg [0:0] andOp_91_in0;
	reg [0:0] andOp_91_in1;
	wire [0:0] andOp_91_out;
	andOp #(.WIDTH(1)) andOp_91(.in0(andOp_91_in0), .in1(andOp_91_in1), .out(andOp_91_out));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] notOp_92_in0;
	wire [0:0] notOp_92_out;
	notOp #(.WIDTH(1)) notOp_92(.in(notOp_92_in0), .out(notOp_92_out));

	reg [0:0] andOp_93_in0;
	reg [0:0] andOp_93_in1;
	wire [0:0] andOp_93_out;
	andOp #(.WIDTH(1)) andOp_93(.in0(andOp_93_in0), .in1(andOp_93_in1), .out(andOp_93_out));

	reg [0:0] andOp_94_in0;
	reg [0:0] andOp_94_in1;
	wire [0:0] andOp_94_out;
	andOp #(.WIDTH(1)) andOp_94(.in0(andOp_94_in0), .in1(andOp_94_in1), .out(andOp_94_out));

	reg [0:0] br_8_happened_in_state_1_in_data;
	wire [0:0] br_8_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_8_happened_in_state_1(.in_data(br_8_happened_in_state_1_in_data), .out_data(br_8_happened_in_state_1_out_data));

	reg [0:0] notOp_95_in0;
	wire [0:0] notOp_95_out;
	notOp #(.WIDTH(1)) notOp_95(.in(notOp_95_in0), .out(notOp_95_out));

	reg [0:0] andOp_96_in0;
	reg [0:0] andOp_96_in1;
	wire [0:0] andOp_96_out;
	andOp #(.WIDTH(1)) andOp_96(.in0(andOp_96_in0), .in1(andOp_96_in1), .out(andOp_96_out));

	reg [0:0] andOp_97_in0;
	reg [0:0] andOp_97_in1;
	wire [0:0] andOp_97_out;
	andOp #(.WIDTH(1)) andOp_97(.in0(andOp_97_in0), .in1(andOp_97_in1), .out(andOp_97_out));

	reg [0:0] br_0_happened_in_state_1_in_data;
	wire [0:0] br_0_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_1(.in_data(br_0_happened_in_state_1_in_data), .out_data(br_0_happened_in_state_1_out_data));

	reg [0:0] notOp_98_in0;
	wire [0:0] notOp_98_out;
	notOp #(.WIDTH(1)) notOp_98(.in(notOp_98_in0), .out(notOp_98_out));

	reg [0:0] andOp_99_in0;
	reg [0:0] andOp_99_in1;
	wire [0:0] andOp_99_out;
	andOp #(.WIDTH(1)) andOp_99(.in0(andOp_99_in0), .in1(andOp_99_in1), .out(andOp_99_out));

	reg [0:0] andOp_100_in0;
	reg [0:0] andOp_100_in1;
	wire [0:0] andOp_100_out;
	andOp #(.WIDTH(1)) andOp_100(.in0(andOp_100_in0), .in1(andOp_100_in1), .out(andOp_100_out));

	reg [0:0] br_3_happened_in_state_1_in_data;
	wire [0:0] br_3_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_1(.in_data(br_3_happened_in_state_1_in_data), .out_data(br_3_happened_in_state_1_out_data));

	reg [0:0] notOp_101_in0;
	wire [0:0] notOp_101_out;
	notOp #(.WIDTH(1)) notOp_101(.in(notOp_101_in0), .out(notOp_101_out));

	reg [0:0] andOp_102_in0;
	reg [0:0] andOp_102_in1;
	wire [0:0] andOp_102_out;
	andOp #(.WIDTH(1)) andOp_102(.in0(andOp_102_in0), .in1(andOp_102_in1), .out(andOp_102_out));

	reg [0:0] andOp_103_in0;
	reg [0:0] andOp_103_in1;
	wire [0:0] andOp_103_out;
	andOp #(.WIDTH(1)) andOp_103(.in0(andOp_103_in0), .in1(andOp_103_in1), .out(andOp_103_out));

	reg [0:0] br_9_happened_in_state_1_in_data;
	wire [0:0] br_9_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_9_happened_in_state_1(.in_data(br_9_happened_in_state_1_in_data), .out_data(br_9_happened_in_state_1_out_data));

	reg [0:0] notOp_104_in0;
	wire [0:0] notOp_104_out;
	notOp #(.WIDTH(1)) notOp_104(.in(notOp_104_in0), .out(notOp_104_out));

	reg [0:0] andOp_105_in0;
	reg [0:0] andOp_105_in1;
	wire [0:0] andOp_105_out;
	andOp #(.WIDTH(1)) andOp_105(.in0(andOp_105_in0), .in1(andOp_105_in1), .out(andOp_105_out));

	reg [0:0] notOp_106_in0;
	wire [0:0] notOp_106_out;
	notOp #(.WIDTH(1)) notOp_106(.in(notOp_106_in0), .out(notOp_106_out));

	reg [0:0] andOp_107_in0;
	reg [0:0] andOp_107_in1;
	wire [0:0] andOp_107_out;
	andOp #(.WIDTH(1)) andOp_107(.in0(andOp_107_in0), .in1(andOp_107_in1), .out(andOp_107_out));

	reg [0:0] andOp_108_in0;
	reg [0:0] andOp_108_in1;
	wire [0:0] andOp_108_out;
	andOp #(.WIDTH(1)) andOp_108(.in0(andOp_108_in0), .in1(andOp_108_in1), .out(andOp_108_out));

	reg [0:0] andOp_109_in0;
	reg [0:0] andOp_109_in1;
	wire [0:0] andOp_109_out;
	andOp #(.WIDTH(1)) andOp_109(.in0(andOp_109_in0), .in1(andOp_109_in1), .out(andOp_109_out));

	reg [0:0] br_10_happened_in_state_2_in_data;
	wire [0:0] br_10_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_2(.in_data(br_10_happened_in_state_2_in_data), .out_data(br_10_happened_in_state_2_out_data));

	reg [0:0] notOp_110_in0;
	wire [0:0] notOp_110_out;
	notOp #(.WIDTH(1)) notOp_110(.in(notOp_110_in0), .out(notOp_110_out));

	reg [0:0] andOp_111_in0;
	reg [0:0] andOp_111_in1;
	wire [0:0] andOp_111_out;
	andOp #(.WIDTH(1)) andOp_111(.in0(andOp_111_in0), .in1(andOp_111_in1), .out(andOp_111_out));

	reg [0:0] andOp_112_in0;
	reg [0:0] andOp_112_in1;
	wire [0:0] andOp_112_out;
	andOp #(.WIDTH(1)) andOp_112(.in0(andOp_112_in0), .in1(andOp_112_in1), .out(andOp_112_out));

	reg [0:0] br_4_happened_in_state_3_in_data;
	wire [0:0] br_4_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_3(.in_data(br_4_happened_in_state_3_in_data), .out_data(br_4_happened_in_state_3_out_data));

	reg [0:0] notOp_113_in0;
	wire [0:0] notOp_113_out;
	notOp #(.WIDTH(1)) notOp_113(.in(notOp_113_in0), .out(notOp_113_out));

	reg [0:0] andOp_114_in0;
	reg [0:0] andOp_114_in1;
	wire [0:0] andOp_114_out;
	andOp #(.WIDTH(1)) andOp_114(.in0(andOp_114_in0), .in1(andOp_114_in1), .out(andOp_114_out));

	reg [0:0] notOp_115_in0;
	wire [0:0] notOp_115_out;
	notOp #(.WIDTH(1)) notOp_115(.in(notOp_115_in0), .out(notOp_115_out));

	reg [0:0] andOp_116_in0;
	reg [0:0] andOp_116_in1;
	wire [0:0] andOp_116_out;
	andOp #(.WIDTH(1)) andOp_116(.in0(andOp_116_in0), .in1(andOp_116_in1), .out(andOp_116_out));

	reg [0:0] andOp_117_in0;
	reg [0:0] andOp_117_in1;
	wire [0:0] andOp_117_out;
	andOp #(.WIDTH(1)) andOp_117(.in0(andOp_117_in0), .in1(andOp_117_in1), .out(andOp_117_out));

	reg [0:0] andOp_118_in0;
	reg [0:0] andOp_118_in1;
	wire [0:0] andOp_118_out;
	andOp #(.WIDTH(1)) andOp_118(.in0(andOp_118_in0), .in1(andOp_118_in1), .out(andOp_118_out));

	reg [0:0] br_10_happened_in_state_3_in_data;
	wire [0:0] br_10_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_3(.in_data(br_10_happened_in_state_3_in_data), .out_data(br_10_happened_in_state_3_out_data));

	reg [0:0] notOp_119_in0;
	wire [0:0] notOp_119_out;
	notOp #(.WIDTH(1)) notOp_119(.in(notOp_119_in0), .out(notOp_119_out));

	reg [0:0] andOp_120_in0;
	reg [0:0] andOp_120_in1;
	wire [0:0] andOp_120_out;
	andOp #(.WIDTH(1)) andOp_120(.in0(andOp_120_in0), .in1(andOp_120_in1), .out(andOp_120_out));

	reg [0:0] andOp_121_in0;
	reg [0:0] andOp_121_in1;
	wire [0:0] andOp_121_out;
	andOp #(.WIDTH(1)) andOp_121(.in0(andOp_121_in0), .in1(andOp_121_in1), .out(andOp_121_out));

	reg [0:0] br_5_happened_in_state_4_in_data;
	wire [0:0] br_5_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_5_happened_in_state_4(.in_data(br_5_happened_in_state_4_in_data), .out_data(br_5_happened_in_state_4_out_data));

	reg [0:0] notOp_122_in0;
	wire [0:0] notOp_122_out;
	notOp #(.WIDTH(1)) notOp_122(.in(notOp_122_in0), .out(notOp_122_out));

	reg [0:0] andOp_123_in0;
	reg [0:0] andOp_123_in1;
	wire [0:0] andOp_123_out;
	andOp #(.WIDTH(1)) andOp_123(.in0(andOp_123_in0), .in1(andOp_123_in1), .out(andOp_123_out));

	reg [0:0] andOp_124_in0;
	reg [0:0] andOp_124_in1;
	wire [0:0] andOp_124_out;
	andOp #(.WIDTH(1)) andOp_124(.in0(andOp_124_in0), .in1(andOp_124_in1), .out(andOp_124_out));

	reg [0:0] br_6_happened_in_state_4_in_data;
	wire [0:0] br_6_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_6_happened_in_state_4(.in_data(br_6_happened_in_state_4_in_data), .out_data(br_6_happened_in_state_4_out_data));

	reg [0:0] notOp_125_in0;
	wire [0:0] notOp_125_out;
	notOp #(.WIDTH(1)) notOp_125(.in(notOp_125_in0), .out(notOp_125_out));

	reg [0:0] andOp_126_in0;
	reg [0:0] andOp_126_in1;
	wire [0:0] andOp_126_out;
	andOp #(.WIDTH(1)) andOp_126(.in0(andOp_126_in0), .in1(andOp_126_in1), .out(andOp_126_out));

	reg [0:0] notOp_127_in0;
	wire [0:0] notOp_127_out;
	notOp #(.WIDTH(1)) notOp_127(.in(notOp_127_in0), .out(notOp_127_out));

	reg [0:0] andOp_128_in0;
	reg [0:0] andOp_128_in1;
	wire [0:0] andOp_128_out;
	andOp #(.WIDTH(1)) andOp_128(.in0(andOp_128_in0), .in1(andOp_128_in1), .out(andOp_128_out));

	reg [0:0] andOp_129_in0;
	reg [0:0] andOp_129_in1;
	wire [0:0] andOp_129_out;
	andOp #(.WIDTH(1)) andOp_129(.in0(andOp_129_in0), .in1(andOp_129_in1), .out(andOp_129_out));

	reg [0:0] andOp_130_in0;
	reg [0:0] andOp_130_in1;
	wire [0:0] andOp_130_out;
	andOp #(.WIDTH(1)) andOp_130(.in0(andOp_130_in0), .in1(andOp_130_in1), .out(andOp_130_out));

	reg [0:0] br_7_happened_in_state_4_in_data;
	wire [0:0] br_7_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_7_happened_in_state_4(.in_data(br_7_happened_in_state_4_in_data), .out_data(br_7_happened_in_state_4_out_data));

	reg [0:0] notOp_131_in0;
	wire [0:0] notOp_131_out;
	notOp #(.WIDTH(1)) notOp_131(.in(notOp_131_in0), .out(notOp_131_out));

	reg [0:0] andOp_132_in0;
	reg [0:0] andOp_132_in1;
	wire [0:0] andOp_132_out;
	andOp #(.WIDTH(1)) andOp_132(.in0(andOp_132_in0), .in1(andOp_132_in1), .out(andOp_132_out));

	reg [0:0] andOp_133_in0;
	reg [0:0] andOp_133_in1;
	wire [0:0] andOp_133_out;
	andOp #(.WIDTH(1)) andOp_133(.in0(andOp_133_in0), .in1(andOp_133_in1), .out(andOp_133_out));

	reg [0:0] br_4_happened_in_state_4_in_data;
	wire [0:0] br_4_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_4(.in_data(br_4_happened_in_state_4_in_data), .out_data(br_4_happened_in_state_4_out_data));

	reg [0:0] notOp_134_in0;
	wire [0:0] notOp_134_out;
	notOp #(.WIDTH(1)) notOp_134(.in(notOp_134_in0), .out(notOp_134_out));

	reg [0:0] andOp_135_in0;
	reg [0:0] andOp_135_in1;
	wire [0:0] andOp_135_out;
	andOp #(.WIDTH(1)) andOp_135(.in0(andOp_135_in0), .in1(andOp_135_in1), .out(andOp_135_out));

	reg [0:0] notOp_136_in0;
	wire [0:0] notOp_136_out;
	notOp #(.WIDTH(1)) notOp_136(.in(notOp_136_in0), .out(notOp_136_out));

	reg [0:0] andOp_137_in0;
	reg [0:0] andOp_137_in1;
	wire [0:0] andOp_137_out;
	andOp #(.WIDTH(1)) andOp_137(.in0(andOp_137_in0), .in1(andOp_137_in1), .out(andOp_137_out));

	reg [0:0] andOp_138_in0;
	reg [0:0] andOp_138_in1;
	wire [0:0] andOp_138_out;
	andOp #(.WIDTH(1)) andOp_138(.in0(andOp_138_in0), .in1(andOp_138_in1), .out(andOp_138_out));

	reg [0:0] andOp_139_in0;
	reg [0:0] andOp_139_in1;
	wire [0:0] andOp_139_out;
	andOp #(.WIDTH(1)) andOp_139(.in0(andOp_139_in0), .in1(andOp_139_in1), .out(andOp_139_out));

	reg [0:0] br_1_happened_in_state_4_in_data;
	wire [0:0] br_1_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened_in_state_4(.in_data(br_1_happened_in_state_4_in_data), .out_data(br_1_happened_in_state_4_out_data));

	reg [0:0] notOp_140_in0;
	wire [0:0] notOp_140_out;
	notOp #(.WIDTH(1)) notOp_140(.in(notOp_140_in0), .out(notOp_140_out));

	reg [31:0] eq_141_in0;
	reg [31:0] eq_141_in1;
	wire [0:0] eq_141_out;
	eq #(.WIDTH(32)) eq_141(.in0(eq_141_in0), .in1(eq_141_in1), .out(eq_141_out));

	reg [31:0] eq_142_in0;
	reg [31:0] eq_142_in1;
	wire [0:0] eq_142_out;
	eq #(.WIDTH(32)) eq_142(.in0(eq_142_in0), .in1(eq_142_in1), .out(eq_142_out));

	reg [0:0] orOp_143_in0;
	reg [0:0] orOp_143_in1;
	wire [0:0] orOp_143_out;
	orOp #(.WIDTH(1)) orOp_143(.in0(orOp_143_in0), .in1(orOp_143_in1), .out(orOp_143_out));

	reg [31:0] eq_144_in0;
	reg [31:0] eq_144_in1;
	wire [0:0] eq_144_out;
	eq #(.WIDTH(32)) eq_144(.in0(eq_144_in0), .in1(eq_144_in1), .out(eq_144_out));

	reg [31:0] eq_145_in0;
	reg [31:0] eq_145_in1;
	wire [0:0] eq_145_out;
	eq #(.WIDTH(32)) eq_145(.in0(eq_145_in0), .in1(eq_145_in1), .out(eq_145_out));

	reg [0:0] orOp_146_in0;
	reg [0:0] orOp_146_in1;
	wire [0:0] orOp_146_out;
	orOp #(.WIDTH(1)) orOp_146(.in0(orOp_146_in0), .in1(orOp_146_in1), .out(orOp_146_out));

	reg [31:0] eq_147_in0;
	reg [31:0] eq_147_in1;
	wire [0:0] eq_147_out;
	eq #(.WIDTH(32)) eq_147(.in0(eq_147_in0), .in1(eq_147_in1), .out(eq_147_out));

	reg [0:0] orOp_148_in0;
	reg [0:0] orOp_148_in1;
	wire [0:0] orOp_148_out;
	orOp #(.WIDTH(1)) orOp_148(.in0(orOp_148_in0), .in1(orOp_148_in1), .out(orOp_148_out));

	reg [31:0] eq_149_in0;
	reg [31:0] eq_149_in1;
	wire [0:0] eq_149_out;
	eq #(.WIDTH(32)) eq_149(.in0(eq_149_in0), .in1(eq_149_in1), .out(eq_149_out));

	reg [31:0] eq_150_in0;
	reg [31:0] eq_150_in1;
	wire [0:0] eq_150_out;
	eq #(.WIDTH(32)) eq_150(.in0(eq_150_in0), .in1(eq_150_in1), .out(eq_150_out));

	reg [0:0] orOp_151_in0;
	reg [0:0] orOp_151_in1;
	wire [0:0] orOp_151_out;
	orOp #(.WIDTH(1)) orOp_151(.in0(orOp_151_in0), .in1(orOp_151_in1), .out(orOp_151_out));

	reg [31:0] eq_152_in0;
	reg [31:0] eq_152_in1;
	wire [0:0] eq_152_out;
	eq #(.WIDTH(32)) eq_152(.in0(eq_152_in0), .in1(eq_152_in1), .out(eq_152_out));

	reg [31:0] eq_153_in0;
	reg [31:0] eq_153_in1;
	wire [0:0] eq_153_out;
	eq #(.WIDTH(32)) eq_153(.in0(eq_153_in0), .in1(eq_153_in1), .out(eq_153_out));

	reg [0:0] orOp_154_in0;
	reg [0:0] orOp_154_in1;
	wire [0:0] orOp_154_out;
	orOp #(.WIDTH(1)) orOp_154(.in0(orOp_154_in0), .in1(orOp_154_in1), .out(orOp_154_out));

	reg [31:0] eq_155_in0;
	reg [31:0] eq_155_in1;
	wire [0:0] eq_155_out;
	eq #(.WIDTH(32)) eq_155(.in0(eq_155_in0), .in1(eq_155_in1), .out(eq_155_out));

	reg [0:0] orOp_156_in0;
	reg [0:0] orOp_156_in1;
	wire [0:0] orOp_156_out;
	orOp #(.WIDTH(1)) orOp_156(.in0(orOp_156_in0), .in1(orOp_156_in1), .out(orOp_156_out));

	reg [31:0] eq_157_in0;
	reg [31:0] eq_157_in1;
	wire [0:0] eq_157_out;
	eq #(.WIDTH(32)) eq_157(.in0(eq_157_in0), .in1(eq_157_in1), .out(eq_157_out));

	reg [0:0] orOp_158_in0;
	reg [0:0] orOp_158_in1;
	wire [0:0] orOp_158_out;
	orOp #(.WIDTH(1)) orOp_158(.in0(orOp_158_in0), .in1(orOp_158_in1), .out(orOp_158_out));

	reg [31:0] eq_159_in0;
	reg [31:0] eq_159_in1;
	wire [0:0] eq_159_out;
	eq #(.WIDTH(32)) eq_159(.in0(eq_159_in0), .in1(eq_159_in1), .out(eq_159_out));

	reg [31:0] eq_160_in0;
	reg [31:0] eq_160_in1;
	wire [0:0] eq_160_out;
	eq #(.WIDTH(32)) eq_160(.in0(eq_160_in0), .in1(eq_160_in1), .out(eq_160_out));

	reg [0:0] orOp_161_in0;
	reg [0:0] orOp_161_in1;
	wire [0:0] orOp_161_out;
	orOp #(.WIDTH(1)) orOp_161(.in0(orOp_161_in0), .in1(orOp_161_in1), .out(orOp_161_out));

	reg [31:0] eq_162_in0;
	reg [31:0] eq_162_in1;
	wire [0:0] eq_162_out;
	eq #(.WIDTH(32)) eq_162(.in0(eq_162_in0), .in1(eq_162_in1), .out(eq_162_out));

	reg [0:0] orOp_163_in0;
	reg [0:0] orOp_163_in1;
	wire [0:0] orOp_163_out;
	orOp #(.WIDTH(1)) orOp_163(.in0(orOp_163_in0), .in1(orOp_163_in1), .out(orOp_163_out));

	reg [31:0] eq_164_in0;
	reg [31:0] eq_164_in1;
	wire [0:0] eq_164_out;
	eq #(.WIDTH(32)) eq_164(.in0(eq_164_in0), .in1(eq_164_in1), .out(eq_164_out));

	reg [31:0] eq_165_in0;
	reg [31:0] eq_165_in1;
	wire [0:0] eq_165_out;
	eq #(.WIDTH(32)) eq_165(.in0(eq_165_in0), .in1(eq_165_in1), .out(eq_165_out));

	reg [0:0] notOp_166_in0;
	wire [0:0] notOp_166_out;
	notOp #(.WIDTH(1)) notOp_166(.in(notOp_166_in0), .out(notOp_166_out));

	reg [0:0] andOp_167_in0;
	reg [0:0] andOp_167_in1;
	wire [0:0] andOp_167_out;
	andOp #(.WIDTH(1)) andOp_167(.in0(andOp_167_in0), .in1(andOp_167_in1), .out(andOp_167_out));

	reg [31:0] eq_168_in0;
	reg [31:0] eq_168_in1;
	wire [0:0] eq_168_out;
	eq #(.WIDTH(32)) eq_168(.in0(eq_168_in0), .in1(eq_168_in1), .out(eq_168_out));

	reg [31:0] eq_169_in0;
	reg [31:0] eq_169_in1;
	wire [0:0] eq_169_out;
	eq #(.WIDTH(32)) eq_169(.in0(eq_169_in0), .in1(eq_169_in1), .out(eq_169_out));

	reg [0:0] notOp_170_in0;
	wire [0:0] notOp_170_out;
	notOp #(.WIDTH(1)) notOp_170(.in(notOp_170_in0), .out(notOp_170_out));

	reg [0:0] andOp_171_in0;
	reg [0:0] andOp_171_in1;
	wire [0:0] andOp_171_out;
	andOp #(.WIDTH(1)) andOp_171(.in0(andOp_171_in0), .in1(andOp_171_in1), .out(andOp_171_out));

	reg [31:0] eq_172_in0;
	reg [31:0] eq_172_in1;
	wire [0:0] eq_172_out;
	eq #(.WIDTH(32)) eq_172(.in0(eq_172_in0), .in1(eq_172_in1), .out(eq_172_out));

	reg [0:0] notOp_173_in0;
	wire [0:0] notOp_173_out;
	notOp #(.WIDTH(1)) notOp_173(.in(notOp_173_in0), .out(notOp_173_out));

	reg [0:0] andOp_174_in0;
	reg [0:0] andOp_174_in1;
	wire [0:0] andOp_174_out;
	andOp #(.WIDTH(1)) andOp_174(.in0(andOp_174_in0), .in1(andOp_174_in1), .out(andOp_174_out));

	reg [31:0] eq_175_in0;
	reg [31:0] eq_175_in1;
	wire [0:0] eq_175_out;
	eq #(.WIDTH(32)) eq_175(.in0(eq_175_in0), .in1(eq_175_in1), .out(eq_175_out));

	reg [31:0] eq_176_in0;
	reg [31:0] eq_176_in1;
	wire [0:0] eq_176_out;
	eq #(.WIDTH(32)) eq_176(.in0(eq_176_in0), .in1(eq_176_in1), .out(eq_176_out));

	reg [0:0] notOp_177_in0;
	wire [0:0] notOp_177_out;
	notOp #(.WIDTH(1)) notOp_177(.in(notOp_177_in0), .out(notOp_177_out));

	reg [0:0] andOp_178_in0;
	reg [0:0] andOp_178_in1;
	wire [0:0] andOp_178_out;
	andOp #(.WIDTH(1)) andOp_178(.in0(andOp_178_in0), .in1(andOp_178_in1), .out(andOp_178_out));

	reg [31:0] eq_179_in0;
	reg [31:0] eq_179_in1;
	wire [0:0] eq_179_out;
	eq #(.WIDTH(32)) eq_179(.in0(eq_179_in0), .in1(eq_179_in1), .out(eq_179_out));

	reg [31:0] eq_180_in0;
	reg [31:0] eq_180_in1;
	wire [0:0] eq_180_out;
	eq #(.WIDTH(32)) eq_180(.in0(eq_180_in0), .in1(eq_180_in1), .out(eq_180_out));

	reg [0:0] notOp_181_in0;
	wire [0:0] notOp_181_out;
	notOp #(.WIDTH(1)) notOp_181(.in(notOp_181_in0), .out(notOp_181_out));

	reg [0:0] andOp_182_in0;
	reg [0:0] andOp_182_in1;
	wire [0:0] andOp_182_out;
	andOp #(.WIDTH(1)) andOp_182(.in0(andOp_182_in0), .in1(andOp_182_in1), .out(andOp_182_out));

	reg [31:0] eq_183_in0;
	reg [31:0] eq_183_in1;
	wire [0:0] eq_183_out;
	eq #(.WIDTH(32)) eq_183(.in0(eq_183_in0), .in1(eq_183_in1), .out(eq_183_out));

	reg [0:0] notOp_184_in0;
	wire [0:0] notOp_184_out;
	notOp #(.WIDTH(1)) notOp_184(.in(notOp_184_in0), .out(notOp_184_out));

	reg [0:0] andOp_185_in0;
	reg [0:0] andOp_185_in1;
	wire [0:0] andOp_185_out;
	andOp #(.WIDTH(1)) andOp_185(.in0(andOp_185_in0), .in1(andOp_185_in1), .out(andOp_185_out));

	reg [31:0] eq_186_in0;
	reg [31:0] eq_186_in1;
	wire [0:0] eq_186_out;
	eq #(.WIDTH(32)) eq_186(.in0(eq_186_in0), .in1(eq_186_in1), .out(eq_186_out));

	reg [0:0] notOp_187_in0;
	wire [0:0] notOp_187_out;
	notOp #(.WIDTH(1)) notOp_187(.in(notOp_187_in0), .out(notOp_187_out));

	reg [0:0] andOp_188_in0;
	reg [0:0] andOp_188_in1;
	wire [0:0] andOp_188_out;
	andOp #(.WIDTH(1)) andOp_188(.in0(andOp_188_in0), .in1(andOp_188_in1), .out(andOp_188_out));

	reg [31:0] eq_189_in0;
	reg [31:0] eq_189_in1;
	wire [0:0] eq_189_out;
	eq #(.WIDTH(32)) eq_189(.in0(eq_189_in0), .in1(eq_189_in1), .out(eq_189_out));

	reg [31:0] eq_190_in0;
	reg [31:0] eq_190_in1;
	wire [0:0] eq_190_out;
	eq #(.WIDTH(32)) eq_190(.in0(eq_190_in0), .in1(eq_190_in1), .out(eq_190_out));

	reg [0:0] notOp_191_in0;
	wire [0:0] notOp_191_out;
	notOp #(.WIDTH(1)) notOp_191(.in(notOp_191_in0), .out(notOp_191_out));

	reg [0:0] andOp_192_in0;
	reg [0:0] andOp_192_in1;
	wire [0:0] andOp_192_out;
	andOp #(.WIDTH(1)) andOp_192(.in0(andOp_192_in0), .in1(andOp_192_in1), .out(andOp_192_out));

	reg [31:0] eq_193_in0;
	reg [31:0] eq_193_in1;
	wire [0:0] eq_193_out;
	eq #(.WIDTH(32)) eq_193(.in0(eq_193_in0), .in1(eq_193_in1), .out(eq_193_out));

	reg [0:0] notOp_194_in0;
	wire [0:0] notOp_194_out;
	notOp #(.WIDTH(1)) notOp_194(.in(notOp_194_in0), .out(notOp_194_out));

	reg [0:0] andOp_195_in0;
	reg [0:0] andOp_195_in1;
	wire [0:0] andOp_195_out;
	andOp #(.WIDTH(1)) andOp_195(.in0(andOp_195_in0), .in1(andOp_195_in1), .out(andOp_195_out));

	reg [0:0] andOp_196_in0;
	reg [0:0] andOp_196_in1;
	wire [0:0] andOp_196_out;
	andOp #(.WIDTH(1)) andOp_196(.in0(andOp_196_in0), .in1(andOp_196_in1), .out(andOp_196_out));

	reg [0:0] andOp_197_in0;
	reg [0:0] andOp_197_in1;
	wire [0:0] andOp_197_out;
	andOp #(.WIDTH(1)) andOp_197(.in0(andOp_197_in0), .in1(andOp_197_in1), .out(andOp_197_out));

	reg [0:0] andOp_198_in0;
	reg [0:0] andOp_198_in1;
	wire [0:0] andOp_198_out;
	andOp #(.WIDTH(1)) andOp_198(.in0(andOp_198_in0), .in1(andOp_198_in1), .out(andOp_198_out));

	reg [0:0] andOp_199_in0;
	reg [0:0] andOp_199_in1;
	wire [0:0] andOp_199_out;
	andOp #(.WIDTH(1)) andOp_199(.in0(andOp_199_in0), .in1(andOp_199_in1), .out(andOp_199_out));

	reg [0:0] andOp_200_in0;
	reg [0:0] andOp_200_in1;
	wire [0:0] andOp_200_out;
	andOp #(.WIDTH(1)) andOp_200(.in0(andOp_200_in0), .in1(andOp_200_in1), .out(andOp_200_out));

	reg [0:0] andOp_201_in0;
	reg [0:0] andOp_201_in1;
	wire [0:0] andOp_201_out;
	andOp #(.WIDTH(1)) andOp_201(.in0(andOp_201_in0), .in1(andOp_201_in1), .out(andOp_201_out));

	reg [0:0] andOp_202_in0;
	reg [0:0] andOp_202_in1;
	wire [0:0] andOp_202_out;
	andOp #(.WIDTH(1)) andOp_202(.in0(andOp_202_in0), .in1(andOp_202_in1), .out(andOp_202_out));

	reg [0:0] andOp_203_in0;
	reg [0:0] andOp_203_in1;
	wire [0:0] andOp_203_out;
	andOp #(.WIDTH(1)) andOp_203(.in0(andOp_203_in0), .in1(andOp_203_in1), .out(andOp_203_out));

	reg [0:0] andOp_204_in0;
	reg [0:0] andOp_204_in1;
	wire [0:0] andOp_204_out;
	andOp #(.WIDTH(1)) andOp_204(.in0(andOp_204_in0), .in1(andOp_204_in1), .out(andOp_204_out));

	reg [0:0] andOp_205_in0;
	reg [0:0] andOp_205_in1;
	wire [0:0] andOp_205_out;
	andOp #(.WIDTH(1)) andOp_205(.in0(andOp_205_in0), .in1(andOp_205_in1), .out(andOp_205_out));

	reg [0:0] andOp_206_in0;
	reg [0:0] andOp_206_in1;
	wire [0:0] andOp_206_out;
	andOp #(.WIDTH(1)) andOp_206(.in0(andOp_206_in0), .in1(andOp_206_in1), .out(andOp_206_out));

	reg [31:0] concat_207_in0;
	reg [31:0] concat_207_in1;
	wire [63:0] concat_207_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_207(.in0(concat_207_in0), .in1(concat_207_in1), .out(concat_207_out));

	reg [31:0] concat_208_in0;
	reg [31:0] concat_208_in1;
	wire [63:0] concat_208_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_208(.in0(concat_208_in0), .in1(concat_208_in1), .out(concat_208_out));

	reg [0:0] andOp_209_in0;
	reg [0:0] andOp_209_in1;
	wire [0:0] andOp_209_out;
	andOp #(.WIDTH(1)) andOp_209(.in0(andOp_209_in0), .in1(andOp_209_in1), .out(andOp_209_out));

	reg [31:0] tmp_output_210_in_data;
	wire [31:0] tmp_output_210_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_210(.in_data(tmp_output_210_in_data), .out_data(tmp_output_210_out_data));

	reg [31:0] eq_211_in0;
	reg [31:0] eq_211_in1;
	wire [0:0] eq_211_out;
	eq #(.WIDTH(32)) eq_211(.in0(eq_211_in0), .in1(eq_211_in1), .out(eq_211_out));

	reg [0:0] andOp_212_in0;
	reg [0:0] andOp_212_in1;
	wire [0:0] andOp_212_out;
	andOp #(.WIDTH(1)) andOp_212(.in0(andOp_212_in0), .in1(andOp_212_in1), .out(andOp_212_out));

	reg [0:0] andOp_213_in0;
	reg [0:0] andOp_213_in1;
	wire [0:0] andOp_213_out;
	andOp #(.WIDTH(1)) andOp_213(.in0(andOp_213_in0), .in1(andOp_213_in1), .out(andOp_213_out));

	reg [0:0] andOp_214_in0;
	reg [0:0] andOp_214_in1;
	wire [0:0] andOp_214_out;
	andOp #(.WIDTH(1)) andOp_214(.in0(andOp_214_in0), .in1(andOp_214_in1), .out(andOp_214_out));

	reg [0:0] andOp_215_in0;
	reg [0:0] andOp_215_in1;
	wire [0:0] andOp_215_out;
	andOp #(.WIDTH(1)) andOp_215(.in0(andOp_215_in0), .in1(andOp_215_in1), .out(andOp_215_out));

	reg [0:0] andOp_216_in0;
	reg [0:0] andOp_216_in1;
	wire [0:0] andOp_216_out;
	andOp #(.WIDTH(1)) andOp_216(.in0(andOp_216_in0), .in1(andOp_216_in1), .out(andOp_216_out));

	reg [0:0] andOp_217_in0;
	reg [0:0] andOp_217_in1;
	wire [0:0] andOp_217_out;
	andOp #(.WIDTH(1)) andOp_217(.in0(andOp_217_in0), .in1(andOp_217_in1), .out(andOp_217_out));

	reg [0:0] andOp_218_in0;
	reg [0:0] andOp_218_in1;
	wire [0:0] andOp_218_out;
	andOp #(.WIDTH(1)) andOp_218(.in0(andOp_218_in0), .in1(andOp_218_in1), .out(andOp_218_out));

	reg [0:0] andOp_219_in0;
	reg [0:0] andOp_219_in1;
	wire [0:0] andOp_219_out;
	andOp #(.WIDTH(1)) andOp_219(.in0(andOp_219_in0), .in1(andOp_219_in1), .out(andOp_219_out));

	reg [0:0] andOp_220_in0;
	reg [0:0] andOp_220_in1;
	wire [0:0] andOp_220_out;
	andOp #(.WIDTH(1)) andOp_220(.in0(andOp_220_in0), .in1(andOp_220_in1), .out(andOp_220_out));

	reg [0:0] andOp_221_in0;
	reg [0:0] andOp_221_in1;
	wire [0:0] andOp_221_out;
	andOp #(.WIDTH(1)) andOp_221(.in0(andOp_221_in0), .in1(andOp_221_in1), .out(andOp_221_out));

	reg [0:0] andOp_222_in0;
	reg [0:0] andOp_222_in1;
	wire [0:0] andOp_222_out;
	andOp #(.WIDTH(1)) andOp_222(.in0(andOp_222_in0), .in1(andOp_222_in1), .out(andOp_222_out));

	reg [0:0] notOp_223_in0;
	wire [0:0] notOp_223_out;
	notOp #(.WIDTH(1)) notOp_223(.in(notOp_223_in0), .out(notOp_223_out));

	reg [0:0] andOp_224_in0;
	reg [0:0] andOp_224_in1;
	wire [0:0] andOp_224_out;
	andOp #(.WIDTH(1)) andOp_224(.in0(andOp_224_in0), .in1(andOp_224_in1), .out(andOp_224_out));

	reg [0:0] notOp_225_in0;
	wire [0:0] notOp_225_out;
	notOp #(.WIDTH(1)) notOp_225(.in(notOp_225_in0), .out(notOp_225_out));

	reg [0:0] andOp_226_in0;
	reg [0:0] andOp_226_in1;
	wire [0:0] andOp_226_out;
	andOp #(.WIDTH(1)) andOp_226(.in0(andOp_226_in0), .in1(andOp_226_in1), .out(andOp_226_out));

	reg [0:0] notOp_227_in0;
	wire [0:0] notOp_227_out;
	notOp #(.WIDTH(1)) notOp_227(.in(notOp_227_in0), .out(notOp_227_out));

	reg [0:0] andOp_228_in0;
	reg [0:0] andOp_228_in1;
	wire [0:0] andOp_228_out;
	andOp #(.WIDTH(1)) andOp_228(.in0(andOp_228_in0), .in1(andOp_228_in1), .out(andOp_228_out));

	reg [0:0] notOp_229_in0;
	wire [0:0] notOp_229_out;
	notOp #(.WIDTH(1)) notOp_229(.in(notOp_229_in0), .out(notOp_229_out));

	reg [0:0] andOp_230_in0;
	reg [0:0] andOp_230_in1;
	wire [0:0] andOp_230_out;
	andOp #(.WIDTH(1)) andOp_230(.in0(andOp_230_in0), .in1(andOp_230_in1), .out(andOp_230_out));

	reg [0:0] notOp_231_in0;
	wire [0:0] notOp_231_out;
	notOp #(.WIDTH(1)) notOp_231(.in(notOp_231_in0), .out(notOp_231_out));

	reg [0:0] andOp_232_in0;
	reg [0:0] andOp_232_in1;
	wire [0:0] andOp_232_out;
	andOp #(.WIDTH(1)) andOp_232(.in0(andOp_232_in0), .in1(andOp_232_in1), .out(andOp_232_out));

	reg [0:0] notOp_233_in0;
	wire [0:0] notOp_233_out;
	notOp #(.WIDTH(1)) notOp_233(.in(notOp_233_in0), .out(notOp_233_out));

	reg [0:0] andOp_234_in0;
	reg [0:0] andOp_234_in1;
	wire [0:0] andOp_234_out;
	andOp #(.WIDTH(1)) andOp_234(.in0(andOp_234_in0), .in1(andOp_234_in1), .out(andOp_234_out));

	reg [0:0] notOp_235_in0;
	wire [0:0] notOp_235_out;
	notOp #(.WIDTH(1)) notOp_235(.in(notOp_235_in0), .out(notOp_235_out));

	reg [0:0] andOp_236_in0;
	reg [0:0] andOp_236_in1;
	wire [0:0] andOp_236_out;
	andOp #(.WIDTH(1)) andOp_236(.in0(andOp_236_in0), .in1(andOp_236_in1), .out(andOp_236_out));

	reg [0:0] notOp_237_in0;
	wire [0:0] notOp_237_out;
	notOp #(.WIDTH(1)) notOp_237(.in(notOp_237_in0), .out(notOp_237_out));

	reg [0:0] andOp_238_in0;
	reg [0:0] andOp_238_in1;
	wire [0:0] andOp_238_out;
	andOp #(.WIDTH(1)) andOp_238(.in0(andOp_238_in0), .in1(andOp_238_in1), .out(andOp_238_out));

	reg [0:0] andOp_239_in0;
	reg [0:0] andOp_239_in1;
	wire [0:0] andOp_239_out;
	andOp #(.WIDTH(1)) andOp_239(.in0(andOp_239_in0), .in1(andOp_239_in1), .out(andOp_239_out));

	reg [0:0] andOp_240_in0;
	reg [0:0] andOp_240_in1;
	wire [0:0] andOp_240_out;
	andOp #(.WIDTH(1)) andOp_240(.in0(andOp_240_in0), .in1(andOp_240_in1), .out(andOp_240_out));

	reg [0:0] andOp_241_in0;
	reg [0:0] andOp_241_in1;
	wire [0:0] andOp_241_out;
	andOp #(.WIDTH(1)) andOp_241(.in0(andOp_241_in0), .in1(andOp_241_in1), .out(andOp_241_out));

	reg [0:0] andOp_242_in0;
	reg [0:0] andOp_242_in1;
	wire [0:0] andOp_242_out;
	andOp #(.WIDTH(1)) andOp_242(.in0(andOp_242_in0), .in1(andOp_242_in1), .out(andOp_242_out));

	reg [31:0] eq_243_in0;
	reg [31:0] eq_243_in1;
	wire [0:0] eq_243_out;
	eq #(.WIDTH(32)) eq_243(.in0(eq_243_in0), .in1(eq_243_in1), .out(eq_243_out));

	reg [0:0] andOp_244_in0;
	reg [0:0] andOp_244_in1;
	wire [0:0] andOp_244_out;
	andOp #(.WIDTH(1)) andOp_244(.in0(andOp_244_in0), .in1(andOp_244_in1), .out(andOp_244_out));

	reg [31:0] eq_245_in0;
	reg [31:0] eq_245_in1;
	wire [0:0] eq_245_out;
	eq #(.WIDTH(32)) eq_245(.in0(eq_245_in0), .in1(eq_245_in1), .out(eq_245_out));

	reg [0:0] andOp_246_in0;
	reg [0:0] andOp_246_in1;
	wire [0:0] andOp_246_out;
	andOp #(.WIDTH(1)) andOp_246(.in0(andOp_246_in0), .in1(andOp_246_in1), .out(andOp_246_out));

	reg [31:0] eq_247_in0;
	reg [31:0] eq_247_in1;
	wire [0:0] eq_247_out;
	eq #(.WIDTH(32)) eq_247(.in0(eq_247_in0), .in1(eq_247_in1), .out(eq_247_out));

	reg [0:0] andOp_248_in0;
	reg [0:0] andOp_248_in1;
	wire [0:0] andOp_248_out;
	andOp #(.WIDTH(1)) andOp_248(.in0(andOp_248_in0), .in1(andOp_248_in1), .out(andOp_248_out));

	reg [31:0] eq_249_in0;
	reg [31:0] eq_249_in1;
	wire [0:0] eq_249_out;
	eq #(.WIDTH(32)) eq_249(.in0(eq_249_in0), .in1(eq_249_in1), .out(eq_249_out));

	reg [0:0] andOp_250_in0;
	reg [0:0] andOp_250_in1;
	wire [0:0] andOp_250_out;
	andOp #(.WIDTH(1)) andOp_250(.in0(andOp_250_in0), .in1(andOp_250_in1), .out(andOp_250_out));

	reg [31:0] eq_251_in0;
	reg [31:0] eq_251_in1;
	wire [0:0] eq_251_out;
	eq #(.WIDTH(32)) eq_251(.in0(eq_251_in0), .in1(eq_251_in1), .out(eq_251_out));

	reg [0:0] andOp_252_in0;
	reg [0:0] andOp_252_in1;
	wire [0:0] andOp_252_out;
	andOp #(.WIDTH(1)) andOp_252(.in0(andOp_252_in0), .in1(andOp_252_in1), .out(andOp_252_out));

	reg [0:0] andOp_253_in0;
	reg [0:0] andOp_253_in1;
	wire [0:0] andOp_253_out;
	andOp #(.WIDTH(1)) andOp_253(.in0(andOp_253_in0), .in1(andOp_253_in1), .out(andOp_253_out));

	reg [31:0] eq_254_in0;
	reg [31:0] eq_254_in1;
	wire [0:0] eq_254_out;
	eq #(.WIDTH(32)) eq_254(.in0(eq_254_in0), .in1(eq_254_in1), .out(eq_254_out));

	reg [0:0] andOp_255_in0;
	reg [0:0] andOp_255_in1;
	wire [0:0] andOp_255_out;
	andOp #(.WIDTH(1)) andOp_255(.in0(andOp_255_in0), .in1(andOp_255_in1), .out(andOp_255_out));

	reg [0:0] notOp_256_in0;
	wire [0:0] notOp_256_out;
	notOp #(.WIDTH(1)) notOp_256(.in(notOp_256_in0), .out(notOp_256_out));

	reg [0:0] andOp_257_in0;
	reg [0:0] andOp_257_in1;
	wire [0:0] andOp_257_out;
	andOp #(.WIDTH(1)) andOp_257(.in0(andOp_257_in0), .in1(andOp_257_in1), .out(andOp_257_out));

	reg [0:0] notOp_258_in0;
	wire [0:0] notOp_258_out;
	notOp #(.WIDTH(1)) notOp_258(.in(notOp_258_in0), .out(notOp_258_out));

	reg [0:0] andOp_259_in0;
	reg [0:0] andOp_259_in1;
	wire [0:0] andOp_259_out;
	andOp #(.WIDTH(1)) andOp_259(.in0(andOp_259_in0), .in1(andOp_259_in1), .out(andOp_259_out));

	reg [0:0] notOp_260_in0;
	wire [0:0] notOp_260_out;
	notOp #(.WIDTH(1)) notOp_260(.in(notOp_260_in0), .out(notOp_260_out));

	reg [0:0] andOp_261_in0;
	reg [0:0] andOp_261_in1;
	wire [0:0] andOp_261_out;
	andOp #(.WIDTH(1)) andOp_261(.in0(andOp_261_in0), .in1(andOp_261_in1), .out(andOp_261_out));

	reg [0:0] andOp_262_in0;
	reg [0:0] andOp_262_in1;
	wire [0:0] andOp_262_out;
	andOp #(.WIDTH(1)) andOp_262(.in0(andOp_262_in0), .in1(andOp_262_in1), .out(andOp_262_out));

	reg [31:0] eq_263_in0;
	reg [31:0] eq_263_in1;
	wire [0:0] eq_263_out;
	eq #(.WIDTH(32)) eq_263(.in0(eq_263_in0), .in1(eq_263_in1), .out(eq_263_out));

	reg [0:0] andOp_264_in0;
	reg [0:0] andOp_264_in1;
	wire [0:0] andOp_264_out;
	andOp #(.WIDTH(1)) andOp_264(.in0(andOp_264_in0), .in1(andOp_264_in1), .out(andOp_264_out));

	reg [0:0] notOp_265_in0;
	wire [0:0] notOp_265_out;
	notOp #(.WIDTH(1)) notOp_265(.in(notOp_265_in0), .out(notOp_265_out));

	reg [0:0] andOp_266_in0;
	reg [0:0] andOp_266_in1;
	wire [0:0] andOp_266_out;
	andOp #(.WIDTH(1)) andOp_266(.in0(andOp_266_in0), .in1(andOp_266_in1), .out(andOp_266_out));

	reg [0:0] notOp_267_in0;
	wire [0:0] notOp_267_out;
	notOp #(.WIDTH(1)) notOp_267(.in(notOp_267_in0), .out(notOp_267_out));

	reg [0:0] andOp_268_in0;
	reg [0:0] andOp_268_in1;
	wire [0:0] andOp_268_out;
	andOp #(.WIDTH(1)) andOp_268(.in0(andOp_268_in0), .in1(andOp_268_in1), .out(andOp_268_out));

	reg [0:0] notOp_269_in0;
	wire [0:0] notOp_269_out;
	notOp #(.WIDTH(1)) notOp_269(.in(notOp_269_in0), .out(notOp_269_out));

	reg [0:0] andOp_270_in0;
	reg [0:0] andOp_270_in1;
	wire [0:0] andOp_270_out;
	andOp #(.WIDTH(1)) andOp_270(.in0(andOp_270_in0), .in1(andOp_270_in1), .out(andOp_270_out));

	reg [0:0] andOp_271_in0;
	reg [0:0] andOp_271_in1;
	wire [0:0] andOp_271_out;
	andOp #(.WIDTH(1)) andOp_271(.in0(andOp_271_in0), .in1(andOp_271_in1), .out(andOp_271_out));

	reg [31:0] eq_272_in0;
	reg [31:0] eq_272_in1;
	wire [0:0] eq_272_out;
	eq #(.WIDTH(32)) eq_272(.in0(eq_272_in0), .in1(eq_272_in1), .out(eq_272_out));

	reg [0:0] andOp_273_in0;
	reg [0:0] andOp_273_in1;
	wire [0:0] andOp_273_out;
	andOp #(.WIDTH(1)) andOp_273(.in0(andOp_273_in0), .in1(andOp_273_in1), .out(andOp_273_out));

	reg [0:0] notOp_274_in0;
	wire [0:0] notOp_274_out;
	notOp #(.WIDTH(1)) notOp_274(.in(notOp_274_in0), .out(notOp_274_out));

	reg [0:0] andOp_275_in0;
	reg [0:0] andOp_275_in1;
	wire [0:0] andOp_275_out;
	andOp #(.WIDTH(1)) andOp_275(.in0(andOp_275_in0), .in1(andOp_275_in1), .out(andOp_275_out));

	reg [0:0] notOp_276_in0;
	wire [0:0] notOp_276_out;
	notOp #(.WIDTH(1)) notOp_276(.in(notOp_276_in0), .out(notOp_276_out));

	reg [0:0] andOp_277_in0;
	reg [0:0] andOp_277_in1;
	wire [0:0] andOp_277_out;
	andOp #(.WIDTH(1)) andOp_277(.in0(andOp_277_in0), .in1(andOp_277_in1), .out(andOp_277_out));

	reg [0:0] notOp_278_in0;
	wire [0:0] notOp_278_out;
	notOp #(.WIDTH(1)) notOp_278(.in(notOp_278_in0), .out(notOp_278_out));

	reg [0:0] andOp_279_in0;
	reg [0:0] andOp_279_in1;
	wire [0:0] andOp_279_out;
	andOp #(.WIDTH(1)) andOp_279(.in0(andOp_279_in0), .in1(andOp_279_in1), .out(andOp_279_out));

	reg [0:0] andOp_280_in0;
	reg [0:0] andOp_280_in1;
	wire [0:0] andOp_280_out;
	andOp #(.WIDTH(1)) andOp_280(.in0(andOp_280_in0), .in1(andOp_280_in1), .out(andOp_280_out));

	reg [31:0] eq_281_in0;
	reg [31:0] eq_281_in1;
	wire [0:0] eq_281_out;
	eq #(.WIDTH(32)) eq_281(.in0(eq_281_in0), .in1(eq_281_in1), .out(eq_281_out));

	reg [0:0] andOp_282_in0;
	reg [0:0] andOp_282_in1;
	wire [0:0] andOp_282_out;
	andOp #(.WIDTH(1)) andOp_282(.in0(andOp_282_in0), .in1(andOp_282_in1), .out(andOp_282_out));

	reg [0:0] notOp_283_in0;
	wire [0:0] notOp_283_out;
	notOp #(.WIDTH(1)) notOp_283(.in(notOp_283_in0), .out(notOp_283_out));

	reg [0:0] andOp_284_in0;
	reg [0:0] andOp_284_in1;
	wire [0:0] andOp_284_out;
	andOp #(.WIDTH(1)) andOp_284(.in0(andOp_284_in0), .in1(andOp_284_in1), .out(andOp_284_out));

	reg [0:0] notOp_285_in0;
	wire [0:0] notOp_285_out;
	notOp #(.WIDTH(1)) notOp_285(.in(notOp_285_in0), .out(notOp_285_out));

	reg [0:0] andOp_286_in0;
	reg [0:0] andOp_286_in1;
	wire [0:0] andOp_286_out;
	andOp #(.WIDTH(1)) andOp_286(.in0(andOp_286_in0), .in1(andOp_286_in1), .out(andOp_286_out));

	reg [0:0] notOp_287_in0;
	wire [0:0] notOp_287_out;
	notOp #(.WIDTH(1)) notOp_287(.in(notOp_287_in0), .out(notOp_287_out));

	reg [0:0] andOp_288_in0;
	reg [0:0] andOp_288_in1;
	wire [0:0] andOp_288_out;
	andOp #(.WIDTH(1)) andOp_288(.in0(andOp_288_in0), .in1(andOp_288_in1), .out(andOp_288_out));

	reg [0:0] andOp_289_in0;
	reg [0:0] andOp_289_in1;
	wire [0:0] andOp_289_out;
	andOp #(.WIDTH(1)) andOp_289(.in0(andOp_289_in0), .in1(andOp_289_in1), .out(andOp_289_out));

	reg [31:0] eq_290_in0;
	reg [31:0] eq_290_in1;
	wire [0:0] eq_290_out;
	eq #(.WIDTH(32)) eq_290(.in0(eq_290_in0), .in1(eq_290_in1), .out(eq_290_out));

	reg [0:0] andOp_291_in0;
	reg [0:0] andOp_291_in1;
	wire [0:0] andOp_291_out;
	andOp #(.WIDTH(1)) andOp_291(.in0(andOp_291_in0), .in1(andOp_291_in1), .out(andOp_291_out));

	reg [0:0] notOp_292_in0;
	wire [0:0] notOp_292_out;
	notOp #(.WIDTH(1)) notOp_292(.in(notOp_292_in0), .out(notOp_292_out));

	reg [0:0] andOp_293_in0;
	reg [0:0] andOp_293_in1;
	wire [0:0] andOp_293_out;
	andOp #(.WIDTH(1)) andOp_293(.in0(andOp_293_in0), .in1(andOp_293_in1), .out(andOp_293_out));

	reg [0:0] notOp_294_in0;
	wire [0:0] notOp_294_out;
	notOp #(.WIDTH(1)) notOp_294(.in(notOp_294_in0), .out(notOp_294_out));

	reg [0:0] andOp_295_in0;
	reg [0:0] andOp_295_in1;
	wire [0:0] andOp_295_out;
	andOp #(.WIDTH(1)) andOp_295(.in0(andOp_295_in0), .in1(andOp_295_in1), .out(andOp_295_out));

	reg [0:0] notOp_296_in0;
	wire [0:0] notOp_296_out;
	notOp #(.WIDTH(1)) notOp_296(.in(notOp_296_in0), .out(notOp_296_out));

	reg [0:0] andOp_297_in0;
	reg [0:0] andOp_297_in1;
	wire [0:0] andOp_297_out;
	andOp #(.WIDTH(1)) andOp_297(.in0(andOp_297_in0), .in1(andOp_297_in1), .out(andOp_297_out));

	reg [0:0] andOp_298_in0;
	reg [0:0] andOp_298_in1;
	wire [0:0] andOp_298_out;
	andOp #(.WIDTH(1)) andOp_298(.in0(andOp_298_in0), .in1(andOp_298_in1), .out(andOp_298_out));

	reg [31:0] eq_299_in0;
	reg [31:0] eq_299_in1;
	wire [0:0] eq_299_out;
	eq #(.WIDTH(32)) eq_299(.in0(eq_299_in0), .in1(eq_299_in1), .out(eq_299_out));

	reg [0:0] andOp_300_in0;
	reg [0:0] andOp_300_in1;
	wire [0:0] andOp_300_out;
	andOp #(.WIDTH(1)) andOp_300(.in0(andOp_300_in0), .in1(andOp_300_in1), .out(andOp_300_out));

	reg [0:0] notOp_301_in0;
	wire [0:0] notOp_301_out;
	notOp #(.WIDTH(1)) notOp_301(.in(notOp_301_in0), .out(notOp_301_out));

	reg [0:0] andOp_302_in0;
	reg [0:0] andOp_302_in1;
	wire [0:0] andOp_302_out;
	andOp #(.WIDTH(1)) andOp_302(.in0(andOp_302_in0), .in1(andOp_302_in1), .out(andOp_302_out));

	reg [0:0] notOp_303_in0;
	wire [0:0] notOp_303_out;
	notOp #(.WIDTH(1)) notOp_303(.in(notOp_303_in0), .out(notOp_303_out));

	reg [0:0] andOp_304_in0;
	reg [0:0] andOp_304_in1;
	wire [0:0] andOp_304_out;
	andOp #(.WIDTH(1)) andOp_304(.in0(andOp_304_in0), .in1(andOp_304_in1), .out(andOp_304_out));

	reg [0:0] notOp_305_in0;
	wire [0:0] notOp_305_out;
	notOp #(.WIDTH(1)) notOp_305(.in(notOp_305_in0), .out(notOp_305_out));

	reg [0:0] andOp_306_in0;
	reg [0:0] andOp_306_in1;
	wire [0:0] andOp_306_out;
	andOp #(.WIDTH(1)) andOp_306(.in0(andOp_306_in0), .in1(andOp_306_in1), .out(andOp_306_out));

	reg [0:0] andOp_307_in0;
	reg [0:0] andOp_307_in1;
	wire [0:0] andOp_307_out;
	andOp #(.WIDTH(1)) andOp_307(.in0(andOp_307_in0), .in1(andOp_307_in1), .out(andOp_307_out));

	reg [31:0] eq_308_in0;
	reg [31:0] eq_308_in1;
	wire [0:0] eq_308_out;
	eq #(.WIDTH(32)) eq_308(.in0(eq_308_in0), .in1(eq_308_in1), .out(eq_308_out));

	reg [0:0] andOp_309_in0;
	reg [0:0] andOp_309_in1;
	wire [0:0] andOp_309_out;
	andOp #(.WIDTH(1)) andOp_309(.in0(andOp_309_in0), .in1(andOp_309_in1), .out(andOp_309_out));

	reg [0:0] notOp_310_in0;
	wire [0:0] notOp_310_out;
	notOp #(.WIDTH(1)) notOp_310(.in(notOp_310_in0), .out(notOp_310_out));

	reg [0:0] andOp_311_in0;
	reg [0:0] andOp_311_in1;
	wire [0:0] andOp_311_out;
	andOp #(.WIDTH(1)) andOp_311(.in0(andOp_311_in0), .in1(andOp_311_in1), .out(andOp_311_out));

	reg [0:0] notOp_312_in0;
	wire [0:0] notOp_312_out;
	notOp #(.WIDTH(1)) notOp_312(.in(notOp_312_in0), .out(notOp_312_out));

	reg [0:0] andOp_313_in0;
	reg [0:0] andOp_313_in1;
	wire [0:0] andOp_313_out;
	andOp #(.WIDTH(1)) andOp_313(.in0(andOp_313_in0), .in1(andOp_313_in1), .out(andOp_313_out));

	reg [0:0] notOp_314_in0;
	wire [0:0] notOp_314_out;
	notOp #(.WIDTH(1)) notOp_314(.in(notOp_314_in0), .out(notOp_314_out));

	reg [0:0] andOp_315_in0;
	reg [0:0] andOp_315_in1;
	wire [0:0] andOp_315_out;
	andOp #(.WIDTH(1)) andOp_315(.in0(andOp_315_in0), .in1(andOp_315_in1), .out(andOp_315_out));

	reg [0:0] andOp_316_in0;
	reg [0:0] andOp_316_in1;
	wire [0:0] andOp_316_out;
	andOp #(.WIDTH(1)) andOp_316(.in0(andOp_316_in0), .in1(andOp_316_in1), .out(andOp_316_out));

	reg [31:0] eq_317_in0;
	reg [31:0] eq_317_in1;
	wire [0:0] eq_317_out;
	eq #(.WIDTH(32)) eq_317(.in0(eq_317_in0), .in1(eq_317_in1), .out(eq_317_out));

	reg [0:0] andOp_318_in0;
	reg [0:0] andOp_318_in1;
	wire [0:0] andOp_318_out;
	andOp #(.WIDTH(1)) andOp_318(.in0(andOp_318_in0), .in1(andOp_318_in1), .out(andOp_318_out));

	reg [0:0] notOp_319_in0;
	wire [0:0] notOp_319_out;
	notOp #(.WIDTH(1)) notOp_319(.in(notOp_319_in0), .out(notOp_319_out));

	reg [0:0] andOp_320_in0;
	reg [0:0] andOp_320_in1;
	wire [0:0] andOp_320_out;
	andOp #(.WIDTH(1)) andOp_320(.in0(andOp_320_in0), .in1(andOp_320_in1), .out(andOp_320_out));

	reg [0:0] notOp_321_in0;
	wire [0:0] notOp_321_out;
	notOp #(.WIDTH(1)) notOp_321(.in(notOp_321_in0), .out(notOp_321_out));

	reg [0:0] andOp_322_in0;
	reg [0:0] andOp_322_in1;
	wire [0:0] andOp_322_out;
	andOp #(.WIDTH(1)) andOp_322(.in0(andOp_322_in0), .in1(andOp_322_in1), .out(andOp_322_out));

	reg [0:0] notOp_323_in0;
	wire [0:0] notOp_323_out;
	notOp #(.WIDTH(1)) notOp_323(.in(notOp_323_in0), .out(notOp_323_out));

	reg [0:0] andOp_324_in0;
	reg [0:0] andOp_324_in1;
	wire [0:0] andOp_324_out;
	andOp #(.WIDTH(1)) andOp_324(.in0(andOp_324_in0), .in1(andOp_324_in1), .out(andOp_324_out));

	reg [0:0] andOp_325_in0;
	reg [0:0] andOp_325_in1;
	wire [0:0] andOp_325_out;
	andOp #(.WIDTH(1)) andOp_325(.in0(andOp_325_in0), .in1(andOp_325_in1), .out(andOp_325_out));

	reg [31:0] eq_326_in0;
	reg [31:0] eq_326_in1;
	wire [0:0] eq_326_out;
	eq #(.WIDTH(32)) eq_326(.in0(eq_326_in0), .in1(eq_326_in1), .out(eq_326_out));

	reg [0:0] andOp_327_in0;
	reg [0:0] andOp_327_in1;
	wire [0:0] andOp_327_out;
	andOp #(.WIDTH(1)) andOp_327(.in0(andOp_327_in0), .in1(andOp_327_in1), .out(andOp_327_out));

	reg [0:0] notOp_328_in0;
	wire [0:0] notOp_328_out;
	notOp #(.WIDTH(1)) notOp_328(.in(notOp_328_in0), .out(notOp_328_out));

	reg [0:0] andOp_329_in0;
	reg [0:0] andOp_329_in1;
	wire [0:0] andOp_329_out;
	andOp #(.WIDTH(1)) andOp_329(.in0(andOp_329_in0), .in1(andOp_329_in1), .out(andOp_329_out));

	reg [0:0] notOp_330_in0;
	wire [0:0] notOp_330_out;
	notOp #(.WIDTH(1)) notOp_330(.in(notOp_330_in0), .out(notOp_330_out));

	reg [0:0] andOp_331_in0;
	reg [0:0] andOp_331_in1;
	wire [0:0] andOp_331_out;
	andOp #(.WIDTH(1)) andOp_331(.in0(andOp_331_in0), .in1(andOp_331_in1), .out(andOp_331_out));

	reg [0:0] notOp_332_in0;
	wire [0:0] notOp_332_out;
	notOp #(.WIDTH(1)) notOp_332(.in(notOp_332_in0), .out(notOp_332_out));

	reg [0:0] andOp_333_in0;
	reg [0:0] andOp_333_in1;
	wire [0:0] andOp_333_out;
	andOp #(.WIDTH(1)) andOp_333(.in0(andOp_333_in0), .in1(andOp_333_in1), .out(andOp_333_out));

	reg [31:0] eq_334_in0;
	reg [31:0] eq_334_in1;
	wire [0:0] eq_334_out;
	eq #(.WIDTH(32)) eq_334(.in0(eq_334_in0), .in1(eq_334_in1), .out(eq_334_out));

	reg [0:0] andOp_335_in0;
	reg [0:0] andOp_335_in1;
	wire [0:0] andOp_335_out;
	andOp #(.WIDTH(1)) andOp_335(.in0(andOp_335_in0), .in1(andOp_335_in1), .out(andOp_335_out));

	reg [31:0] eq_336_in0;
	reg [31:0] eq_336_in1;
	wire [0:0] eq_336_out;
	eq #(.WIDTH(32)) eq_336(.in0(eq_336_in0), .in1(eq_336_in1), .out(eq_336_out));

	reg [0:0] andOp_337_in0;
	reg [0:0] andOp_337_in1;
	wire [0:0] andOp_337_out;
	andOp #(.WIDTH(1)) andOp_337(.in0(andOp_337_in0), .in1(andOp_337_in1), .out(andOp_337_out));

	reg [31:0] eq_338_in0;
	reg [31:0] eq_338_in1;
	wire [0:0] eq_338_out;
	eq #(.WIDTH(32)) eq_338(.in0(eq_338_in0), .in1(eq_338_in1), .out(eq_338_out));

	reg [0:0] andOp_339_in0;
	reg [0:0] andOp_339_in1;
	wire [0:0] andOp_339_out;
	andOp #(.WIDTH(1)) andOp_339(.in0(andOp_339_in0), .in1(andOp_339_in1), .out(andOp_339_out));

	reg [31:0] eq_340_in0;
	reg [31:0] eq_340_in1;
	wire [0:0] eq_340_out;
	eq #(.WIDTH(32)) eq_340(.in0(eq_340_in0), .in1(eq_340_in1), .out(eq_340_out));

	reg [0:0] andOp_341_in0;
	reg [0:0] andOp_341_in1;
	wire [0:0] andOp_341_out;
	andOp #(.WIDTH(1)) andOp_341(.in0(andOp_341_in0), .in1(andOp_341_in1), .out(andOp_341_out));

	reg [31:0] eq_342_in0;
	reg [31:0] eq_342_in1;
	wire [0:0] eq_342_out;
	eq #(.WIDTH(32)) eq_342(.in0(eq_342_in0), .in1(eq_342_in1), .out(eq_342_out));

	reg [0:0] andOp_343_in0;
	reg [0:0] andOp_343_in1;
	wire [0:0] andOp_343_out;
	andOp #(.WIDTH(1)) andOp_343(.in0(andOp_343_in0), .in1(andOp_343_in1), .out(andOp_343_out));

	reg [0:0] andOp_344_in0;
	reg [0:0] andOp_344_in1;
	wire [0:0] andOp_344_out;
	andOp #(.WIDTH(1)) andOp_344(.in0(andOp_344_in0), .in1(andOp_344_in1), .out(andOp_344_out));

	reg [31:0] eq_345_in0;
	reg [31:0] eq_345_in1;
	wire [0:0] eq_345_out;
	eq #(.WIDTH(32)) eq_345(.in0(eq_345_in0), .in1(eq_345_in1), .out(eq_345_out));

	reg [0:0] andOp_346_in0;
	reg [0:0] andOp_346_in1;
	wire [0:0] andOp_346_out;
	andOp #(.WIDTH(1)) andOp_346(.in0(andOp_346_in0), .in1(andOp_346_in1), .out(andOp_346_out));

	reg [0:0] notOp_347_in0;
	wire [0:0] notOp_347_out;
	notOp #(.WIDTH(1)) notOp_347(.in(notOp_347_in0), .out(notOp_347_out));

	reg [0:0] andOp_348_in0;
	reg [0:0] andOp_348_in1;
	wire [0:0] andOp_348_out;
	andOp #(.WIDTH(1)) andOp_348(.in0(andOp_348_in0), .in1(andOp_348_in1), .out(andOp_348_out));

	reg [0:0] notOp_349_in0;
	wire [0:0] notOp_349_out;
	notOp #(.WIDTH(1)) notOp_349(.in(notOp_349_in0), .out(notOp_349_out));

	reg [0:0] andOp_350_in0;
	reg [0:0] andOp_350_in1;
	wire [0:0] andOp_350_out;
	andOp #(.WIDTH(1)) andOp_350(.in0(andOp_350_in0), .in1(andOp_350_in1), .out(andOp_350_out));

	reg [0:0] notOp_351_in0;
	wire [0:0] notOp_351_out;
	notOp #(.WIDTH(1)) notOp_351(.in(notOp_351_in0), .out(notOp_351_out));

	reg [0:0] andOp_352_in0;
	reg [0:0] andOp_352_in1;
	wire [0:0] andOp_352_out;
	andOp #(.WIDTH(1)) andOp_352(.in0(andOp_352_in0), .in1(andOp_352_in1), .out(andOp_352_out));

	reg [0:0] andOp_353_in0;
	reg [0:0] andOp_353_in1;
	wire [0:0] andOp_353_out;
	andOp #(.WIDTH(1)) andOp_353(.in0(andOp_353_in0), .in1(andOp_353_in1), .out(andOp_353_out));

	reg [31:0] eq_354_in0;
	reg [31:0] eq_354_in1;
	wire [0:0] eq_354_out;
	eq #(.WIDTH(32)) eq_354(.in0(eq_354_in0), .in1(eq_354_in1), .out(eq_354_out));

	reg [0:0] andOp_355_in0;
	reg [0:0] andOp_355_in1;
	wire [0:0] andOp_355_out;
	andOp #(.WIDTH(1)) andOp_355(.in0(andOp_355_in0), .in1(andOp_355_in1), .out(andOp_355_out));

	reg [0:0] notOp_356_in0;
	wire [0:0] notOp_356_out;
	notOp #(.WIDTH(1)) notOp_356(.in(notOp_356_in0), .out(notOp_356_out));

	reg [0:0] andOp_357_in0;
	reg [0:0] andOp_357_in1;
	wire [0:0] andOp_357_out;
	andOp #(.WIDTH(1)) andOp_357(.in0(andOp_357_in0), .in1(andOp_357_in1), .out(andOp_357_out));

	reg [0:0] notOp_358_in0;
	wire [0:0] notOp_358_out;
	notOp #(.WIDTH(1)) notOp_358(.in(notOp_358_in0), .out(notOp_358_out));

	reg [0:0] andOp_359_in0;
	reg [0:0] andOp_359_in1;
	wire [0:0] andOp_359_out;
	andOp #(.WIDTH(1)) andOp_359(.in0(andOp_359_in0), .in1(andOp_359_in1), .out(andOp_359_out));

	reg [0:0] notOp_360_in0;
	wire [0:0] notOp_360_out;
	notOp #(.WIDTH(1)) notOp_360(.in(notOp_360_in0), .out(notOp_360_out));

	reg [0:0] andOp_361_in0;
	reg [0:0] andOp_361_in1;
	wire [0:0] andOp_361_out;
	andOp #(.WIDTH(1)) andOp_361(.in0(andOp_361_in0), .in1(andOp_361_in1), .out(andOp_361_out));

	reg [0:0] andOp_362_in0;
	reg [0:0] andOp_362_in1;
	wire [0:0] andOp_362_out;
	andOp #(.WIDTH(1)) andOp_362(.in0(andOp_362_in0), .in1(andOp_362_in1), .out(andOp_362_out));

	reg [31:0] eq_363_in0;
	reg [31:0] eq_363_in1;
	wire [0:0] eq_363_out;
	eq #(.WIDTH(32)) eq_363(.in0(eq_363_in0), .in1(eq_363_in1), .out(eq_363_out));

	reg [0:0] andOp_364_in0;
	reg [0:0] andOp_364_in1;
	wire [0:0] andOp_364_out;
	andOp #(.WIDTH(1)) andOp_364(.in0(andOp_364_in0), .in1(andOp_364_in1), .out(andOp_364_out));

	reg [0:0] notOp_365_in0;
	wire [0:0] notOp_365_out;
	notOp #(.WIDTH(1)) notOp_365(.in(notOp_365_in0), .out(notOp_365_out));

	reg [0:0] andOp_366_in0;
	reg [0:0] andOp_366_in1;
	wire [0:0] andOp_366_out;
	andOp #(.WIDTH(1)) andOp_366(.in0(andOp_366_in0), .in1(andOp_366_in1), .out(andOp_366_out));

	reg [0:0] notOp_367_in0;
	wire [0:0] notOp_367_out;
	notOp #(.WIDTH(1)) notOp_367(.in(notOp_367_in0), .out(notOp_367_out));

	reg [0:0] andOp_368_in0;
	reg [0:0] andOp_368_in1;
	wire [0:0] andOp_368_out;
	andOp #(.WIDTH(1)) andOp_368(.in0(andOp_368_in0), .in1(andOp_368_in1), .out(andOp_368_out));

	reg [0:0] notOp_369_in0;
	wire [0:0] notOp_369_out;
	notOp #(.WIDTH(1)) notOp_369(.in(notOp_369_in0), .out(notOp_369_out));

	reg [0:0] andOp_370_in0;
	reg [0:0] andOp_370_in1;
	wire [0:0] andOp_370_out;
	andOp #(.WIDTH(1)) andOp_370(.in0(andOp_370_in0), .in1(andOp_370_in1), .out(andOp_370_out));

	reg [0:0] andOp_371_in0;
	reg [0:0] andOp_371_in1;
	wire [0:0] andOp_371_out;
	andOp #(.WIDTH(1)) andOp_371(.in0(andOp_371_in0), .in1(andOp_371_in1), .out(andOp_371_out));

	reg [31:0] eq_372_in0;
	reg [31:0] eq_372_in1;
	wire [0:0] eq_372_out;
	eq #(.WIDTH(32)) eq_372(.in0(eq_372_in0), .in1(eq_372_in1), .out(eq_372_out));

	reg [0:0] andOp_373_in0;
	reg [0:0] andOp_373_in1;
	wire [0:0] andOp_373_out;
	andOp #(.WIDTH(1)) andOp_373(.in0(andOp_373_in0), .in1(andOp_373_in1), .out(andOp_373_out));

	reg [0:0] notOp_374_in0;
	wire [0:0] notOp_374_out;
	notOp #(.WIDTH(1)) notOp_374(.in(notOp_374_in0), .out(notOp_374_out));

	reg [0:0] andOp_375_in0;
	reg [0:0] andOp_375_in1;
	wire [0:0] andOp_375_out;
	andOp #(.WIDTH(1)) andOp_375(.in0(andOp_375_in0), .in1(andOp_375_in1), .out(andOp_375_out));

	reg [0:0] notOp_376_in0;
	wire [0:0] notOp_376_out;
	notOp #(.WIDTH(1)) notOp_376(.in(notOp_376_in0), .out(notOp_376_out));

	reg [0:0] andOp_377_in0;
	reg [0:0] andOp_377_in1;
	wire [0:0] andOp_377_out;
	andOp #(.WIDTH(1)) andOp_377(.in0(andOp_377_in0), .in1(andOp_377_in1), .out(andOp_377_out));

	reg [0:0] notOp_378_in0;
	wire [0:0] notOp_378_out;
	notOp #(.WIDTH(1)) notOp_378(.in(notOp_378_in0), .out(notOp_378_out));

	reg [0:0] andOp_379_in0;
	reg [0:0] andOp_379_in1;
	wire [0:0] andOp_379_out;
	andOp #(.WIDTH(1)) andOp_379(.in0(andOp_379_in0), .in1(andOp_379_in1), .out(andOp_379_out));

	reg [0:0] andOp_380_in0;
	reg [0:0] andOp_380_in1;
	wire [0:0] andOp_380_out;
	andOp #(.WIDTH(1)) andOp_380(.in0(andOp_380_in0), .in1(andOp_380_in1), .out(andOp_380_out));

	reg [31:0] eq_381_in0;
	reg [31:0] eq_381_in1;
	wire [0:0] eq_381_out;
	eq #(.WIDTH(32)) eq_381(.in0(eq_381_in0), .in1(eq_381_in1), .out(eq_381_out));

	reg [0:0] andOp_382_in0;
	reg [0:0] andOp_382_in1;
	wire [0:0] andOp_382_out;
	andOp #(.WIDTH(1)) andOp_382(.in0(andOp_382_in0), .in1(andOp_382_in1), .out(andOp_382_out));

	reg [0:0] notOp_383_in0;
	wire [0:0] notOp_383_out;
	notOp #(.WIDTH(1)) notOp_383(.in(notOp_383_in0), .out(notOp_383_out));

	reg [0:0] andOp_384_in0;
	reg [0:0] andOp_384_in1;
	wire [0:0] andOp_384_out;
	andOp #(.WIDTH(1)) andOp_384(.in0(andOp_384_in0), .in1(andOp_384_in1), .out(andOp_384_out));

	reg [0:0] notOp_385_in0;
	wire [0:0] notOp_385_out;
	notOp #(.WIDTH(1)) notOp_385(.in(notOp_385_in0), .out(notOp_385_out));

	reg [0:0] andOp_386_in0;
	reg [0:0] andOp_386_in1;
	wire [0:0] andOp_386_out;
	andOp #(.WIDTH(1)) andOp_386(.in0(andOp_386_in0), .in1(andOp_386_in1), .out(andOp_386_out));

	reg [0:0] notOp_387_in0;
	wire [0:0] notOp_387_out;
	notOp #(.WIDTH(1)) notOp_387(.in(notOp_387_in0), .out(notOp_387_out));

	reg [0:0] andOp_388_in0;
	reg [0:0] andOp_388_in1;
	wire [0:0] andOp_388_out;
	andOp #(.WIDTH(1)) andOp_388(.in0(andOp_388_in0), .in1(andOp_388_in1), .out(andOp_388_out));

	reg [0:0] andOp_389_in0;
	reg [0:0] andOp_389_in1;
	wire [0:0] andOp_389_out;
	andOp #(.WIDTH(1)) andOp_389(.in0(andOp_389_in0), .in1(andOp_389_in1), .out(andOp_389_out));

	reg [31:0] eq_390_in0;
	reg [31:0] eq_390_in1;
	wire [0:0] eq_390_out;
	eq #(.WIDTH(32)) eq_390(.in0(eq_390_in0), .in1(eq_390_in1), .out(eq_390_out));

	reg [0:0] andOp_391_in0;
	reg [0:0] andOp_391_in1;
	wire [0:0] andOp_391_out;
	andOp #(.WIDTH(1)) andOp_391(.in0(andOp_391_in0), .in1(andOp_391_in1), .out(andOp_391_out));

	reg [0:0] notOp_392_in0;
	wire [0:0] notOp_392_out;
	notOp #(.WIDTH(1)) notOp_392(.in(notOp_392_in0), .out(notOp_392_out));

	reg [0:0] andOp_393_in0;
	reg [0:0] andOp_393_in1;
	wire [0:0] andOp_393_out;
	andOp #(.WIDTH(1)) andOp_393(.in0(andOp_393_in0), .in1(andOp_393_in1), .out(andOp_393_out));

	reg [0:0] notOp_394_in0;
	wire [0:0] notOp_394_out;
	notOp #(.WIDTH(1)) notOp_394(.in(notOp_394_in0), .out(notOp_394_out));

	reg [0:0] andOp_395_in0;
	reg [0:0] andOp_395_in1;
	wire [0:0] andOp_395_out;
	andOp #(.WIDTH(1)) andOp_395(.in0(andOp_395_in0), .in1(andOp_395_in1), .out(andOp_395_out));

	reg [0:0] notOp_396_in0;
	wire [0:0] notOp_396_out;
	notOp #(.WIDTH(1)) notOp_396(.in(notOp_396_in0), .out(notOp_396_out));

	reg [0:0] andOp_397_in0;
	reg [0:0] andOp_397_in1;
	wire [0:0] andOp_397_out;
	andOp #(.WIDTH(1)) andOp_397(.in0(andOp_397_in0), .in1(andOp_397_in1), .out(andOp_397_out));

	reg [0:0] andOp_398_in0;
	reg [0:0] andOp_398_in1;
	wire [0:0] andOp_398_out;
	andOp #(.WIDTH(1)) andOp_398(.in0(andOp_398_in0), .in1(andOp_398_in1), .out(andOp_398_out));

	reg [31:0] eq_399_in0;
	reg [31:0] eq_399_in1;
	wire [0:0] eq_399_out;
	eq #(.WIDTH(32)) eq_399(.in0(eq_399_in0), .in1(eq_399_in1), .out(eq_399_out));

	reg [0:0] andOp_400_in0;
	reg [0:0] andOp_400_in1;
	wire [0:0] andOp_400_out;
	andOp #(.WIDTH(1)) andOp_400(.in0(andOp_400_in0), .in1(andOp_400_in1), .out(andOp_400_out));

	reg [0:0] notOp_401_in0;
	wire [0:0] notOp_401_out;
	notOp #(.WIDTH(1)) notOp_401(.in(notOp_401_in0), .out(notOp_401_out));

	reg [0:0] andOp_402_in0;
	reg [0:0] andOp_402_in1;
	wire [0:0] andOp_402_out;
	andOp #(.WIDTH(1)) andOp_402(.in0(andOp_402_in0), .in1(andOp_402_in1), .out(andOp_402_out));

	reg [0:0] notOp_403_in0;
	wire [0:0] notOp_403_out;
	notOp #(.WIDTH(1)) notOp_403(.in(notOp_403_in0), .out(notOp_403_out));

	reg [0:0] andOp_404_in0;
	reg [0:0] andOp_404_in1;
	wire [0:0] andOp_404_out;
	andOp #(.WIDTH(1)) andOp_404(.in0(andOp_404_in0), .in1(andOp_404_in1), .out(andOp_404_out));

	reg [0:0] notOp_405_in0;
	wire [0:0] notOp_405_out;
	notOp #(.WIDTH(1)) notOp_405(.in(notOp_405_in0), .out(notOp_405_out));

	reg [0:0] andOp_406_in0;
	reg [0:0] andOp_406_in1;
	wire [0:0] andOp_406_out;
	andOp #(.WIDTH(1)) andOp_406(.in0(andOp_406_in0), .in1(andOp_406_in1), .out(andOp_406_out));

	reg [0:0] andOp_407_in0;
	reg [0:0] andOp_407_in1;
	wire [0:0] andOp_407_out;
	andOp #(.WIDTH(1)) andOp_407(.in0(andOp_407_in0), .in1(andOp_407_in1), .out(andOp_407_out));

	reg [31:0] eq_408_in0;
	reg [31:0] eq_408_in1;
	wire [0:0] eq_408_out;
	eq #(.WIDTH(32)) eq_408(.in0(eq_408_in0), .in1(eq_408_in1), .out(eq_408_out));

	reg [0:0] andOp_409_in0;
	reg [0:0] andOp_409_in1;
	wire [0:0] andOp_409_out;
	andOp #(.WIDTH(1)) andOp_409(.in0(andOp_409_in0), .in1(andOp_409_in1), .out(andOp_409_out));

	reg [0:0] notOp_410_in0;
	wire [0:0] notOp_410_out;
	notOp #(.WIDTH(1)) notOp_410(.in(notOp_410_in0), .out(notOp_410_out));

	reg [0:0] andOp_411_in0;
	reg [0:0] andOp_411_in1;
	wire [0:0] andOp_411_out;
	andOp #(.WIDTH(1)) andOp_411(.in0(andOp_411_in0), .in1(andOp_411_in1), .out(andOp_411_out));

	reg [0:0] notOp_412_in0;
	wire [0:0] notOp_412_out;
	notOp #(.WIDTH(1)) notOp_412(.in(notOp_412_in0), .out(notOp_412_out));

	reg [0:0] andOp_413_in0;
	reg [0:0] andOp_413_in1;
	wire [0:0] andOp_413_out;
	andOp #(.WIDTH(1)) andOp_413(.in0(andOp_413_in0), .in1(andOp_413_in1), .out(andOp_413_out));

	reg [0:0] notOp_414_in0;
	wire [0:0] notOp_414_out;
	notOp #(.WIDTH(1)) notOp_414(.in(notOp_414_in0), .out(notOp_414_out));

	reg [0:0] andOp_415_in0;
	reg [0:0] andOp_415_in1;
	wire [0:0] andOp_415_out;
	andOp #(.WIDTH(1)) andOp_415(.in0(andOp_415_in0), .in1(andOp_415_in1), .out(andOp_415_out));

	reg [0:0] andOp_416_in0;
	reg [0:0] andOp_416_in1;
	wire [0:0] andOp_416_out;
	andOp #(.WIDTH(1)) andOp_416(.in0(andOp_416_in0), .in1(andOp_416_in1), .out(andOp_416_out));

	reg [31:0] eq_417_in0;
	reg [31:0] eq_417_in1;
	wire [0:0] eq_417_out;
	eq #(.WIDTH(32)) eq_417(.in0(eq_417_in0), .in1(eq_417_in1), .out(eq_417_out));

	reg [0:0] andOp_418_in0;
	reg [0:0] andOp_418_in1;
	wire [0:0] andOp_418_out;
	andOp #(.WIDTH(1)) andOp_418(.in0(andOp_418_in0), .in1(andOp_418_in1), .out(andOp_418_out));

	reg [0:0] notOp_419_in0;
	wire [0:0] notOp_419_out;
	notOp #(.WIDTH(1)) notOp_419(.in(notOp_419_in0), .out(notOp_419_out));

	reg [0:0] andOp_420_in0;
	reg [0:0] andOp_420_in1;
	wire [0:0] andOp_420_out;
	andOp #(.WIDTH(1)) andOp_420(.in0(andOp_420_in0), .in1(andOp_420_in1), .out(andOp_420_out));

	reg [0:0] notOp_421_in0;
	wire [0:0] notOp_421_out;
	notOp #(.WIDTH(1)) notOp_421(.in(notOp_421_in0), .out(notOp_421_out));

	reg [0:0] andOp_422_in0;
	reg [0:0] andOp_422_in1;
	wire [0:0] andOp_422_out;
	andOp #(.WIDTH(1)) andOp_422(.in0(andOp_422_in0), .in1(andOp_422_in1), .out(andOp_422_out));

	reg [0:0] notOp_423_in0;
	wire [0:0] notOp_423_out;
	notOp #(.WIDTH(1)) notOp_423(.in(notOp_423_in0), .out(notOp_423_out));

	reg [0:0] andOp_424_in0;
	reg [0:0] andOp_424_in1;
	wire [0:0] andOp_424_out;
	andOp #(.WIDTH(1)) andOp_424(.in0(andOp_424_in0), .in1(andOp_424_in1), .out(andOp_424_out));

	reg [31:0] eq_425_in0;
	reg [31:0] eq_425_in1;
	wire [0:0] eq_425_out;
	eq #(.WIDTH(32)) eq_425(.in0(eq_425_in0), .in1(eq_425_in1), .out(eq_425_out));

	reg [0:0] andOp_426_in0;
	reg [0:0] andOp_426_in1;
	wire [0:0] andOp_426_out;
	andOp #(.WIDTH(1)) andOp_426(.in0(andOp_426_in0), .in1(andOp_426_in1), .out(andOp_426_out));

	reg [31:0] eq_427_in0;
	reg [31:0] eq_427_in1;
	wire [0:0] eq_427_out;
	eq #(.WIDTH(32)) eq_427(.in0(eq_427_in0), .in1(eq_427_in1), .out(eq_427_out));

	reg [0:0] andOp_428_in0;
	reg [0:0] andOp_428_in1;
	wire [0:0] andOp_428_out;
	andOp #(.WIDTH(1)) andOp_428(.in0(andOp_428_in0), .in1(andOp_428_in1), .out(andOp_428_out));

	reg [31:0] eq_429_in0;
	reg [31:0] eq_429_in1;
	wire [0:0] eq_429_out;
	eq #(.WIDTH(32)) eq_429(.in0(eq_429_in0), .in1(eq_429_in1), .out(eq_429_out));

	reg [0:0] andOp_430_in0;
	reg [0:0] andOp_430_in1;
	wire [0:0] andOp_430_out;
	andOp #(.WIDTH(1)) andOp_430(.in0(andOp_430_in0), .in1(andOp_430_in1), .out(andOp_430_out));

	reg [31:0] eq_431_in0;
	reg [31:0] eq_431_in1;
	wire [0:0] eq_431_out;
	eq #(.WIDTH(32)) eq_431(.in0(eq_431_in0), .in1(eq_431_in1), .out(eq_431_out));

	reg [0:0] andOp_432_in0;
	reg [0:0] andOp_432_in1;
	wire [0:0] andOp_432_out;
	andOp #(.WIDTH(1)) andOp_432(.in0(andOp_432_in0), .in1(andOp_432_in1), .out(andOp_432_out));

	reg [31:0] eq_433_in0;
	reg [31:0] eq_433_in1;
	wire [0:0] eq_433_out;
	eq #(.WIDTH(32)) eq_433(.in0(eq_433_in0), .in1(eq_433_in1), .out(eq_433_out));

	reg [0:0] andOp_434_in0;
	reg [0:0] andOp_434_in1;
	wire [0:0] andOp_434_out;
	andOp #(.WIDTH(1)) andOp_434(.in0(andOp_434_in0), .in1(andOp_434_in1), .out(andOp_434_out));

	reg [0:0] andOp_435_in0;
	reg [0:0] andOp_435_in1;
	wire [0:0] andOp_435_out;
	andOp #(.WIDTH(1)) andOp_435(.in0(andOp_435_in0), .in1(andOp_435_in1), .out(andOp_435_out));

	reg [31:0] eq_436_in0;
	reg [31:0] eq_436_in1;
	wire [0:0] eq_436_out;
	eq #(.WIDTH(32)) eq_436(.in0(eq_436_in0), .in1(eq_436_in1), .out(eq_436_out));

	reg [0:0] andOp_437_in0;
	reg [0:0] andOp_437_in1;
	wire [0:0] andOp_437_out;
	andOp #(.WIDTH(1)) andOp_437(.in0(andOp_437_in0), .in1(andOp_437_in1), .out(andOp_437_out));

	reg [0:0] notOp_438_in0;
	wire [0:0] notOp_438_out;
	notOp #(.WIDTH(1)) notOp_438(.in(notOp_438_in0), .out(notOp_438_out));

	reg [0:0] andOp_439_in0;
	reg [0:0] andOp_439_in1;
	wire [0:0] andOp_439_out;
	andOp #(.WIDTH(1)) andOp_439(.in0(andOp_439_in0), .in1(andOp_439_in1), .out(andOp_439_out));

	reg [0:0] notOp_440_in0;
	wire [0:0] notOp_440_out;
	notOp #(.WIDTH(1)) notOp_440(.in(notOp_440_in0), .out(notOp_440_out));

	reg [0:0] andOp_441_in0;
	reg [0:0] andOp_441_in1;
	wire [0:0] andOp_441_out;
	andOp #(.WIDTH(1)) andOp_441(.in0(andOp_441_in0), .in1(andOp_441_in1), .out(andOp_441_out));

	reg [0:0] notOp_442_in0;
	wire [0:0] notOp_442_out;
	notOp #(.WIDTH(1)) notOp_442(.in(notOp_442_in0), .out(notOp_442_out));

	reg [0:0] andOp_443_in0;
	reg [0:0] andOp_443_in1;
	wire [0:0] andOp_443_out;
	andOp #(.WIDTH(1)) andOp_443(.in0(andOp_443_in0), .in1(andOp_443_in1), .out(andOp_443_out));

	reg [0:0] andOp_444_in0;
	reg [0:0] andOp_444_in1;
	wire [0:0] andOp_444_out;
	andOp #(.WIDTH(1)) andOp_444(.in0(andOp_444_in0), .in1(andOp_444_in1), .out(andOp_444_out));

	reg [31:0] eq_445_in0;
	reg [31:0] eq_445_in1;
	wire [0:0] eq_445_out;
	eq #(.WIDTH(32)) eq_445(.in0(eq_445_in0), .in1(eq_445_in1), .out(eq_445_out));

	reg [0:0] andOp_446_in0;
	reg [0:0] andOp_446_in1;
	wire [0:0] andOp_446_out;
	andOp #(.WIDTH(1)) andOp_446(.in0(andOp_446_in0), .in1(andOp_446_in1), .out(andOp_446_out));

	reg [0:0] notOp_447_in0;
	wire [0:0] notOp_447_out;
	notOp #(.WIDTH(1)) notOp_447(.in(notOp_447_in0), .out(notOp_447_out));

	reg [0:0] andOp_448_in0;
	reg [0:0] andOp_448_in1;
	wire [0:0] andOp_448_out;
	andOp #(.WIDTH(1)) andOp_448(.in0(andOp_448_in0), .in1(andOp_448_in1), .out(andOp_448_out));

	reg [0:0] notOp_449_in0;
	wire [0:0] notOp_449_out;
	notOp #(.WIDTH(1)) notOp_449(.in(notOp_449_in0), .out(notOp_449_out));

	reg [0:0] andOp_450_in0;
	reg [0:0] andOp_450_in1;
	wire [0:0] andOp_450_out;
	andOp #(.WIDTH(1)) andOp_450(.in0(andOp_450_in0), .in1(andOp_450_in1), .out(andOp_450_out));

	reg [0:0] notOp_451_in0;
	wire [0:0] notOp_451_out;
	notOp #(.WIDTH(1)) notOp_451(.in(notOp_451_in0), .out(notOp_451_out));

	reg [0:0] andOp_452_in0;
	reg [0:0] andOp_452_in1;
	wire [0:0] andOp_452_out;
	andOp #(.WIDTH(1)) andOp_452(.in0(andOp_452_in0), .in1(andOp_452_in1), .out(andOp_452_out));

	reg [0:0] andOp_453_in0;
	reg [0:0] andOp_453_in1;
	wire [0:0] andOp_453_out;
	andOp #(.WIDTH(1)) andOp_453(.in0(andOp_453_in0), .in1(andOp_453_in1), .out(andOp_453_out));

	reg [31:0] eq_454_in0;
	reg [31:0] eq_454_in1;
	wire [0:0] eq_454_out;
	eq #(.WIDTH(32)) eq_454(.in0(eq_454_in0), .in1(eq_454_in1), .out(eq_454_out));

	reg [0:0] andOp_455_in0;
	reg [0:0] andOp_455_in1;
	wire [0:0] andOp_455_out;
	andOp #(.WIDTH(1)) andOp_455(.in0(andOp_455_in0), .in1(andOp_455_in1), .out(andOp_455_out));

	reg [0:0] notOp_456_in0;
	wire [0:0] notOp_456_out;
	notOp #(.WIDTH(1)) notOp_456(.in(notOp_456_in0), .out(notOp_456_out));

	reg [0:0] andOp_457_in0;
	reg [0:0] andOp_457_in1;
	wire [0:0] andOp_457_out;
	andOp #(.WIDTH(1)) andOp_457(.in0(andOp_457_in0), .in1(andOp_457_in1), .out(andOp_457_out));

	reg [0:0] notOp_458_in0;
	wire [0:0] notOp_458_out;
	notOp #(.WIDTH(1)) notOp_458(.in(notOp_458_in0), .out(notOp_458_out));

	reg [0:0] andOp_459_in0;
	reg [0:0] andOp_459_in1;
	wire [0:0] andOp_459_out;
	andOp #(.WIDTH(1)) andOp_459(.in0(andOp_459_in0), .in1(andOp_459_in1), .out(andOp_459_out));

	reg [0:0] notOp_460_in0;
	wire [0:0] notOp_460_out;
	notOp #(.WIDTH(1)) notOp_460(.in(notOp_460_in0), .out(notOp_460_out));

	reg [0:0] andOp_461_in0;
	reg [0:0] andOp_461_in1;
	wire [0:0] andOp_461_out;
	andOp #(.WIDTH(1)) andOp_461(.in0(andOp_461_in0), .in1(andOp_461_in1), .out(andOp_461_out));

	reg [0:0] andOp_462_in0;
	reg [0:0] andOp_462_in1;
	wire [0:0] andOp_462_out;
	andOp #(.WIDTH(1)) andOp_462(.in0(andOp_462_in0), .in1(andOp_462_in1), .out(andOp_462_out));

	reg [31:0] eq_463_in0;
	reg [31:0] eq_463_in1;
	wire [0:0] eq_463_out;
	eq #(.WIDTH(32)) eq_463(.in0(eq_463_in0), .in1(eq_463_in1), .out(eq_463_out));

	reg [0:0] andOp_464_in0;
	reg [0:0] andOp_464_in1;
	wire [0:0] andOp_464_out;
	andOp #(.WIDTH(1)) andOp_464(.in0(andOp_464_in0), .in1(andOp_464_in1), .out(andOp_464_out));

	reg [0:0] notOp_465_in0;
	wire [0:0] notOp_465_out;
	notOp #(.WIDTH(1)) notOp_465(.in(notOp_465_in0), .out(notOp_465_out));

	reg [0:0] andOp_466_in0;
	reg [0:0] andOp_466_in1;
	wire [0:0] andOp_466_out;
	andOp #(.WIDTH(1)) andOp_466(.in0(andOp_466_in0), .in1(andOp_466_in1), .out(andOp_466_out));

	reg [0:0] notOp_467_in0;
	wire [0:0] notOp_467_out;
	notOp #(.WIDTH(1)) notOp_467(.in(notOp_467_in0), .out(notOp_467_out));

	reg [0:0] andOp_468_in0;
	reg [0:0] andOp_468_in1;
	wire [0:0] andOp_468_out;
	andOp #(.WIDTH(1)) andOp_468(.in0(andOp_468_in0), .in1(andOp_468_in1), .out(andOp_468_out));

	reg [0:0] notOp_469_in0;
	wire [0:0] notOp_469_out;
	notOp #(.WIDTH(1)) notOp_469(.in(notOp_469_in0), .out(notOp_469_out));

	reg [0:0] andOp_470_in0;
	reg [0:0] andOp_470_in1;
	wire [0:0] andOp_470_out;
	andOp #(.WIDTH(1)) andOp_470(.in0(andOp_470_in0), .in1(andOp_470_in1), .out(andOp_470_out));

	reg [0:0] andOp_471_in0;
	reg [0:0] andOp_471_in1;
	wire [0:0] andOp_471_out;
	andOp #(.WIDTH(1)) andOp_471(.in0(andOp_471_in0), .in1(andOp_471_in1), .out(andOp_471_out));

	reg [31:0] eq_472_in0;
	reg [31:0] eq_472_in1;
	wire [0:0] eq_472_out;
	eq #(.WIDTH(32)) eq_472(.in0(eq_472_in0), .in1(eq_472_in1), .out(eq_472_out));

	reg [0:0] andOp_473_in0;
	reg [0:0] andOp_473_in1;
	wire [0:0] andOp_473_out;
	andOp #(.WIDTH(1)) andOp_473(.in0(andOp_473_in0), .in1(andOp_473_in1), .out(andOp_473_out));

	reg [0:0] notOp_474_in0;
	wire [0:0] notOp_474_out;
	notOp #(.WIDTH(1)) notOp_474(.in(notOp_474_in0), .out(notOp_474_out));

	reg [0:0] andOp_475_in0;
	reg [0:0] andOp_475_in1;
	wire [0:0] andOp_475_out;
	andOp #(.WIDTH(1)) andOp_475(.in0(andOp_475_in0), .in1(andOp_475_in1), .out(andOp_475_out));

	reg [0:0] notOp_476_in0;
	wire [0:0] notOp_476_out;
	notOp #(.WIDTH(1)) notOp_476(.in(notOp_476_in0), .out(notOp_476_out));

	reg [0:0] andOp_477_in0;
	reg [0:0] andOp_477_in1;
	wire [0:0] andOp_477_out;
	andOp #(.WIDTH(1)) andOp_477(.in0(andOp_477_in0), .in1(andOp_477_in1), .out(andOp_477_out));

	reg [0:0] notOp_478_in0;
	wire [0:0] notOp_478_out;
	notOp #(.WIDTH(1)) notOp_478(.in(notOp_478_in0), .out(notOp_478_out));

	reg [0:0] andOp_479_in0;
	reg [0:0] andOp_479_in1;
	wire [0:0] andOp_479_out;
	andOp #(.WIDTH(1)) andOp_479(.in0(andOp_479_in0), .in1(andOp_479_in1), .out(andOp_479_out));

	reg [0:0] andOp_480_in0;
	reg [0:0] andOp_480_in1;
	wire [0:0] andOp_480_out;
	andOp #(.WIDTH(1)) andOp_480(.in0(andOp_480_in0), .in1(andOp_480_in1), .out(andOp_480_out));

	reg [31:0] eq_481_in0;
	reg [31:0] eq_481_in1;
	wire [0:0] eq_481_out;
	eq #(.WIDTH(32)) eq_481(.in0(eq_481_in0), .in1(eq_481_in1), .out(eq_481_out));

	reg [0:0] andOp_482_in0;
	reg [0:0] andOp_482_in1;
	wire [0:0] andOp_482_out;
	andOp #(.WIDTH(1)) andOp_482(.in0(andOp_482_in0), .in1(andOp_482_in1), .out(andOp_482_out));

	reg [0:0] notOp_483_in0;
	wire [0:0] notOp_483_out;
	notOp #(.WIDTH(1)) notOp_483(.in(notOp_483_in0), .out(notOp_483_out));

	reg [0:0] andOp_484_in0;
	reg [0:0] andOp_484_in1;
	wire [0:0] andOp_484_out;
	andOp #(.WIDTH(1)) andOp_484(.in0(andOp_484_in0), .in1(andOp_484_in1), .out(andOp_484_out));

	reg [0:0] notOp_485_in0;
	wire [0:0] notOp_485_out;
	notOp #(.WIDTH(1)) notOp_485(.in(notOp_485_in0), .out(notOp_485_out));

	reg [0:0] andOp_486_in0;
	reg [0:0] andOp_486_in1;
	wire [0:0] andOp_486_out;
	andOp #(.WIDTH(1)) andOp_486(.in0(andOp_486_in0), .in1(andOp_486_in1), .out(andOp_486_out));

	reg [0:0] notOp_487_in0;
	wire [0:0] notOp_487_out;
	notOp #(.WIDTH(1)) notOp_487(.in(notOp_487_in0), .out(notOp_487_out));

	reg [0:0] andOp_488_in0;
	reg [0:0] andOp_488_in1;
	wire [0:0] andOp_488_out;
	andOp #(.WIDTH(1)) andOp_488(.in0(andOp_488_in0), .in1(andOp_488_in1), .out(andOp_488_out));

	reg [0:0] andOp_489_in0;
	reg [0:0] andOp_489_in1;
	wire [0:0] andOp_489_out;
	andOp #(.WIDTH(1)) andOp_489(.in0(andOp_489_in0), .in1(andOp_489_in1), .out(andOp_489_out));

	reg [31:0] eq_490_in0;
	reg [31:0] eq_490_in1;
	wire [0:0] eq_490_out;
	eq #(.WIDTH(32)) eq_490(.in0(eq_490_in0), .in1(eq_490_in1), .out(eq_490_out));

	reg [0:0] andOp_491_in0;
	reg [0:0] andOp_491_in1;
	wire [0:0] andOp_491_out;
	andOp #(.WIDTH(1)) andOp_491(.in0(andOp_491_in0), .in1(andOp_491_in1), .out(andOp_491_out));

	reg [0:0] notOp_492_in0;
	wire [0:0] notOp_492_out;
	notOp #(.WIDTH(1)) notOp_492(.in(notOp_492_in0), .out(notOp_492_out));

	reg [0:0] andOp_493_in0;
	reg [0:0] andOp_493_in1;
	wire [0:0] andOp_493_out;
	andOp #(.WIDTH(1)) andOp_493(.in0(andOp_493_in0), .in1(andOp_493_in1), .out(andOp_493_out));

	reg [0:0] notOp_494_in0;
	wire [0:0] notOp_494_out;
	notOp #(.WIDTH(1)) notOp_494(.in(notOp_494_in0), .out(notOp_494_out));

	reg [0:0] andOp_495_in0;
	reg [0:0] andOp_495_in1;
	wire [0:0] andOp_495_out;
	andOp #(.WIDTH(1)) andOp_495(.in0(andOp_495_in0), .in1(andOp_495_in1), .out(andOp_495_out));

	reg [0:0] notOp_496_in0;
	wire [0:0] notOp_496_out;
	notOp #(.WIDTH(1)) notOp_496(.in(notOp_496_in0), .out(notOp_496_out));

	reg [0:0] andOp_497_in0;
	reg [0:0] andOp_497_in1;
	wire [0:0] andOp_497_out;
	andOp #(.WIDTH(1)) andOp_497(.in0(andOp_497_in0), .in1(andOp_497_in1), .out(andOp_497_out));

	reg [0:0] andOp_498_in0;
	reg [0:0] andOp_498_in1;
	wire [0:0] andOp_498_out;
	andOp #(.WIDTH(1)) andOp_498(.in0(andOp_498_in0), .in1(andOp_498_in1), .out(andOp_498_out));

	reg [31:0] eq_499_in0;
	reg [31:0] eq_499_in1;
	wire [0:0] eq_499_out;
	eq #(.WIDTH(32)) eq_499(.in0(eq_499_in0), .in1(eq_499_in1), .out(eq_499_out));

	reg [0:0] andOp_500_in0;
	reg [0:0] andOp_500_in1;
	wire [0:0] andOp_500_out;
	andOp #(.WIDTH(1)) andOp_500(.in0(andOp_500_in0), .in1(andOp_500_in1), .out(andOp_500_out));

	reg [0:0] notOp_501_in0;
	wire [0:0] notOp_501_out;
	notOp #(.WIDTH(1)) notOp_501(.in(notOp_501_in0), .out(notOp_501_out));

	reg [0:0] andOp_502_in0;
	reg [0:0] andOp_502_in1;
	wire [0:0] andOp_502_out;
	andOp #(.WIDTH(1)) andOp_502(.in0(andOp_502_in0), .in1(andOp_502_in1), .out(andOp_502_out));

	reg [0:0] notOp_503_in0;
	wire [0:0] notOp_503_out;
	notOp #(.WIDTH(1)) notOp_503(.in(notOp_503_in0), .out(notOp_503_out));

	reg [0:0] andOp_504_in0;
	reg [0:0] andOp_504_in1;
	wire [0:0] andOp_504_out;
	andOp #(.WIDTH(1)) andOp_504(.in0(andOp_504_in0), .in1(andOp_504_in1), .out(andOp_504_out));

	reg [0:0] notOp_505_in0;
	wire [0:0] notOp_505_out;
	notOp #(.WIDTH(1)) notOp_505(.in(notOp_505_in0), .out(notOp_505_out));

	reg [0:0] andOp_506_in0;
	reg [0:0] andOp_506_in1;
	wire [0:0] andOp_506_out;
	andOp #(.WIDTH(1)) andOp_506(.in0(andOp_506_in0), .in1(andOp_506_in1), .out(andOp_506_out));

	reg [0:0] andOp_507_in0;
	reg [0:0] andOp_507_in1;
	wire [0:0] andOp_507_out;
	andOp #(.WIDTH(1)) andOp_507(.in0(andOp_507_in0), .in1(andOp_507_in1), .out(andOp_507_out));

	reg [31:0] eq_508_in0;
	reg [31:0] eq_508_in1;
	wire [0:0] eq_508_out;
	eq #(.WIDTH(32)) eq_508(.in0(eq_508_in0), .in1(eq_508_in1), .out(eq_508_out));

	reg [0:0] andOp_509_in0;
	reg [0:0] andOp_509_in1;
	wire [0:0] andOp_509_out;
	andOp #(.WIDTH(1)) andOp_509(.in0(andOp_509_in0), .in1(andOp_509_in1), .out(andOp_509_out));

	reg [0:0] notOp_510_in0;
	wire [0:0] notOp_510_out;
	notOp #(.WIDTH(1)) notOp_510(.in(notOp_510_in0), .out(notOp_510_out));

	reg [0:0] andOp_511_in0;
	reg [0:0] andOp_511_in1;
	wire [0:0] andOp_511_out;
	andOp #(.WIDTH(1)) andOp_511(.in0(andOp_511_in0), .in1(andOp_511_in1), .out(andOp_511_out));

	reg [0:0] notOp_512_in0;
	wire [0:0] notOp_512_out;
	notOp #(.WIDTH(1)) notOp_512(.in(notOp_512_in0), .out(notOp_512_out));

	reg [0:0] andOp_513_in0;
	reg [0:0] andOp_513_in1;
	wire [0:0] andOp_513_out;
	andOp #(.WIDTH(1)) andOp_513(.in0(andOp_513_in0), .in1(andOp_513_in1), .out(andOp_513_out));

	reg [0:0] notOp_514_in0;
	wire [0:0] notOp_514_out;
	notOp #(.WIDTH(1)) notOp_514(.in(notOp_514_in0), .out(notOp_514_out));

	reg [0:0] andOp_515_in0;
	reg [0:0] andOp_515_in1;
	wire [0:0] andOp_515_out;
	andOp #(.WIDTH(1)) andOp_515(.in0(andOp_515_in0), .in1(andOp_515_in1), .out(andOp_515_out));

	reg [31:0] eq_516_in0;
	reg [31:0] eq_516_in1;
	wire [0:0] eq_516_out;
	eq #(.WIDTH(32)) eq_516(.in0(eq_516_in0), .in1(eq_516_in1), .out(eq_516_out));

	reg [0:0] andOp_517_in0;
	reg [0:0] andOp_517_in1;
	wire [0:0] andOp_517_out;
	andOp #(.WIDTH(1)) andOp_517(.in0(andOp_517_in0), .in1(andOp_517_in1), .out(andOp_517_out));

	reg [31:0] eq_518_in0;
	reg [31:0] eq_518_in1;
	wire [0:0] eq_518_out;
	eq #(.WIDTH(32)) eq_518(.in0(eq_518_in0), .in1(eq_518_in1), .out(eq_518_out));

	reg [0:0] andOp_519_in0;
	reg [0:0] andOp_519_in1;
	wire [0:0] andOp_519_out;
	andOp #(.WIDTH(1)) andOp_519(.in0(andOp_519_in0), .in1(andOp_519_in1), .out(andOp_519_out));

	reg [31:0] eq_520_in0;
	reg [31:0] eq_520_in1;
	wire [0:0] eq_520_out;
	eq #(.WIDTH(32)) eq_520(.in0(eq_520_in0), .in1(eq_520_in1), .out(eq_520_out));

	reg [0:0] andOp_521_in0;
	reg [0:0] andOp_521_in1;
	wire [0:0] andOp_521_out;
	andOp #(.WIDTH(1)) andOp_521(.in0(andOp_521_in0), .in1(andOp_521_in1), .out(andOp_521_out));

	reg [31:0] eq_522_in0;
	reg [31:0] eq_522_in1;
	wire [0:0] eq_522_out;
	eq #(.WIDTH(32)) eq_522(.in0(eq_522_in0), .in1(eq_522_in1), .out(eq_522_out));

	reg [0:0] andOp_523_in0;
	reg [0:0] andOp_523_in1;
	wire [0:0] andOp_523_out;
	andOp #(.WIDTH(1)) andOp_523(.in0(andOp_523_in0), .in1(andOp_523_in1), .out(andOp_523_out));

	reg [31:0] eq_524_in0;
	reg [31:0] eq_524_in1;
	wire [0:0] eq_524_out;
	eq #(.WIDTH(32)) eq_524(.in0(eq_524_in0), .in1(eq_524_in1), .out(eq_524_out));

	reg [0:0] andOp_525_in0;
	reg [0:0] andOp_525_in1;
	wire [0:0] andOp_525_out;
	andOp #(.WIDTH(1)) andOp_525(.in0(andOp_525_in0), .in1(andOp_525_in1), .out(andOp_525_out));

	reg [0:0] andOp_526_in0;
	reg [0:0] andOp_526_in1;
	wire [0:0] andOp_526_out;
	andOp #(.WIDTH(1)) andOp_526(.in0(andOp_526_in0), .in1(andOp_526_in1), .out(andOp_526_out));

	reg [31:0] eq_527_in0;
	reg [31:0] eq_527_in1;
	wire [0:0] eq_527_out;
	eq #(.WIDTH(32)) eq_527(.in0(eq_527_in0), .in1(eq_527_in1), .out(eq_527_out));

	reg [0:0] andOp_528_in0;
	reg [0:0] andOp_528_in1;
	wire [0:0] andOp_528_out;
	andOp #(.WIDTH(1)) andOp_528(.in0(andOp_528_in0), .in1(andOp_528_in1), .out(andOp_528_out));

	reg [0:0] notOp_529_in0;
	wire [0:0] notOp_529_out;
	notOp #(.WIDTH(1)) notOp_529(.in(notOp_529_in0), .out(notOp_529_out));

	reg [0:0] andOp_530_in0;
	reg [0:0] andOp_530_in1;
	wire [0:0] andOp_530_out;
	andOp #(.WIDTH(1)) andOp_530(.in0(andOp_530_in0), .in1(andOp_530_in1), .out(andOp_530_out));

	reg [0:0] notOp_531_in0;
	wire [0:0] notOp_531_out;
	notOp #(.WIDTH(1)) notOp_531(.in(notOp_531_in0), .out(notOp_531_out));

	reg [0:0] andOp_532_in0;
	reg [0:0] andOp_532_in1;
	wire [0:0] andOp_532_out;
	andOp #(.WIDTH(1)) andOp_532(.in0(andOp_532_in0), .in1(andOp_532_in1), .out(andOp_532_out));

	reg [0:0] notOp_533_in0;
	wire [0:0] notOp_533_out;
	notOp #(.WIDTH(1)) notOp_533(.in(notOp_533_in0), .out(notOp_533_out));

	reg [0:0] andOp_534_in0;
	reg [0:0] andOp_534_in1;
	wire [0:0] andOp_534_out;
	andOp #(.WIDTH(1)) andOp_534(.in0(andOp_534_in0), .in1(andOp_534_in1), .out(andOp_534_out));

	reg [0:0] andOp_535_in0;
	reg [0:0] andOp_535_in1;
	wire [0:0] andOp_535_out;
	andOp #(.WIDTH(1)) andOp_535(.in0(andOp_535_in0), .in1(andOp_535_in1), .out(andOp_535_out));

	reg [31:0] eq_536_in0;
	reg [31:0] eq_536_in1;
	wire [0:0] eq_536_out;
	eq #(.WIDTH(32)) eq_536(.in0(eq_536_in0), .in1(eq_536_in1), .out(eq_536_out));

	reg [0:0] andOp_537_in0;
	reg [0:0] andOp_537_in1;
	wire [0:0] andOp_537_out;
	andOp #(.WIDTH(1)) andOp_537(.in0(andOp_537_in0), .in1(andOp_537_in1), .out(andOp_537_out));

	reg [0:0] notOp_538_in0;
	wire [0:0] notOp_538_out;
	notOp #(.WIDTH(1)) notOp_538(.in(notOp_538_in0), .out(notOp_538_out));

	reg [0:0] andOp_539_in0;
	reg [0:0] andOp_539_in1;
	wire [0:0] andOp_539_out;
	andOp #(.WIDTH(1)) andOp_539(.in0(andOp_539_in0), .in1(andOp_539_in1), .out(andOp_539_out));

	reg [0:0] notOp_540_in0;
	wire [0:0] notOp_540_out;
	notOp #(.WIDTH(1)) notOp_540(.in(notOp_540_in0), .out(notOp_540_out));

	reg [0:0] andOp_541_in0;
	reg [0:0] andOp_541_in1;
	wire [0:0] andOp_541_out;
	andOp #(.WIDTH(1)) andOp_541(.in0(andOp_541_in0), .in1(andOp_541_in1), .out(andOp_541_out));

	reg [0:0] notOp_542_in0;
	wire [0:0] notOp_542_out;
	notOp #(.WIDTH(1)) notOp_542(.in(notOp_542_in0), .out(notOp_542_out));

	reg [0:0] andOp_543_in0;
	reg [0:0] andOp_543_in1;
	wire [0:0] andOp_543_out;
	andOp #(.WIDTH(1)) andOp_543(.in0(andOp_543_in0), .in1(andOp_543_in1), .out(andOp_543_out));

	reg [0:0] andOp_544_in0;
	reg [0:0] andOp_544_in1;
	wire [0:0] andOp_544_out;
	andOp #(.WIDTH(1)) andOp_544(.in0(andOp_544_in0), .in1(andOp_544_in1), .out(andOp_544_out));

	reg [31:0] eq_545_in0;
	reg [31:0] eq_545_in1;
	wire [0:0] eq_545_out;
	eq #(.WIDTH(32)) eq_545(.in0(eq_545_in0), .in1(eq_545_in1), .out(eq_545_out));

	reg [0:0] andOp_546_in0;
	reg [0:0] andOp_546_in1;
	wire [0:0] andOp_546_out;
	andOp #(.WIDTH(1)) andOp_546(.in0(andOp_546_in0), .in1(andOp_546_in1), .out(andOp_546_out));

	reg [0:0] notOp_547_in0;
	wire [0:0] notOp_547_out;
	notOp #(.WIDTH(1)) notOp_547(.in(notOp_547_in0), .out(notOp_547_out));

	reg [0:0] andOp_548_in0;
	reg [0:0] andOp_548_in1;
	wire [0:0] andOp_548_out;
	andOp #(.WIDTH(1)) andOp_548(.in0(andOp_548_in0), .in1(andOp_548_in1), .out(andOp_548_out));

	reg [0:0] notOp_549_in0;
	wire [0:0] notOp_549_out;
	notOp #(.WIDTH(1)) notOp_549(.in(notOp_549_in0), .out(notOp_549_out));

	reg [0:0] andOp_550_in0;
	reg [0:0] andOp_550_in1;
	wire [0:0] andOp_550_out;
	andOp #(.WIDTH(1)) andOp_550(.in0(andOp_550_in0), .in1(andOp_550_in1), .out(andOp_550_out));

	reg [0:0] notOp_551_in0;
	wire [0:0] notOp_551_out;
	notOp #(.WIDTH(1)) notOp_551(.in(notOp_551_in0), .out(notOp_551_out));

	reg [0:0] andOp_552_in0;
	reg [0:0] andOp_552_in1;
	wire [0:0] andOp_552_out;
	andOp #(.WIDTH(1)) andOp_552(.in0(andOp_552_in0), .in1(andOp_552_in1), .out(andOp_552_out));

	reg [0:0] andOp_553_in0;
	reg [0:0] andOp_553_in1;
	wire [0:0] andOp_553_out;
	andOp #(.WIDTH(1)) andOp_553(.in0(andOp_553_in0), .in1(andOp_553_in1), .out(andOp_553_out));

	reg [31:0] eq_554_in0;
	reg [31:0] eq_554_in1;
	wire [0:0] eq_554_out;
	eq #(.WIDTH(32)) eq_554(.in0(eq_554_in0), .in1(eq_554_in1), .out(eq_554_out));

	reg [0:0] andOp_555_in0;
	reg [0:0] andOp_555_in1;
	wire [0:0] andOp_555_out;
	andOp #(.WIDTH(1)) andOp_555(.in0(andOp_555_in0), .in1(andOp_555_in1), .out(andOp_555_out));

	reg [0:0] notOp_556_in0;
	wire [0:0] notOp_556_out;
	notOp #(.WIDTH(1)) notOp_556(.in(notOp_556_in0), .out(notOp_556_out));

	reg [0:0] andOp_557_in0;
	reg [0:0] andOp_557_in1;
	wire [0:0] andOp_557_out;
	andOp #(.WIDTH(1)) andOp_557(.in0(andOp_557_in0), .in1(andOp_557_in1), .out(andOp_557_out));

	reg [0:0] notOp_558_in0;
	wire [0:0] notOp_558_out;
	notOp #(.WIDTH(1)) notOp_558(.in(notOp_558_in0), .out(notOp_558_out));

	reg [0:0] andOp_559_in0;
	reg [0:0] andOp_559_in1;
	wire [0:0] andOp_559_out;
	andOp #(.WIDTH(1)) andOp_559(.in0(andOp_559_in0), .in1(andOp_559_in1), .out(andOp_559_out));

	reg [0:0] notOp_560_in0;
	wire [0:0] notOp_560_out;
	notOp #(.WIDTH(1)) notOp_560(.in(notOp_560_in0), .out(notOp_560_out));

	reg [0:0] andOp_561_in0;
	reg [0:0] andOp_561_in1;
	wire [0:0] andOp_561_out;
	andOp #(.WIDTH(1)) andOp_561(.in0(andOp_561_in0), .in1(andOp_561_in1), .out(andOp_561_out));

	reg [0:0] andOp_562_in0;
	reg [0:0] andOp_562_in1;
	wire [0:0] andOp_562_out;
	andOp #(.WIDTH(1)) andOp_562(.in0(andOp_562_in0), .in1(andOp_562_in1), .out(andOp_562_out));

	reg [31:0] eq_563_in0;
	reg [31:0] eq_563_in1;
	wire [0:0] eq_563_out;
	eq #(.WIDTH(32)) eq_563(.in0(eq_563_in0), .in1(eq_563_in1), .out(eq_563_out));

	reg [0:0] andOp_564_in0;
	reg [0:0] andOp_564_in1;
	wire [0:0] andOp_564_out;
	andOp #(.WIDTH(1)) andOp_564(.in0(andOp_564_in0), .in1(andOp_564_in1), .out(andOp_564_out));

	reg [0:0] notOp_565_in0;
	wire [0:0] notOp_565_out;
	notOp #(.WIDTH(1)) notOp_565(.in(notOp_565_in0), .out(notOp_565_out));

	reg [0:0] andOp_566_in0;
	reg [0:0] andOp_566_in1;
	wire [0:0] andOp_566_out;
	andOp #(.WIDTH(1)) andOp_566(.in0(andOp_566_in0), .in1(andOp_566_in1), .out(andOp_566_out));

	reg [0:0] notOp_567_in0;
	wire [0:0] notOp_567_out;
	notOp #(.WIDTH(1)) notOp_567(.in(notOp_567_in0), .out(notOp_567_out));

	reg [0:0] andOp_568_in0;
	reg [0:0] andOp_568_in1;
	wire [0:0] andOp_568_out;
	andOp #(.WIDTH(1)) andOp_568(.in0(andOp_568_in0), .in1(andOp_568_in1), .out(andOp_568_out));

	reg [0:0] notOp_569_in0;
	wire [0:0] notOp_569_out;
	notOp #(.WIDTH(1)) notOp_569(.in(notOp_569_in0), .out(notOp_569_out));

	reg [0:0] andOp_570_in0;
	reg [0:0] andOp_570_in1;
	wire [0:0] andOp_570_out;
	andOp #(.WIDTH(1)) andOp_570(.in0(andOp_570_in0), .in1(andOp_570_in1), .out(andOp_570_out));

	reg [0:0] andOp_571_in0;
	reg [0:0] andOp_571_in1;
	wire [0:0] andOp_571_out;
	andOp #(.WIDTH(1)) andOp_571(.in0(andOp_571_in0), .in1(andOp_571_in1), .out(andOp_571_out));

	reg [31:0] eq_572_in0;
	reg [31:0] eq_572_in1;
	wire [0:0] eq_572_out;
	eq #(.WIDTH(32)) eq_572(.in0(eq_572_in0), .in1(eq_572_in1), .out(eq_572_out));

	reg [0:0] andOp_573_in0;
	reg [0:0] andOp_573_in1;
	wire [0:0] andOp_573_out;
	andOp #(.WIDTH(1)) andOp_573(.in0(andOp_573_in0), .in1(andOp_573_in1), .out(andOp_573_out));

	reg [0:0] notOp_574_in0;
	wire [0:0] notOp_574_out;
	notOp #(.WIDTH(1)) notOp_574(.in(notOp_574_in0), .out(notOp_574_out));

	reg [0:0] andOp_575_in0;
	reg [0:0] andOp_575_in1;
	wire [0:0] andOp_575_out;
	andOp #(.WIDTH(1)) andOp_575(.in0(andOp_575_in0), .in1(andOp_575_in1), .out(andOp_575_out));

	reg [0:0] notOp_576_in0;
	wire [0:0] notOp_576_out;
	notOp #(.WIDTH(1)) notOp_576(.in(notOp_576_in0), .out(notOp_576_out));

	reg [0:0] andOp_577_in0;
	reg [0:0] andOp_577_in1;
	wire [0:0] andOp_577_out;
	andOp #(.WIDTH(1)) andOp_577(.in0(andOp_577_in0), .in1(andOp_577_in1), .out(andOp_577_out));

	reg [0:0] notOp_578_in0;
	wire [0:0] notOp_578_out;
	notOp #(.WIDTH(1)) notOp_578(.in(notOp_578_in0), .out(notOp_578_out));

	reg [0:0] andOp_579_in0;
	reg [0:0] andOp_579_in1;
	wire [0:0] andOp_579_out;
	andOp #(.WIDTH(1)) andOp_579(.in0(andOp_579_in0), .in1(andOp_579_in1), .out(andOp_579_out));

	reg [0:0] andOp_580_in0;
	reg [0:0] andOp_580_in1;
	wire [0:0] andOp_580_out;
	andOp #(.WIDTH(1)) andOp_580(.in0(andOp_580_in0), .in1(andOp_580_in1), .out(andOp_580_out));

	reg [31:0] eq_581_in0;
	reg [31:0] eq_581_in1;
	wire [0:0] eq_581_out;
	eq #(.WIDTH(32)) eq_581(.in0(eq_581_in0), .in1(eq_581_in1), .out(eq_581_out));

	reg [0:0] andOp_582_in0;
	reg [0:0] andOp_582_in1;
	wire [0:0] andOp_582_out;
	andOp #(.WIDTH(1)) andOp_582(.in0(andOp_582_in0), .in1(andOp_582_in1), .out(andOp_582_out));

	reg [0:0] notOp_583_in0;
	wire [0:0] notOp_583_out;
	notOp #(.WIDTH(1)) notOp_583(.in(notOp_583_in0), .out(notOp_583_out));

	reg [0:0] andOp_584_in0;
	reg [0:0] andOp_584_in1;
	wire [0:0] andOp_584_out;
	andOp #(.WIDTH(1)) andOp_584(.in0(andOp_584_in0), .in1(andOp_584_in1), .out(andOp_584_out));

	reg [0:0] notOp_585_in0;
	wire [0:0] notOp_585_out;
	notOp #(.WIDTH(1)) notOp_585(.in(notOp_585_in0), .out(notOp_585_out));

	reg [0:0] andOp_586_in0;
	reg [0:0] andOp_586_in1;
	wire [0:0] andOp_586_out;
	andOp #(.WIDTH(1)) andOp_586(.in0(andOp_586_in0), .in1(andOp_586_in1), .out(andOp_586_out));

	reg [0:0] notOp_587_in0;
	wire [0:0] notOp_587_out;
	notOp #(.WIDTH(1)) notOp_587(.in(notOp_587_in0), .out(notOp_587_out));

	reg [0:0] andOp_588_in0;
	reg [0:0] andOp_588_in1;
	wire [0:0] andOp_588_out;
	andOp #(.WIDTH(1)) andOp_588(.in0(andOp_588_in0), .in1(andOp_588_in1), .out(andOp_588_out));

	reg [0:0] andOp_589_in0;
	reg [0:0] andOp_589_in1;
	wire [0:0] andOp_589_out;
	andOp #(.WIDTH(1)) andOp_589(.in0(andOp_589_in0), .in1(andOp_589_in1), .out(andOp_589_out));

	reg [31:0] eq_590_in0;
	reg [31:0] eq_590_in1;
	wire [0:0] eq_590_out;
	eq #(.WIDTH(32)) eq_590(.in0(eq_590_in0), .in1(eq_590_in1), .out(eq_590_out));

	reg [0:0] andOp_591_in0;
	reg [0:0] andOp_591_in1;
	wire [0:0] andOp_591_out;
	andOp #(.WIDTH(1)) andOp_591(.in0(andOp_591_in0), .in1(andOp_591_in1), .out(andOp_591_out));

	reg [0:0] notOp_592_in0;
	wire [0:0] notOp_592_out;
	notOp #(.WIDTH(1)) notOp_592(.in(notOp_592_in0), .out(notOp_592_out));

	reg [0:0] andOp_593_in0;
	reg [0:0] andOp_593_in1;
	wire [0:0] andOp_593_out;
	andOp #(.WIDTH(1)) andOp_593(.in0(andOp_593_in0), .in1(andOp_593_in1), .out(andOp_593_out));

	reg [0:0] notOp_594_in0;
	wire [0:0] notOp_594_out;
	notOp #(.WIDTH(1)) notOp_594(.in(notOp_594_in0), .out(notOp_594_out));

	reg [0:0] andOp_595_in0;
	reg [0:0] andOp_595_in1;
	wire [0:0] andOp_595_out;
	andOp #(.WIDTH(1)) andOp_595(.in0(andOp_595_in0), .in1(andOp_595_in1), .out(andOp_595_out));

	reg [0:0] notOp_596_in0;
	wire [0:0] notOp_596_out;
	notOp #(.WIDTH(1)) notOp_596(.in(notOp_596_in0), .out(notOp_596_out));

	reg [0:0] andOp_597_in0;
	reg [0:0] andOp_597_in1;
	wire [0:0] andOp_597_out;
	andOp #(.WIDTH(1)) andOp_597(.in0(andOp_597_in0), .in1(andOp_597_in1), .out(andOp_597_out));

	reg [0:0] andOp_598_in0;
	reg [0:0] andOp_598_in1;
	wire [0:0] andOp_598_out;
	andOp #(.WIDTH(1)) andOp_598(.in0(andOp_598_in0), .in1(andOp_598_in1), .out(andOp_598_out));

	reg [31:0] eq_599_in0;
	reg [31:0] eq_599_in1;
	wire [0:0] eq_599_out;
	eq #(.WIDTH(32)) eq_599(.in0(eq_599_in0), .in1(eq_599_in1), .out(eq_599_out));

	reg [0:0] andOp_600_in0;
	reg [0:0] andOp_600_in1;
	wire [0:0] andOp_600_out;
	andOp #(.WIDTH(1)) andOp_600(.in0(andOp_600_in0), .in1(andOp_600_in1), .out(andOp_600_out));

	reg [0:0] notOp_601_in0;
	wire [0:0] notOp_601_out;
	notOp #(.WIDTH(1)) notOp_601(.in(notOp_601_in0), .out(notOp_601_out));

	reg [0:0] andOp_602_in0;
	reg [0:0] andOp_602_in1;
	wire [0:0] andOp_602_out;
	andOp #(.WIDTH(1)) andOp_602(.in0(andOp_602_in0), .in1(andOp_602_in1), .out(andOp_602_out));

	reg [0:0] notOp_603_in0;
	wire [0:0] notOp_603_out;
	notOp #(.WIDTH(1)) notOp_603(.in(notOp_603_in0), .out(notOp_603_out));

	reg [0:0] andOp_604_in0;
	reg [0:0] andOp_604_in1;
	wire [0:0] andOp_604_out;
	andOp #(.WIDTH(1)) andOp_604(.in0(andOp_604_in0), .in1(andOp_604_in1), .out(andOp_604_out));

	reg [0:0] notOp_605_in0;
	wire [0:0] notOp_605_out;
	notOp #(.WIDTH(1)) notOp_605(.in(notOp_605_in0), .out(notOp_605_out));

	reg [0:0] andOp_606_in0;
	reg [0:0] andOp_606_in1;
	wire [0:0] andOp_606_out;
	andOp #(.WIDTH(1)) andOp_606(.in0(andOp_606_in0), .in1(andOp_606_in1), .out(andOp_606_out));

	reg [31:0] eq_607_in0;
	reg [31:0] eq_607_in1;
	wire [0:0] eq_607_out;
	eq #(.WIDTH(32)) eq_607(.in0(eq_607_in0), .in1(eq_607_in1), .out(eq_607_out));

	reg [0:0] andOp_608_in0;
	reg [0:0] andOp_608_in1;
	wire [0:0] andOp_608_out;
	andOp #(.WIDTH(1)) andOp_608(.in0(andOp_608_in0), .in1(andOp_608_in1), .out(andOp_608_out));

	reg [31:0] eq_609_in0;
	reg [31:0] eq_609_in1;
	wire [0:0] eq_609_out;
	eq #(.WIDTH(32)) eq_609(.in0(eq_609_in0), .in1(eq_609_in1), .out(eq_609_out));

	reg [0:0] andOp_610_in0;
	reg [0:0] andOp_610_in1;
	wire [0:0] andOp_610_out;
	andOp #(.WIDTH(1)) andOp_610(.in0(andOp_610_in0), .in1(andOp_610_in1), .out(andOp_610_out));

	reg [31:0] eq_611_in0;
	reg [31:0] eq_611_in1;
	wire [0:0] eq_611_out;
	eq #(.WIDTH(32)) eq_611(.in0(eq_611_in0), .in1(eq_611_in1), .out(eq_611_out));

	reg [0:0] andOp_612_in0;
	reg [0:0] andOp_612_in1;
	wire [0:0] andOp_612_out;
	andOp #(.WIDTH(1)) andOp_612(.in0(andOp_612_in0), .in1(andOp_612_in1), .out(andOp_612_out));

	reg [31:0] eq_613_in0;
	reg [31:0] eq_613_in1;
	wire [0:0] eq_613_out;
	eq #(.WIDTH(32)) eq_613(.in0(eq_613_in0), .in1(eq_613_in1), .out(eq_613_out));

	reg [0:0] andOp_614_in0;
	reg [0:0] andOp_614_in1;
	wire [0:0] andOp_614_out;
	andOp #(.WIDTH(1)) andOp_614(.in0(andOp_614_in0), .in1(andOp_614_in1), .out(andOp_614_out));

	reg [31:0] eq_615_in0;
	reg [31:0] eq_615_in1;
	wire [0:0] eq_615_out;
	eq #(.WIDTH(32)) eq_615(.in0(eq_615_in0), .in1(eq_615_in1), .out(eq_615_out));

	reg [0:0] andOp_616_in0;
	reg [0:0] andOp_616_in1;
	wire [0:0] andOp_616_out;
	andOp #(.WIDTH(1)) andOp_616(.in0(andOp_616_in0), .in1(andOp_616_in1), .out(andOp_616_out));

	reg [0:0] andOp_617_in0;
	reg [0:0] andOp_617_in1;
	wire [0:0] andOp_617_out;
	andOp #(.WIDTH(1)) andOp_617(.in0(andOp_617_in0), .in1(andOp_617_in1), .out(andOp_617_out));

	reg [31:0] eq_618_in0;
	reg [31:0] eq_618_in1;
	wire [0:0] eq_618_out;
	eq #(.WIDTH(32)) eq_618(.in0(eq_618_in0), .in1(eq_618_in1), .out(eq_618_out));

	reg [0:0] andOp_619_in0;
	reg [0:0] andOp_619_in1;
	wire [0:0] andOp_619_out;
	andOp #(.WIDTH(1)) andOp_619(.in0(andOp_619_in0), .in1(andOp_619_in1), .out(andOp_619_out));

	reg [0:0] notOp_620_in0;
	wire [0:0] notOp_620_out;
	notOp #(.WIDTH(1)) notOp_620(.in(notOp_620_in0), .out(notOp_620_out));

	reg [0:0] andOp_621_in0;
	reg [0:0] andOp_621_in1;
	wire [0:0] andOp_621_out;
	andOp #(.WIDTH(1)) andOp_621(.in0(andOp_621_in0), .in1(andOp_621_in1), .out(andOp_621_out));

	reg [0:0] notOp_622_in0;
	wire [0:0] notOp_622_out;
	notOp #(.WIDTH(1)) notOp_622(.in(notOp_622_in0), .out(notOp_622_out));

	reg [0:0] andOp_623_in0;
	reg [0:0] andOp_623_in1;
	wire [0:0] andOp_623_out;
	andOp #(.WIDTH(1)) andOp_623(.in0(andOp_623_in0), .in1(andOp_623_in1), .out(andOp_623_out));

	reg [0:0] notOp_624_in0;
	wire [0:0] notOp_624_out;
	notOp #(.WIDTH(1)) notOp_624(.in(notOp_624_in0), .out(notOp_624_out));

	reg [0:0] andOp_625_in0;
	reg [0:0] andOp_625_in1;
	wire [0:0] andOp_625_out;
	andOp #(.WIDTH(1)) andOp_625(.in0(andOp_625_in0), .in1(andOp_625_in1), .out(andOp_625_out));

	reg [0:0] andOp_626_in0;
	reg [0:0] andOp_626_in1;
	wire [0:0] andOp_626_out;
	andOp #(.WIDTH(1)) andOp_626(.in0(andOp_626_in0), .in1(andOp_626_in1), .out(andOp_626_out));

	reg [31:0] eq_627_in0;
	reg [31:0] eq_627_in1;
	wire [0:0] eq_627_out;
	eq #(.WIDTH(32)) eq_627(.in0(eq_627_in0), .in1(eq_627_in1), .out(eq_627_out));

	reg [0:0] andOp_628_in0;
	reg [0:0] andOp_628_in1;
	wire [0:0] andOp_628_out;
	andOp #(.WIDTH(1)) andOp_628(.in0(andOp_628_in0), .in1(andOp_628_in1), .out(andOp_628_out));

	reg [0:0] notOp_629_in0;
	wire [0:0] notOp_629_out;
	notOp #(.WIDTH(1)) notOp_629(.in(notOp_629_in0), .out(notOp_629_out));

	reg [0:0] andOp_630_in0;
	reg [0:0] andOp_630_in1;
	wire [0:0] andOp_630_out;
	andOp #(.WIDTH(1)) andOp_630(.in0(andOp_630_in0), .in1(andOp_630_in1), .out(andOp_630_out));

	reg [0:0] notOp_631_in0;
	wire [0:0] notOp_631_out;
	notOp #(.WIDTH(1)) notOp_631(.in(notOp_631_in0), .out(notOp_631_out));

	reg [0:0] andOp_632_in0;
	reg [0:0] andOp_632_in1;
	wire [0:0] andOp_632_out;
	andOp #(.WIDTH(1)) andOp_632(.in0(andOp_632_in0), .in1(andOp_632_in1), .out(andOp_632_out));

	reg [0:0] notOp_633_in0;
	wire [0:0] notOp_633_out;
	notOp #(.WIDTH(1)) notOp_633(.in(notOp_633_in0), .out(notOp_633_out));

	reg [0:0] andOp_634_in0;
	reg [0:0] andOp_634_in1;
	wire [0:0] andOp_634_out;
	andOp #(.WIDTH(1)) andOp_634(.in0(andOp_634_in0), .in1(andOp_634_in1), .out(andOp_634_out));

	reg [0:0] andOp_635_in0;
	reg [0:0] andOp_635_in1;
	wire [0:0] andOp_635_out;
	andOp #(.WIDTH(1)) andOp_635(.in0(andOp_635_in0), .in1(andOp_635_in1), .out(andOp_635_out));

	reg [31:0] eq_636_in0;
	reg [31:0] eq_636_in1;
	wire [0:0] eq_636_out;
	eq #(.WIDTH(32)) eq_636(.in0(eq_636_in0), .in1(eq_636_in1), .out(eq_636_out));

	reg [0:0] andOp_637_in0;
	reg [0:0] andOp_637_in1;
	wire [0:0] andOp_637_out;
	andOp #(.WIDTH(1)) andOp_637(.in0(andOp_637_in0), .in1(andOp_637_in1), .out(andOp_637_out));

	reg [0:0] notOp_638_in0;
	wire [0:0] notOp_638_out;
	notOp #(.WIDTH(1)) notOp_638(.in(notOp_638_in0), .out(notOp_638_out));

	reg [0:0] andOp_639_in0;
	reg [0:0] andOp_639_in1;
	wire [0:0] andOp_639_out;
	andOp #(.WIDTH(1)) andOp_639(.in0(andOp_639_in0), .in1(andOp_639_in1), .out(andOp_639_out));

	reg [0:0] notOp_640_in0;
	wire [0:0] notOp_640_out;
	notOp #(.WIDTH(1)) notOp_640(.in(notOp_640_in0), .out(notOp_640_out));

	reg [0:0] andOp_641_in0;
	reg [0:0] andOp_641_in1;
	wire [0:0] andOp_641_out;
	andOp #(.WIDTH(1)) andOp_641(.in0(andOp_641_in0), .in1(andOp_641_in1), .out(andOp_641_out));

	reg [0:0] notOp_642_in0;
	wire [0:0] notOp_642_out;
	notOp #(.WIDTH(1)) notOp_642(.in(notOp_642_in0), .out(notOp_642_out));

	reg [0:0] andOp_643_in0;
	reg [0:0] andOp_643_in1;
	wire [0:0] andOp_643_out;
	andOp #(.WIDTH(1)) andOp_643(.in0(andOp_643_in0), .in1(andOp_643_in1), .out(andOp_643_out));

	reg [0:0] andOp_644_in0;
	reg [0:0] andOp_644_in1;
	wire [0:0] andOp_644_out;
	andOp #(.WIDTH(1)) andOp_644(.in0(andOp_644_in0), .in1(andOp_644_in1), .out(andOp_644_out));

	reg [31:0] eq_645_in0;
	reg [31:0] eq_645_in1;
	wire [0:0] eq_645_out;
	eq #(.WIDTH(32)) eq_645(.in0(eq_645_in0), .in1(eq_645_in1), .out(eq_645_out));

	reg [0:0] andOp_646_in0;
	reg [0:0] andOp_646_in1;
	wire [0:0] andOp_646_out;
	andOp #(.WIDTH(1)) andOp_646(.in0(andOp_646_in0), .in1(andOp_646_in1), .out(andOp_646_out));

	reg [0:0] notOp_647_in0;
	wire [0:0] notOp_647_out;
	notOp #(.WIDTH(1)) notOp_647(.in(notOp_647_in0), .out(notOp_647_out));

	reg [0:0] andOp_648_in0;
	reg [0:0] andOp_648_in1;
	wire [0:0] andOp_648_out;
	andOp #(.WIDTH(1)) andOp_648(.in0(andOp_648_in0), .in1(andOp_648_in1), .out(andOp_648_out));

	reg [0:0] notOp_649_in0;
	wire [0:0] notOp_649_out;
	notOp #(.WIDTH(1)) notOp_649(.in(notOp_649_in0), .out(notOp_649_out));

	reg [0:0] andOp_650_in0;
	reg [0:0] andOp_650_in1;
	wire [0:0] andOp_650_out;
	andOp #(.WIDTH(1)) andOp_650(.in0(andOp_650_in0), .in1(andOp_650_in1), .out(andOp_650_out));

	reg [0:0] notOp_651_in0;
	wire [0:0] notOp_651_out;
	notOp #(.WIDTH(1)) notOp_651(.in(notOp_651_in0), .out(notOp_651_out));

	reg [0:0] andOp_652_in0;
	reg [0:0] andOp_652_in1;
	wire [0:0] andOp_652_out;
	andOp #(.WIDTH(1)) andOp_652(.in0(andOp_652_in0), .in1(andOp_652_in1), .out(andOp_652_out));

	reg [0:0] andOp_653_in0;
	reg [0:0] andOp_653_in1;
	wire [0:0] andOp_653_out;
	andOp #(.WIDTH(1)) andOp_653(.in0(andOp_653_in0), .in1(andOp_653_in1), .out(andOp_653_out));

	reg [31:0] eq_654_in0;
	reg [31:0] eq_654_in1;
	wire [0:0] eq_654_out;
	eq #(.WIDTH(32)) eq_654(.in0(eq_654_in0), .in1(eq_654_in1), .out(eq_654_out));

	reg [0:0] andOp_655_in0;
	reg [0:0] andOp_655_in1;
	wire [0:0] andOp_655_out;
	andOp #(.WIDTH(1)) andOp_655(.in0(andOp_655_in0), .in1(andOp_655_in1), .out(andOp_655_out));

	reg [0:0] notOp_656_in0;
	wire [0:0] notOp_656_out;
	notOp #(.WIDTH(1)) notOp_656(.in(notOp_656_in0), .out(notOp_656_out));

	reg [0:0] andOp_657_in0;
	reg [0:0] andOp_657_in1;
	wire [0:0] andOp_657_out;
	andOp #(.WIDTH(1)) andOp_657(.in0(andOp_657_in0), .in1(andOp_657_in1), .out(andOp_657_out));

	reg [0:0] notOp_658_in0;
	wire [0:0] notOp_658_out;
	notOp #(.WIDTH(1)) notOp_658(.in(notOp_658_in0), .out(notOp_658_out));

	reg [0:0] andOp_659_in0;
	reg [0:0] andOp_659_in1;
	wire [0:0] andOp_659_out;
	andOp #(.WIDTH(1)) andOp_659(.in0(andOp_659_in0), .in1(andOp_659_in1), .out(andOp_659_out));

	reg [0:0] notOp_660_in0;
	wire [0:0] notOp_660_out;
	notOp #(.WIDTH(1)) notOp_660(.in(notOp_660_in0), .out(notOp_660_out));

	reg [0:0] andOp_661_in0;
	reg [0:0] andOp_661_in1;
	wire [0:0] andOp_661_out;
	andOp #(.WIDTH(1)) andOp_661(.in0(andOp_661_in0), .in1(andOp_661_in1), .out(andOp_661_out));

	reg [0:0] andOp_662_in0;
	reg [0:0] andOp_662_in1;
	wire [0:0] andOp_662_out;
	andOp #(.WIDTH(1)) andOp_662(.in0(andOp_662_in0), .in1(andOp_662_in1), .out(andOp_662_out));

	reg [31:0] eq_663_in0;
	reg [31:0] eq_663_in1;
	wire [0:0] eq_663_out;
	eq #(.WIDTH(32)) eq_663(.in0(eq_663_in0), .in1(eq_663_in1), .out(eq_663_out));

	reg [0:0] andOp_664_in0;
	reg [0:0] andOp_664_in1;
	wire [0:0] andOp_664_out;
	andOp #(.WIDTH(1)) andOp_664(.in0(andOp_664_in0), .in1(andOp_664_in1), .out(andOp_664_out));

	reg [0:0] notOp_665_in0;
	wire [0:0] notOp_665_out;
	notOp #(.WIDTH(1)) notOp_665(.in(notOp_665_in0), .out(notOp_665_out));

	reg [0:0] andOp_666_in0;
	reg [0:0] andOp_666_in1;
	wire [0:0] andOp_666_out;
	andOp #(.WIDTH(1)) andOp_666(.in0(andOp_666_in0), .in1(andOp_666_in1), .out(andOp_666_out));

	reg [0:0] notOp_667_in0;
	wire [0:0] notOp_667_out;
	notOp #(.WIDTH(1)) notOp_667(.in(notOp_667_in0), .out(notOp_667_out));

	reg [0:0] andOp_668_in0;
	reg [0:0] andOp_668_in1;
	wire [0:0] andOp_668_out;
	andOp #(.WIDTH(1)) andOp_668(.in0(andOp_668_in0), .in1(andOp_668_in1), .out(andOp_668_out));

	reg [0:0] notOp_669_in0;
	wire [0:0] notOp_669_out;
	notOp #(.WIDTH(1)) notOp_669(.in(notOp_669_in0), .out(notOp_669_out));

	reg [0:0] andOp_670_in0;
	reg [0:0] andOp_670_in1;
	wire [0:0] andOp_670_out;
	andOp #(.WIDTH(1)) andOp_670(.in0(andOp_670_in0), .in1(andOp_670_in1), .out(andOp_670_out));

	reg [0:0] andOp_671_in0;
	reg [0:0] andOp_671_in1;
	wire [0:0] andOp_671_out;
	andOp #(.WIDTH(1)) andOp_671(.in0(andOp_671_in0), .in1(andOp_671_in1), .out(andOp_671_out));

	reg [31:0] eq_672_in0;
	reg [31:0] eq_672_in1;
	wire [0:0] eq_672_out;
	eq #(.WIDTH(32)) eq_672(.in0(eq_672_in0), .in1(eq_672_in1), .out(eq_672_out));

	reg [0:0] andOp_673_in0;
	reg [0:0] andOp_673_in1;
	wire [0:0] andOp_673_out;
	andOp #(.WIDTH(1)) andOp_673(.in0(andOp_673_in0), .in1(andOp_673_in1), .out(andOp_673_out));

	reg [0:0] notOp_674_in0;
	wire [0:0] notOp_674_out;
	notOp #(.WIDTH(1)) notOp_674(.in(notOp_674_in0), .out(notOp_674_out));

	reg [0:0] andOp_675_in0;
	reg [0:0] andOp_675_in1;
	wire [0:0] andOp_675_out;
	andOp #(.WIDTH(1)) andOp_675(.in0(andOp_675_in0), .in1(andOp_675_in1), .out(andOp_675_out));

	reg [0:0] notOp_676_in0;
	wire [0:0] notOp_676_out;
	notOp #(.WIDTH(1)) notOp_676(.in(notOp_676_in0), .out(notOp_676_out));

	reg [0:0] andOp_677_in0;
	reg [0:0] andOp_677_in1;
	wire [0:0] andOp_677_out;
	andOp #(.WIDTH(1)) andOp_677(.in0(andOp_677_in0), .in1(andOp_677_in1), .out(andOp_677_out));

	reg [0:0] notOp_678_in0;
	wire [0:0] notOp_678_out;
	notOp #(.WIDTH(1)) notOp_678(.in(notOp_678_in0), .out(notOp_678_out));

	reg [0:0] andOp_679_in0;
	reg [0:0] andOp_679_in1;
	wire [0:0] andOp_679_out;
	andOp #(.WIDTH(1)) andOp_679(.in0(andOp_679_in0), .in1(andOp_679_in1), .out(andOp_679_out));

	reg [0:0] andOp_680_in0;
	reg [0:0] andOp_680_in1;
	wire [0:0] andOp_680_out;
	andOp #(.WIDTH(1)) andOp_680(.in0(andOp_680_in0), .in1(andOp_680_in1), .out(andOp_680_out));

	reg [31:0] eq_681_in0;
	reg [31:0] eq_681_in1;
	wire [0:0] eq_681_out;
	eq #(.WIDTH(32)) eq_681(.in0(eq_681_in0), .in1(eq_681_in1), .out(eq_681_out));

	reg [0:0] andOp_682_in0;
	reg [0:0] andOp_682_in1;
	wire [0:0] andOp_682_out;
	andOp #(.WIDTH(1)) andOp_682(.in0(andOp_682_in0), .in1(andOp_682_in1), .out(andOp_682_out));

	reg [0:0] notOp_683_in0;
	wire [0:0] notOp_683_out;
	notOp #(.WIDTH(1)) notOp_683(.in(notOp_683_in0), .out(notOp_683_out));

	reg [0:0] andOp_684_in0;
	reg [0:0] andOp_684_in1;
	wire [0:0] andOp_684_out;
	andOp #(.WIDTH(1)) andOp_684(.in0(andOp_684_in0), .in1(andOp_684_in1), .out(andOp_684_out));

	reg [0:0] notOp_685_in0;
	wire [0:0] notOp_685_out;
	notOp #(.WIDTH(1)) notOp_685(.in(notOp_685_in0), .out(notOp_685_out));

	reg [0:0] andOp_686_in0;
	reg [0:0] andOp_686_in1;
	wire [0:0] andOp_686_out;
	andOp #(.WIDTH(1)) andOp_686(.in0(andOp_686_in0), .in1(andOp_686_in1), .out(andOp_686_out));

	reg [0:0] notOp_687_in0;
	wire [0:0] notOp_687_out;
	notOp #(.WIDTH(1)) notOp_687(.in(notOp_687_in0), .out(notOp_687_out));

	reg [0:0] andOp_688_in0;
	reg [0:0] andOp_688_in1;
	wire [0:0] andOp_688_out;
	andOp #(.WIDTH(1)) andOp_688(.in0(andOp_688_in0), .in1(andOp_688_in1), .out(andOp_688_out));

	reg [0:0] andOp_689_in0;
	reg [0:0] andOp_689_in1;
	wire [0:0] andOp_689_out;
	andOp #(.WIDTH(1)) andOp_689(.in0(andOp_689_in0), .in1(andOp_689_in1), .out(andOp_689_out));

	reg [31:0] eq_690_in0;
	reg [31:0] eq_690_in1;
	wire [0:0] eq_690_out;
	eq #(.WIDTH(32)) eq_690(.in0(eq_690_in0), .in1(eq_690_in1), .out(eq_690_out));

	reg [0:0] andOp_691_in0;
	reg [0:0] andOp_691_in1;
	wire [0:0] andOp_691_out;
	andOp #(.WIDTH(1)) andOp_691(.in0(andOp_691_in0), .in1(andOp_691_in1), .out(andOp_691_out));

	reg [0:0] notOp_692_in0;
	wire [0:0] notOp_692_out;
	notOp #(.WIDTH(1)) notOp_692(.in(notOp_692_in0), .out(notOp_692_out));

	reg [0:0] andOp_693_in0;
	reg [0:0] andOp_693_in1;
	wire [0:0] andOp_693_out;
	andOp #(.WIDTH(1)) andOp_693(.in0(andOp_693_in0), .in1(andOp_693_in1), .out(andOp_693_out));

	reg [0:0] notOp_694_in0;
	wire [0:0] notOp_694_out;
	notOp #(.WIDTH(1)) notOp_694(.in(notOp_694_in0), .out(notOp_694_out));

	reg [0:0] andOp_695_in0;
	reg [0:0] andOp_695_in1;
	wire [0:0] andOp_695_out;
	andOp #(.WIDTH(1)) andOp_695(.in0(andOp_695_in0), .in1(andOp_695_in1), .out(andOp_695_out));

	reg [0:0] notOp_696_in0;
	wire [0:0] notOp_696_out;
	notOp #(.WIDTH(1)) notOp_696(.in(notOp_696_in0), .out(notOp_696_out));

	reg [0:0] andOp_697_in0;
	reg [0:0] andOp_697_in1;
	wire [0:0] andOp_697_out;
	andOp #(.WIDTH(1)) andOp_697(.in0(andOp_697_in0), .in1(andOp_697_in1), .out(andOp_697_out));

	// End Functional Units

	reg [31:0] add_tmp_5;
	reg [31:0] call_tmp_2;
	reg [0:0] data_store_0_0;
	reg [31:0] data_store_0_10;
	reg [0:0] data_store_0_12;
	reg [31:0] data_store_0_14;
	reg [0:0] data_store_0_16;
	reg [31:0] data_store_0_2;
	reg [31:0] data_store_0_4;
	reg [31:0] data_store_0_6;
	reg [31:0] data_store_0_8;
	reg [0:0] data_store_1_18;
	reg [31:0] data_store_1_20;
	reg [31:0] data_store_1_22;
	reg [31:0] data_store_1_24;
	reg [31:0] data_store_1_26;
	reg [31:0] data_store_1_28;
	reg [0:0] data_store_1_30;
	reg [31:0] data_store_1_32;
	reg [0:0] data_store_1_34;
	reg [0:0] data_store_2_36;
	reg [31:0] data_store_2_38;
	reg [31:0] data_store_2_40;
	reg [31:0] data_store_2_42;
	reg [31:0] data_store_2_44;
	reg [31:0] data_store_2_46;
	reg [0:0] data_store_2_48;
	reg [31:0] data_store_2_50;
	reg [0:0] data_store_2_52;
	reg [0:0] data_store_3_54;
	reg [31:0] data_store_3_56;
	reg [31:0] data_store_3_58;
	reg [31:0] data_store_3_60;
	reg [31:0] data_store_3_62;
	reg [31:0] data_store_3_64;
	reg [0:0] data_store_3_66;
	reg [31:0] data_store_3_68;
	reg [0:0] data_store_3_70;
	reg [0:0] data_store_4_72;
	reg [31:0] data_store_4_74;
	reg [31:0] data_store_4_76;
	reg [31:0] data_store_4_78;
	reg [31:0] data_store_4_80;
	reg [31:0] data_store_4_82;
	reg [0:0] data_store_4_84;
	reg [31:0] data_store_4_86;
	reg [0:0] data_store_4_88;
	reg [31:0] global_state;
	reg [0:0] icmp_tmp_6;
	reg [31:0] phi_tmp_1;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_3_last_state;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;
	reg [31:0] state_4_last_state;

	// controller for add_add_14.add_in0_add_14
	// controller for add_add_14.add_in1_add_14
	// Insensitive connections
	always @(*) begin
		add_in0_add_14 = valid ? rdata_ram_0 : rdata_ram_0;
		add_in1_add_14 = valid ? tmp_output_210_out_data : tmp_output_210_out_data;
	end
	// controller for add_add_16.add_in0_add_16
	// controller for add_add_16.add_in1_add_16
	// Insensitive connections
	always @(*) begin
		add_in0_add_16 = valid ? data_in_3_59_out_data : data_in_3_59_out_data;
		add_in1_add_16 = valid ? 32'd1 : 32'd1;
	end
	// controller for andOp_100.andOp_100_in0
	// controller for andOp_100.andOp_100_in1
	// Insensitive connections
	always @(*) begin
		andOp_100_in0 = valid ? andOp_99_out : andOp_99_out;
		andOp_100_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_102.andOp_102_in0
	// controller for andOp_102.andOp_102_in1
	// Insensitive connections
	always @(*) begin
		andOp_102_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
		andOp_102_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_103.andOp_103_in0
	// controller for andOp_103.andOp_103_in1
	// Insensitive connections
	always @(*) begin
		andOp_103_in0 = valid ? andOp_102_out : andOp_102_out;
		andOp_103_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_105.andOp_105_in0
	// controller for andOp_105.andOp_105_in1
	// Insensitive connections
	always @(*) begin
		andOp_105_in0 = valid ? andOp_103_out : andOp_103_out;
		andOp_105_in1 = valid ? in_read_ready : in_read_ready;
	end
	// controller for andOp_107.andOp_107_in0
	// controller for andOp_107.andOp_107_in1
	// Insensitive connections
	always @(*) begin
		andOp_107_in0 = valid ? andOp_103_out : andOp_103_out;
		andOp_107_in1 = valid ? notOp_106_out : notOp_106_out;
	end
	// controller for andOp_108.andOp_108_in0
	// controller for andOp_108.andOp_108_in1
	// Insensitive connections
	always @(*) begin
		andOp_108_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_108_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_109.andOp_109_in0
	// controller for andOp_109.andOp_109_in1
	// Insensitive connections
	always @(*) begin
		andOp_109_in0 = valid ? andOp_108_out : andOp_108_out;
		andOp_109_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_111.andOp_111_in0
	// controller for andOp_111.andOp_111_in1
	// Insensitive connections
	always @(*) begin
		andOp_111_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_111_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_112.andOp_112_in0
	// controller for andOp_112.andOp_112_in1
	// Insensitive connections
	always @(*) begin
		andOp_112_in0 = valid ? andOp_111_out : andOp_111_out;
		andOp_112_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_114.andOp_114_in0
	// controller for andOp_114.andOp_114_in1
	// Insensitive connections
	always @(*) begin
		andOp_114_in0 = valid ? andOp_112_out : andOp_112_out;
		andOp_114_in1 = valid ? data_in_4_85_out_data : data_in_4_85_out_data;
	end
	// controller for andOp_116.andOp_116_in0
	// controller for andOp_116.andOp_116_in1
	// Insensitive connections
	always @(*) begin
		andOp_116_in0 = valid ? andOp_112_out : andOp_112_out;
		andOp_116_in1 = valid ? notOp_115_out : notOp_115_out;
	end
	// controller for andOp_117.andOp_117_in0
	// controller for andOp_117.andOp_117_in1
	// Insensitive connections
	always @(*) begin
		andOp_117_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_117_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_118.andOp_118_in0
	// controller for andOp_118.andOp_118_in1
	// Insensitive connections
	always @(*) begin
		andOp_118_in0 = valid ? andOp_117_out : andOp_117_out;
		andOp_118_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_120.andOp_120_in0
	// controller for andOp_120.andOp_120_in1
	// Insensitive connections
	always @(*) begin
		andOp_120_in0 = valid ? bb_5_active_in_state_4_out_data : bb_5_active_in_state_4_out_data;
		andOp_120_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_121.andOp_121_in0
	// controller for andOp_121.andOp_121_in1
	// Insensitive connections
	always @(*) begin
		andOp_121_in0 = valid ? andOp_120_out : andOp_120_out;
		andOp_121_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_123.andOp_123_in0
	// controller for andOp_123.andOp_123_in1
	// Insensitive connections
	always @(*) begin
		andOp_123_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
		andOp_123_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_124.andOp_124_in0
	// controller for andOp_124.andOp_124_in1
	// Insensitive connections
	always @(*) begin
		andOp_124_in0 = valid ? andOp_123_out : andOp_123_out;
		andOp_124_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_126.andOp_126_in0
	// controller for andOp_126.andOp_126_in1
	// Insensitive connections
	always @(*) begin
		andOp_126_in0 = valid ? andOp_124_out : andOp_124_out;
		andOp_126_in1 = valid ? out_write_ready : out_write_ready;
	end
	// controller for andOp_128.andOp_128_in0
	// controller for andOp_128.andOp_128_in1
	// Insensitive connections
	always @(*) begin
		andOp_128_in0 = valid ? andOp_124_out : andOp_124_out;
		andOp_128_in1 = valid ? notOp_127_out : notOp_127_out;
	end
	// controller for andOp_129.andOp_129_in0
	// controller for andOp_129.andOp_129_in1
	// Insensitive connections
	always @(*) begin
		andOp_129_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_129_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_130.andOp_130_in0
	// controller for andOp_130.andOp_130_in1
	// Insensitive connections
	always @(*) begin
		andOp_130_in0 = valid ? andOp_129_out : andOp_129_out;
		andOp_130_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_132.andOp_132_in0
	// controller for andOp_132.andOp_132_in1
	// Insensitive connections
	always @(*) begin
		andOp_132_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_132_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_133.andOp_133_in0
	// controller for andOp_133.andOp_133_in1
	// Insensitive connections
	always @(*) begin
		andOp_133_in0 = valid ? andOp_132_out : andOp_132_out;
		andOp_133_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_135.andOp_135_in0
	// controller for andOp_135.andOp_135_in1
	// Insensitive connections
	always @(*) begin
		andOp_135_in0 = valid ? andOp_133_out : andOp_133_out;
		andOp_135_in1 = valid ? data_in_4_85_out_data : data_in_4_85_out_data;
	end
	// controller for andOp_137.andOp_137_in0
	// controller for andOp_137.andOp_137_in1
	// Insensitive connections
	always @(*) begin
		andOp_137_in0 = valid ? andOp_133_out : andOp_133_out;
		andOp_137_in1 = valid ? notOp_136_out : notOp_136_out;
	end
	// controller for andOp_138.andOp_138_in0
	// controller for andOp_138.andOp_138_in1
	// Insensitive connections
	always @(*) begin
		andOp_138_in0 = valid ? bb_1_active_in_state_4_out_data : bb_1_active_in_state_4_out_data;
		andOp_138_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_139.andOp_139_in0
	// controller for andOp_139.andOp_139_in1
	// Insensitive connections
	always @(*) begin
		andOp_139_in0 = valid ? andOp_138_out : andOp_138_out;
		andOp_139_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_167.andOp_167_in0
	// controller for andOp_167.andOp_167_in1
	// Insensitive connections
	always @(*) begin
		andOp_167_in0 = valid ? notOp_166_out : notOp_166_out;
		andOp_167_in1 = valid ? andOp_100_out : andOp_100_out;
	end
	// controller for andOp_171.andOp_171_in0
	// controller for andOp_171.andOp_171_in1
	// Insensitive connections
	always @(*) begin
		andOp_171_in0 = valid ? notOp_170_out : notOp_170_out;
		andOp_171_in1 = valid ? andOp_91_out : andOp_91_out;
	end
	// controller for andOp_174.andOp_174_in0
	// controller for andOp_174.andOp_174_in1
	// Insensitive connections
	always @(*) begin
		andOp_174_in0 = valid ? notOp_173_out : notOp_173_out;
		andOp_174_in1 = valid ? andOp_94_out : andOp_94_out;
	end
	// controller for andOp_178.andOp_178_in0
	// controller for andOp_178.andOp_178_in1
	// Insensitive connections
	always @(*) begin
		andOp_178_in0 = valid ? notOp_177_out : notOp_177_out;
		andOp_178_in1 = valid ? andOp_109_out : andOp_109_out;
	end
	// controller for andOp_182.andOp_182_in0
	// controller for andOp_182.andOp_182_in1
	// Insensitive connections
	always @(*) begin
		andOp_182_in0 = valid ? notOp_181_out : notOp_181_out;
		andOp_182_in1 = valid ? andOp_139_out : andOp_139_out;
	end
	// controller for andOp_185.andOp_185_in0
	// controller for andOp_185.andOp_185_in1
	// Insensitive connections
	always @(*) begin
		andOp_185_in0 = valid ? notOp_184_out : notOp_184_out;
		andOp_185_in1 = valid ? andOp_121_out : andOp_121_out;
	end
	// controller for andOp_188.andOp_188_in0
	// controller for andOp_188.andOp_188_in1
	// Insensitive connections
	always @(*) begin
		andOp_188_in0 = valid ? notOp_187_out : notOp_187_out;
		andOp_188_in1 = valid ? andOp_126_out : andOp_126_out;
	end
	// controller for andOp_192.andOp_192_in0
	// controller for andOp_192.andOp_192_in1
	// Insensitive connections
	always @(*) begin
		andOp_192_in0 = valid ? notOp_191_out : notOp_191_out;
		andOp_192_in1 = valid ? andOp_130_out : andOp_130_out;
	end
	// controller for andOp_195.andOp_195_in0
	// controller for andOp_195.andOp_195_in1
	// Insensitive connections
	always @(*) begin
		andOp_195_in0 = valid ? notOp_194_out : notOp_194_out;
		andOp_195_in1 = valid ? andOp_114_out : andOp_114_out;
	end
	// controller for andOp_196.andOp_196_in0
	// controller for andOp_196.andOp_196_in1
	// Insensitive connections
	always @(*) begin
		andOp_196_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_196_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_197.andOp_197_in0
	// controller for andOp_197.andOp_197_in1
	// Insensitive connections
	always @(*) begin
		andOp_197_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_197_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_198.andOp_198_in0
	// controller for andOp_198.andOp_198_in1
	// Insensitive connections
	always @(*) begin
		andOp_198_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_198_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_199.andOp_199_in0
	// controller for andOp_199.andOp_199_in1
	// Insensitive connections
	always @(*) begin
		andOp_199_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_199_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_200.andOp_200_in0
	// controller for andOp_200.andOp_200_in1
	// Insensitive connections
	always @(*) begin
		andOp_200_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_200_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_201.andOp_201_in0
	// controller for andOp_201.andOp_201_in1
	// Insensitive connections
	always @(*) begin
		andOp_201_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_201_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_202.andOp_202_in0
	// controller for andOp_202.andOp_202_in1
	// Insensitive connections
	always @(*) begin
		andOp_202_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_202_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_203.andOp_203_in0
	// controller for andOp_203.andOp_203_in1
	// Insensitive connections
	always @(*) begin
		andOp_203_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
		andOp_203_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_204.andOp_204_in0
	// controller for andOp_204.andOp_204_in1
	// Insensitive connections
	always @(*) begin
		andOp_204_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_204_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_205.andOp_205_in0
	// controller for andOp_205.andOp_205_in1
	// Insensitive connections
	always @(*) begin
		andOp_205_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_205_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_206.andOp_206_in0
	// controller for andOp_206.andOp_206_in1
	// Insensitive connections
	always @(*) begin
		andOp_206_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_206_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_209.andOp_209_in0
	// controller for andOp_209.andOp_209_in1
	// Insensitive connections
	always @(*) begin
		andOp_209_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_209_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_212.andOp_212_in0
	// controller for andOp_212.andOp_212_in1
	// Insensitive connections
	always @(*) begin
		andOp_212_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_212_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_213.andOp_213_in0
	// controller for andOp_213.andOp_213_in1
	// Insensitive connections
	always @(*) begin
		andOp_213_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_213_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_214.andOp_214_in0
	// controller for andOp_214.andOp_214_in1
	// Insensitive connections
	always @(*) begin
		andOp_214_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_214_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_215.andOp_215_in0
	// controller for andOp_215.andOp_215_in1
	// Insensitive connections
	always @(*) begin
		andOp_215_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_215_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_216.andOp_216_in0
	// controller for andOp_216.andOp_216_in1
	// Insensitive connections
	always @(*) begin
		andOp_216_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
		andOp_216_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_217.andOp_217_in0
	// controller for andOp_217.andOp_217_in1
	// Insensitive connections
	always @(*) begin
		andOp_217_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_217_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_218.andOp_218_in0
	// controller for andOp_218.andOp_218_in1
	// Insensitive connections
	always @(*) begin
		andOp_218_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_218_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_219.andOp_219_in0
	// controller for andOp_219.andOp_219_in1
	// Insensitive connections
	always @(*) begin
		andOp_219_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_219_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_220.andOp_220_in0
	// controller for andOp_220.andOp_220_in1
	// Insensitive connections
	always @(*) begin
		andOp_220_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_220_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_221.andOp_221_in0
	// controller for andOp_221.andOp_221_in1
	// Insensitive connections
	always @(*) begin
		andOp_221_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_221_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_222.andOp_222_in0
	// controller for andOp_222.andOp_222_in1
	// Insensitive connections
	always @(*) begin
		andOp_222_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_222_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_224.andOp_224_in0
	// controller for andOp_224.andOp_224_in1
	// Insensitive connections
	always @(*) begin
		andOp_224_in0 = valid ? notOp_223_out : notOp_223_out;
		andOp_224_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_226.andOp_226_in0
	// controller for andOp_226.andOp_226_in1
	// Insensitive connections
	always @(*) begin
		andOp_226_in0 = valid ? notOp_225_out : notOp_225_out;
		andOp_226_in1 = valid ? andOp_224_out : andOp_224_out;
	end
	// controller for andOp_228.andOp_228_in0
	// controller for andOp_228.andOp_228_in1
	// Insensitive connections
	always @(*) begin
		andOp_228_in0 = valid ? notOp_227_out : notOp_227_out;
		andOp_228_in1 = valid ? andOp_226_out : andOp_226_out;
	end
	// controller for andOp_230.andOp_230_in0
	// controller for andOp_230.andOp_230_in1
	// Insensitive connections
	always @(*) begin
		andOp_230_in0 = valid ? notOp_229_out : notOp_229_out;
		andOp_230_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_232.andOp_232_in0
	// controller for andOp_232.andOp_232_in1
	// Insensitive connections
	always @(*) begin
		andOp_232_in0 = valid ? notOp_231_out : notOp_231_out;
		andOp_232_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_234.andOp_234_in0
	// controller for andOp_234.andOp_234_in1
	// Insensitive connections
	always @(*) begin
		andOp_234_in0 = valid ? notOp_233_out : notOp_233_out;
		andOp_234_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_236.andOp_236_in0
	// controller for andOp_236.andOp_236_in1
	// Insensitive connections
	always @(*) begin
		andOp_236_in0 = valid ? notOp_235_out : notOp_235_out;
		andOp_236_in1 = valid ? andOp_234_out : andOp_234_out;
	end
	// controller for andOp_238.andOp_238_in0
	// controller for andOp_238.andOp_238_in1
	// Insensitive connections
	always @(*) begin
		andOp_238_in0 = valid ? notOp_237_out : notOp_237_out;
		andOp_238_in1 = valid ? andOp_236_out : andOp_236_out;
	end
	// controller for andOp_239.andOp_239_in0
	// controller for andOp_239.andOp_239_in1
	// Insensitive connections
	always @(*) begin
		andOp_239_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_239_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_240.andOp_240_in0
	// controller for andOp_240.andOp_240_in1
	// Insensitive connections
	always @(*) begin
		andOp_240_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_240_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_241.andOp_241_in0
	// controller for andOp_241.andOp_241_in1
	// Insensitive connections
	always @(*) begin
		andOp_241_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_241_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_242.andOp_242_in0
	// controller for andOp_242.andOp_242_in1
	// Insensitive connections
	always @(*) begin
		andOp_242_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_242_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_244.andOp_244_in0
	// controller for andOp_244.andOp_244_in1
	// Insensitive connections
	always @(*) begin
		andOp_244_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_244_in1 = valid ? eq_243_out : eq_243_out;
	end
	// controller for andOp_246.andOp_246_in0
	// controller for andOp_246.andOp_246_in1
	// Insensitive connections
	always @(*) begin
		andOp_246_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_246_in1 = valid ? eq_245_out : eq_245_out;
	end
	// controller for andOp_248.andOp_248_in0
	// controller for andOp_248.andOp_248_in1
	// Insensitive connections
	always @(*) begin
		andOp_248_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_248_in1 = valid ? eq_247_out : eq_247_out;
	end
	// controller for andOp_250.andOp_250_in0
	// controller for andOp_250.andOp_250_in1
	// Insensitive connections
	always @(*) begin
		andOp_250_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_250_in1 = valid ? eq_249_out : eq_249_out;
	end
	// controller for andOp_252.andOp_252_in0
	// controller for andOp_252.andOp_252_in1
	// Insensitive connections
	always @(*) begin
		andOp_252_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_252_in1 = valid ? eq_251_out : eq_251_out;
	end
	// controller for andOp_253.andOp_253_in0
	// controller for andOp_253.andOp_253_in1
	// Insensitive connections
	always @(*) begin
		andOp_253_in0 = valid ? 1'd0 : 1'd0;
		andOp_253_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_255.andOp_255_in0
	// controller for andOp_255.andOp_255_in1
	// Insensitive connections
	always @(*) begin
		andOp_255_in0 = valid ? andOp_253_out : andOp_253_out;
		andOp_255_in1 = valid ? eq_254_out : eq_254_out;
	end
	// controller for andOp_257.andOp_257_in0
	// controller for andOp_257.andOp_257_in1
	// Insensitive connections
	always @(*) begin
		andOp_257_in0 = valid ? andOp_253_out : andOp_253_out;
		andOp_257_in1 = valid ? notOp_256_out : notOp_256_out;
	end
	// controller for andOp_259.andOp_259_in0
	// controller for andOp_259.andOp_259_in1
	// Insensitive connections
	always @(*) begin
		andOp_259_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_259_in1 = valid ? notOp_258_out : notOp_258_out;
	end
	// controller for andOp_261.andOp_261_in0
	// controller for andOp_261.andOp_261_in1
	// Insensitive connections
	always @(*) begin
		andOp_261_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_261_in1 = valid ? notOp_260_out : notOp_260_out;
	end
	// controller for andOp_262.andOp_262_in0
	// controller for andOp_262.andOp_262_in1
	// Insensitive connections
	always @(*) begin
		andOp_262_in0 = valid ? 1'd0 : 1'd0;
		andOp_262_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_264.andOp_264_in0
	// controller for andOp_264.andOp_264_in1
	// Insensitive connections
	always @(*) begin
		andOp_264_in0 = valid ? andOp_262_out : andOp_262_out;
		andOp_264_in1 = valid ? eq_263_out : eq_263_out;
	end
	// controller for andOp_266.andOp_266_in0
	// controller for andOp_266.andOp_266_in1
	// Insensitive connections
	always @(*) begin
		andOp_266_in0 = valid ? andOp_262_out : andOp_262_out;
		andOp_266_in1 = valid ? notOp_265_out : notOp_265_out;
	end
	// controller for andOp_268.andOp_268_in0
	// controller for andOp_268.andOp_268_in1
	// Insensitive connections
	always @(*) begin
		andOp_268_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_268_in1 = valid ? notOp_267_out : notOp_267_out;
	end
	// controller for andOp_270.andOp_270_in0
	// controller for andOp_270.andOp_270_in1
	// Insensitive connections
	always @(*) begin
		andOp_270_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_270_in1 = valid ? notOp_269_out : notOp_269_out;
	end
	// controller for andOp_271.andOp_271_in0
	// controller for andOp_271.andOp_271_in1
	// Insensitive connections
	always @(*) begin
		andOp_271_in0 = valid ? 1'd0 : 1'd0;
		andOp_271_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_273.andOp_273_in0
	// controller for andOp_273.andOp_273_in1
	// Insensitive connections
	always @(*) begin
		andOp_273_in0 = valid ? andOp_271_out : andOp_271_out;
		andOp_273_in1 = valid ? eq_272_out : eq_272_out;
	end
	// controller for andOp_275.andOp_275_in0
	// controller for andOp_275.andOp_275_in1
	// Insensitive connections
	always @(*) begin
		andOp_275_in0 = valid ? andOp_271_out : andOp_271_out;
		andOp_275_in1 = valid ? notOp_274_out : notOp_274_out;
	end
	// controller for andOp_277.andOp_277_in0
	// controller for andOp_277.andOp_277_in1
	// Insensitive connections
	always @(*) begin
		andOp_277_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_277_in1 = valid ? notOp_276_out : notOp_276_out;
	end
	// controller for andOp_279.andOp_279_in0
	// controller for andOp_279.andOp_279_in1
	// Insensitive connections
	always @(*) begin
		andOp_279_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_279_in1 = valid ? notOp_278_out : notOp_278_out;
	end
	// controller for andOp_280.andOp_280_in0
	// controller for andOp_280.andOp_280_in1
	// Insensitive connections
	always @(*) begin
		andOp_280_in0 = valid ? 1'd0 : 1'd0;
		andOp_280_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_282.andOp_282_in0
	// controller for andOp_282.andOp_282_in1
	// Insensitive connections
	always @(*) begin
		andOp_282_in0 = valid ? andOp_280_out : andOp_280_out;
		andOp_282_in1 = valid ? eq_281_out : eq_281_out;
	end
	// controller for andOp_284.andOp_284_in0
	// controller for andOp_284.andOp_284_in1
	// Insensitive connections
	always @(*) begin
		andOp_284_in0 = valid ? andOp_280_out : andOp_280_out;
		andOp_284_in1 = valid ? notOp_283_out : notOp_283_out;
	end
	// controller for andOp_286.andOp_286_in0
	// controller for andOp_286.andOp_286_in1
	// Insensitive connections
	always @(*) begin
		andOp_286_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_286_in1 = valid ? notOp_285_out : notOp_285_out;
	end
	// controller for andOp_288.andOp_288_in0
	// controller for andOp_288.andOp_288_in1
	// Insensitive connections
	always @(*) begin
		andOp_288_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_288_in1 = valid ? notOp_287_out : notOp_287_out;
	end
	// controller for andOp_289.andOp_289_in0
	// controller for andOp_289.andOp_289_in1
	// Insensitive connections
	always @(*) begin
		andOp_289_in0 = valid ? 1'd0 : 1'd0;
		andOp_289_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_291.andOp_291_in0
	// controller for andOp_291.andOp_291_in1
	// Insensitive connections
	always @(*) begin
		andOp_291_in0 = valid ? andOp_289_out : andOp_289_out;
		andOp_291_in1 = valid ? eq_290_out : eq_290_out;
	end
	// controller for andOp_293.andOp_293_in0
	// controller for andOp_293.andOp_293_in1
	// Insensitive connections
	always @(*) begin
		andOp_293_in0 = valid ? andOp_289_out : andOp_289_out;
		andOp_293_in1 = valid ? notOp_292_out : notOp_292_out;
	end
	// controller for andOp_295.andOp_295_in0
	// controller for andOp_295.andOp_295_in1
	// Insensitive connections
	always @(*) begin
		andOp_295_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_295_in1 = valid ? notOp_294_out : notOp_294_out;
	end
	// controller for andOp_297.andOp_297_in0
	// controller for andOp_297.andOp_297_in1
	// Insensitive connections
	always @(*) begin
		andOp_297_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_297_in1 = valid ? notOp_296_out : notOp_296_out;
	end
	// controller for andOp_298.andOp_298_in0
	// controller for andOp_298.andOp_298_in1
	// Insensitive connections
	always @(*) begin
		andOp_298_in0 = valid ? 1'd0 : 1'd0;
		andOp_298_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_300.andOp_300_in0
	// controller for andOp_300.andOp_300_in1
	// Insensitive connections
	always @(*) begin
		andOp_300_in0 = valid ? andOp_298_out : andOp_298_out;
		andOp_300_in1 = valid ? eq_299_out : eq_299_out;
	end
	// controller for andOp_302.andOp_302_in0
	// controller for andOp_302.andOp_302_in1
	// Insensitive connections
	always @(*) begin
		andOp_302_in0 = valid ? andOp_298_out : andOp_298_out;
		andOp_302_in1 = valid ? notOp_301_out : notOp_301_out;
	end
	// controller for andOp_304.andOp_304_in0
	// controller for andOp_304.andOp_304_in1
	// Insensitive connections
	always @(*) begin
		andOp_304_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_304_in1 = valid ? notOp_303_out : notOp_303_out;
	end
	// controller for andOp_306.andOp_306_in0
	// controller for andOp_306.andOp_306_in1
	// Insensitive connections
	always @(*) begin
		andOp_306_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_306_in1 = valid ? notOp_305_out : notOp_305_out;
	end
	// controller for andOp_307.andOp_307_in0
	// controller for andOp_307.andOp_307_in1
	// Insensitive connections
	always @(*) begin
		andOp_307_in0 = valid ? 1'd0 : 1'd0;
		andOp_307_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_309.andOp_309_in0
	// controller for andOp_309.andOp_309_in1
	// Insensitive connections
	always @(*) begin
		andOp_309_in0 = valid ? andOp_307_out : andOp_307_out;
		andOp_309_in1 = valid ? eq_308_out : eq_308_out;
	end
	// controller for andOp_311.andOp_311_in0
	// controller for andOp_311.andOp_311_in1
	// Insensitive connections
	always @(*) begin
		andOp_311_in0 = valid ? andOp_307_out : andOp_307_out;
		andOp_311_in1 = valid ? notOp_310_out : notOp_310_out;
	end
	// controller for andOp_313.andOp_313_in0
	// controller for andOp_313.andOp_313_in1
	// Insensitive connections
	always @(*) begin
		andOp_313_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_313_in1 = valid ? notOp_312_out : notOp_312_out;
	end
	// controller for andOp_315.andOp_315_in0
	// controller for andOp_315.andOp_315_in1
	// Insensitive connections
	always @(*) begin
		andOp_315_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_315_in1 = valid ? notOp_314_out : notOp_314_out;
	end
	// controller for andOp_316.andOp_316_in0
	// controller for andOp_316.andOp_316_in1
	// Insensitive connections
	always @(*) begin
		andOp_316_in0 = valid ? 1'd0 : 1'd0;
		andOp_316_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_318.andOp_318_in0
	// controller for andOp_318.andOp_318_in1
	// Insensitive connections
	always @(*) begin
		andOp_318_in0 = valid ? andOp_316_out : andOp_316_out;
		andOp_318_in1 = valid ? eq_317_out : eq_317_out;
	end
	// controller for andOp_320.andOp_320_in0
	// controller for andOp_320.andOp_320_in1
	// Insensitive connections
	always @(*) begin
		andOp_320_in0 = valid ? andOp_316_out : andOp_316_out;
		andOp_320_in1 = valid ? notOp_319_out : notOp_319_out;
	end
	// controller for andOp_322.andOp_322_in0
	// controller for andOp_322.andOp_322_in1
	// Insensitive connections
	always @(*) begin
		andOp_322_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_322_in1 = valid ? notOp_321_out : notOp_321_out;
	end
	// controller for andOp_324.andOp_324_in0
	// controller for andOp_324.andOp_324_in1
	// Insensitive connections
	always @(*) begin
		andOp_324_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_324_in1 = valid ? notOp_323_out : notOp_323_out;
	end
	// controller for andOp_325.andOp_325_in0
	// controller for andOp_325.andOp_325_in1
	// Insensitive connections
	always @(*) begin
		andOp_325_in0 = valid ? 1'd0 : 1'd0;
		andOp_325_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_327.andOp_327_in0
	// controller for andOp_327.andOp_327_in1
	// Insensitive connections
	always @(*) begin
		andOp_327_in0 = valid ? andOp_325_out : andOp_325_out;
		andOp_327_in1 = valid ? eq_326_out : eq_326_out;
	end
	// controller for andOp_329.andOp_329_in0
	// controller for andOp_329.andOp_329_in1
	// Insensitive connections
	always @(*) begin
		andOp_329_in0 = valid ? andOp_325_out : andOp_325_out;
		andOp_329_in1 = valid ? notOp_328_out : notOp_328_out;
	end
	// controller for andOp_331.andOp_331_in0
	// controller for andOp_331.andOp_331_in1
	// Insensitive connections
	always @(*) begin
		andOp_331_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_331_in1 = valid ? notOp_330_out : notOp_330_out;
	end
	// controller for andOp_333.andOp_333_in0
	// controller for andOp_333.andOp_333_in1
	// Insensitive connections
	always @(*) begin
		andOp_333_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_333_in1 = valid ? notOp_332_out : notOp_332_out;
	end
	// controller for andOp_335.andOp_335_in0
	// controller for andOp_335.andOp_335_in1
	// Insensitive connections
	always @(*) begin
		andOp_335_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_335_in1 = valid ? eq_334_out : eq_334_out;
	end
	// controller for andOp_337.andOp_337_in0
	// controller for andOp_337.andOp_337_in1
	// Insensitive connections
	always @(*) begin
		andOp_337_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_337_in1 = valid ? eq_336_out : eq_336_out;
	end
	// controller for andOp_339.andOp_339_in0
	// controller for andOp_339.andOp_339_in1
	// Insensitive connections
	always @(*) begin
		andOp_339_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_339_in1 = valid ? eq_338_out : eq_338_out;
	end
	// controller for andOp_341.andOp_341_in0
	// controller for andOp_341.andOp_341_in1
	// Insensitive connections
	always @(*) begin
		andOp_341_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_341_in1 = valid ? eq_340_out : eq_340_out;
	end
	// controller for andOp_343.andOp_343_in0
	// controller for andOp_343.andOp_343_in1
	// Insensitive connections
	always @(*) begin
		andOp_343_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_343_in1 = valid ? eq_342_out : eq_342_out;
	end
	// controller for andOp_344.andOp_344_in0
	// controller for andOp_344.andOp_344_in1
	// Insensitive connections
	always @(*) begin
		andOp_344_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
		andOp_344_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_346.andOp_346_in0
	// controller for andOp_346.andOp_346_in1
	// Insensitive connections
	always @(*) begin
		andOp_346_in0 = valid ? andOp_344_out : andOp_344_out;
		andOp_346_in1 = valid ? eq_345_out : eq_345_out;
	end
	// controller for andOp_348.andOp_348_in0
	// controller for andOp_348.andOp_348_in1
	// Insensitive connections
	always @(*) begin
		andOp_348_in0 = valid ? andOp_344_out : andOp_344_out;
		andOp_348_in1 = valid ? notOp_347_out : notOp_347_out;
	end
	// controller for andOp_350.andOp_350_in0
	// controller for andOp_350.andOp_350_in1
	// Insensitive connections
	always @(*) begin
		andOp_350_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_350_in1 = valid ? notOp_349_out : notOp_349_out;
	end
	// controller for andOp_352.andOp_352_in0
	// controller for andOp_352.andOp_352_in1
	// Insensitive connections
	always @(*) begin
		andOp_352_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_352_in1 = valid ? notOp_351_out : notOp_351_out;
	end
	// controller for andOp_353.andOp_353_in0
	// controller for andOp_353.andOp_353_in1
	// Insensitive connections
	always @(*) begin
		andOp_353_in0 = valid ? 1'd0 : 1'd0;
		andOp_353_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_355.andOp_355_in0
	// controller for andOp_355.andOp_355_in1
	// Insensitive connections
	always @(*) begin
		andOp_355_in0 = valid ? andOp_353_out : andOp_353_out;
		andOp_355_in1 = valid ? eq_354_out : eq_354_out;
	end
	// controller for andOp_357.andOp_357_in0
	// controller for andOp_357.andOp_357_in1
	// Insensitive connections
	always @(*) begin
		andOp_357_in0 = valid ? andOp_353_out : andOp_353_out;
		andOp_357_in1 = valid ? notOp_356_out : notOp_356_out;
	end
	// controller for andOp_359.andOp_359_in0
	// controller for andOp_359.andOp_359_in1
	// Insensitive connections
	always @(*) begin
		andOp_359_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_359_in1 = valid ? notOp_358_out : notOp_358_out;
	end
	// controller for andOp_361.andOp_361_in0
	// controller for andOp_361.andOp_361_in1
	// Insensitive connections
	always @(*) begin
		andOp_361_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_361_in1 = valid ? notOp_360_out : notOp_360_out;
	end
	// controller for andOp_362.andOp_362_in0
	// controller for andOp_362.andOp_362_in1
	// Insensitive connections
	always @(*) begin
		andOp_362_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_362_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_364.andOp_364_in0
	// controller for andOp_364.andOp_364_in1
	// Insensitive connections
	always @(*) begin
		andOp_364_in0 = valid ? andOp_362_out : andOp_362_out;
		andOp_364_in1 = valid ? eq_363_out : eq_363_out;
	end
	// controller for andOp_366.andOp_366_in0
	// controller for andOp_366.andOp_366_in1
	// Insensitive connections
	always @(*) begin
		andOp_366_in0 = valid ? andOp_362_out : andOp_362_out;
		andOp_366_in1 = valid ? notOp_365_out : notOp_365_out;
	end
	// controller for andOp_368.andOp_368_in0
	// controller for andOp_368.andOp_368_in1
	// Insensitive connections
	always @(*) begin
		andOp_368_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_368_in1 = valid ? notOp_367_out : notOp_367_out;
	end
	// controller for andOp_370.andOp_370_in0
	// controller for andOp_370.andOp_370_in1
	// Insensitive connections
	always @(*) begin
		andOp_370_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_370_in1 = valid ? notOp_369_out : notOp_369_out;
	end
	// controller for andOp_371.andOp_371_in0
	// controller for andOp_371.andOp_371_in1
	// Insensitive connections
	always @(*) begin
		andOp_371_in0 = valid ? 1'd0 : 1'd0;
		andOp_371_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_373.andOp_373_in0
	// controller for andOp_373.andOp_373_in1
	// Insensitive connections
	always @(*) begin
		andOp_373_in0 = valid ? andOp_371_out : andOp_371_out;
		andOp_373_in1 = valid ? eq_372_out : eq_372_out;
	end
	// controller for andOp_375.andOp_375_in0
	// controller for andOp_375.andOp_375_in1
	// Insensitive connections
	always @(*) begin
		andOp_375_in0 = valid ? andOp_371_out : andOp_371_out;
		andOp_375_in1 = valid ? notOp_374_out : notOp_374_out;
	end
	// controller for andOp_377.andOp_377_in0
	// controller for andOp_377.andOp_377_in1
	// Insensitive connections
	always @(*) begin
		andOp_377_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_377_in1 = valid ? notOp_376_out : notOp_376_out;
	end
	// controller for andOp_379.andOp_379_in0
	// controller for andOp_379.andOp_379_in1
	// Insensitive connections
	always @(*) begin
		andOp_379_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_379_in1 = valid ? notOp_378_out : notOp_378_out;
	end
	// controller for andOp_380.andOp_380_in0
	// controller for andOp_380.andOp_380_in1
	// Insensitive connections
	always @(*) begin
		andOp_380_in0 = valid ? 1'd0 : 1'd0;
		andOp_380_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_382.andOp_382_in0
	// controller for andOp_382.andOp_382_in1
	// Insensitive connections
	always @(*) begin
		andOp_382_in0 = valid ? andOp_380_out : andOp_380_out;
		andOp_382_in1 = valid ? eq_381_out : eq_381_out;
	end
	// controller for andOp_384.andOp_384_in0
	// controller for andOp_384.andOp_384_in1
	// Insensitive connections
	always @(*) begin
		andOp_384_in0 = valid ? andOp_380_out : andOp_380_out;
		andOp_384_in1 = valid ? notOp_383_out : notOp_383_out;
	end
	// controller for andOp_386.andOp_386_in0
	// controller for andOp_386.andOp_386_in1
	// Insensitive connections
	always @(*) begin
		andOp_386_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_386_in1 = valid ? notOp_385_out : notOp_385_out;
	end
	// controller for andOp_388.andOp_388_in0
	// controller for andOp_388.andOp_388_in1
	// Insensitive connections
	always @(*) begin
		andOp_388_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_388_in1 = valid ? notOp_387_out : notOp_387_out;
	end
	// controller for andOp_389.andOp_389_in0
	// controller for andOp_389.andOp_389_in1
	// Insensitive connections
	always @(*) begin
		andOp_389_in0 = valid ? 1'd0 : 1'd0;
		andOp_389_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_391.andOp_391_in0
	// controller for andOp_391.andOp_391_in1
	// Insensitive connections
	always @(*) begin
		andOp_391_in0 = valid ? andOp_389_out : andOp_389_out;
		andOp_391_in1 = valid ? eq_390_out : eq_390_out;
	end
	// controller for andOp_393.andOp_393_in0
	// controller for andOp_393.andOp_393_in1
	// Insensitive connections
	always @(*) begin
		andOp_393_in0 = valid ? andOp_389_out : andOp_389_out;
		andOp_393_in1 = valid ? notOp_392_out : notOp_392_out;
	end
	// controller for andOp_395.andOp_395_in0
	// controller for andOp_395.andOp_395_in1
	// Insensitive connections
	always @(*) begin
		andOp_395_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_395_in1 = valid ? notOp_394_out : notOp_394_out;
	end
	// controller for andOp_397.andOp_397_in0
	// controller for andOp_397.andOp_397_in1
	// Insensitive connections
	always @(*) begin
		andOp_397_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_397_in1 = valid ? notOp_396_out : notOp_396_out;
	end
	// controller for andOp_398.andOp_398_in0
	// controller for andOp_398.andOp_398_in1
	// Insensitive connections
	always @(*) begin
		andOp_398_in0 = valid ? 1'd0 : 1'd0;
		andOp_398_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_400.andOp_400_in0
	// controller for andOp_400.andOp_400_in1
	// Insensitive connections
	always @(*) begin
		andOp_400_in0 = valid ? andOp_398_out : andOp_398_out;
		andOp_400_in1 = valid ? eq_399_out : eq_399_out;
	end
	// controller for andOp_402.andOp_402_in0
	// controller for andOp_402.andOp_402_in1
	// Insensitive connections
	always @(*) begin
		andOp_402_in0 = valid ? andOp_398_out : andOp_398_out;
		andOp_402_in1 = valid ? notOp_401_out : notOp_401_out;
	end
	// controller for andOp_404.andOp_404_in0
	// controller for andOp_404.andOp_404_in1
	// Insensitive connections
	always @(*) begin
		andOp_404_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_404_in1 = valid ? notOp_403_out : notOp_403_out;
	end
	// controller for andOp_406.andOp_406_in0
	// controller for andOp_406.andOp_406_in1
	// Insensitive connections
	always @(*) begin
		andOp_406_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_406_in1 = valid ? notOp_405_out : notOp_405_out;
	end
	// controller for andOp_407.andOp_407_in0
	// controller for andOp_407.andOp_407_in1
	// Insensitive connections
	always @(*) begin
		andOp_407_in0 = valid ? 1'd0 : 1'd0;
		andOp_407_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_409.andOp_409_in0
	// controller for andOp_409.andOp_409_in1
	// Insensitive connections
	always @(*) begin
		andOp_409_in0 = valid ? andOp_407_out : andOp_407_out;
		andOp_409_in1 = valid ? eq_408_out : eq_408_out;
	end
	// controller for andOp_411.andOp_411_in0
	// controller for andOp_411.andOp_411_in1
	// Insensitive connections
	always @(*) begin
		andOp_411_in0 = valid ? andOp_407_out : andOp_407_out;
		andOp_411_in1 = valid ? notOp_410_out : notOp_410_out;
	end
	// controller for andOp_413.andOp_413_in0
	// controller for andOp_413.andOp_413_in1
	// Insensitive connections
	always @(*) begin
		andOp_413_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_413_in1 = valid ? notOp_412_out : notOp_412_out;
	end
	// controller for andOp_415.andOp_415_in0
	// controller for andOp_415.andOp_415_in1
	// Insensitive connections
	always @(*) begin
		andOp_415_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_415_in1 = valid ? notOp_414_out : notOp_414_out;
	end
	// controller for andOp_416.andOp_416_in0
	// controller for andOp_416.andOp_416_in1
	// Insensitive connections
	always @(*) begin
		andOp_416_in0 = valid ? 1'd0 : 1'd0;
		andOp_416_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_418.andOp_418_in0
	// controller for andOp_418.andOp_418_in1
	// Insensitive connections
	always @(*) begin
		andOp_418_in0 = valid ? andOp_416_out : andOp_416_out;
		andOp_418_in1 = valid ? eq_417_out : eq_417_out;
	end
	// controller for andOp_420.andOp_420_in0
	// controller for andOp_420.andOp_420_in1
	// Insensitive connections
	always @(*) begin
		andOp_420_in0 = valid ? andOp_416_out : andOp_416_out;
		andOp_420_in1 = valid ? notOp_419_out : notOp_419_out;
	end
	// controller for andOp_422.andOp_422_in0
	// controller for andOp_422.andOp_422_in1
	// Insensitive connections
	always @(*) begin
		andOp_422_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_422_in1 = valid ? notOp_421_out : notOp_421_out;
	end
	// controller for andOp_424.andOp_424_in0
	// controller for andOp_424.andOp_424_in1
	// Insensitive connections
	always @(*) begin
		andOp_424_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_424_in1 = valid ? notOp_423_out : notOp_423_out;
	end
	// controller for andOp_426.andOp_426_in0
	// controller for andOp_426.andOp_426_in1
	// Insensitive connections
	always @(*) begin
		andOp_426_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_426_in1 = valid ? eq_425_out : eq_425_out;
	end
	// controller for andOp_428.andOp_428_in0
	// controller for andOp_428.andOp_428_in1
	// Insensitive connections
	always @(*) begin
		andOp_428_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_428_in1 = valid ? eq_427_out : eq_427_out;
	end
	// controller for andOp_430.andOp_430_in0
	// controller for andOp_430.andOp_430_in1
	// Insensitive connections
	always @(*) begin
		andOp_430_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_430_in1 = valid ? eq_429_out : eq_429_out;
	end
	// controller for andOp_432.andOp_432_in0
	// controller for andOp_432.andOp_432_in1
	// Insensitive connections
	always @(*) begin
		andOp_432_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_432_in1 = valid ? eq_431_out : eq_431_out;
	end
	// controller for andOp_434.andOp_434_in0
	// controller for andOp_434.andOp_434_in1
	// Insensitive connections
	always @(*) begin
		andOp_434_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_434_in1 = valid ? eq_433_out : eq_433_out;
	end
	// controller for andOp_435.andOp_435_in0
	// controller for andOp_435.andOp_435_in1
	// Insensitive connections
	always @(*) begin
		andOp_435_in0 = valid ? 1'd0 : 1'd0;
		andOp_435_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_437.andOp_437_in0
	// controller for andOp_437.andOp_437_in1
	// Insensitive connections
	always @(*) begin
		andOp_437_in0 = valid ? andOp_435_out : andOp_435_out;
		andOp_437_in1 = valid ? eq_436_out : eq_436_out;
	end
	// controller for andOp_439.andOp_439_in0
	// controller for andOp_439.andOp_439_in1
	// Insensitive connections
	always @(*) begin
		andOp_439_in0 = valid ? andOp_435_out : andOp_435_out;
		andOp_439_in1 = valid ? notOp_438_out : notOp_438_out;
	end
	// controller for andOp_441.andOp_441_in0
	// controller for andOp_441.andOp_441_in1
	// Insensitive connections
	always @(*) begin
		andOp_441_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_441_in1 = valid ? notOp_440_out : notOp_440_out;
	end
	// controller for andOp_443.andOp_443_in0
	// controller for andOp_443.andOp_443_in1
	// Insensitive connections
	always @(*) begin
		andOp_443_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_443_in1 = valid ? notOp_442_out : notOp_442_out;
	end
	// controller for andOp_444.andOp_444_in0
	// controller for andOp_444.andOp_444_in1
	// Insensitive connections
	always @(*) begin
		andOp_444_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_444_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_446.andOp_446_in0
	// controller for andOp_446.andOp_446_in1
	// Insensitive connections
	always @(*) begin
		andOp_446_in0 = valid ? andOp_444_out : andOp_444_out;
		andOp_446_in1 = valid ? eq_445_out : eq_445_out;
	end
	// controller for andOp_448.andOp_448_in0
	// controller for andOp_448.andOp_448_in1
	// Insensitive connections
	always @(*) begin
		andOp_448_in0 = valid ? andOp_444_out : andOp_444_out;
		andOp_448_in1 = valid ? notOp_447_out : notOp_447_out;
	end
	// controller for andOp_450.andOp_450_in0
	// controller for andOp_450.andOp_450_in1
	// Insensitive connections
	always @(*) begin
		andOp_450_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_450_in1 = valid ? notOp_449_out : notOp_449_out;
	end
	// controller for andOp_452.andOp_452_in0
	// controller for andOp_452.andOp_452_in1
	// Insensitive connections
	always @(*) begin
		andOp_452_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_452_in1 = valid ? notOp_451_out : notOp_451_out;
	end
	// controller for andOp_453.andOp_453_in0
	// controller for andOp_453.andOp_453_in1
	// Insensitive connections
	always @(*) begin
		andOp_453_in0 = valid ? 1'd0 : 1'd0;
		andOp_453_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_455.andOp_455_in0
	// controller for andOp_455.andOp_455_in1
	// Insensitive connections
	always @(*) begin
		andOp_455_in0 = valid ? andOp_453_out : andOp_453_out;
		andOp_455_in1 = valid ? eq_454_out : eq_454_out;
	end
	// controller for andOp_457.andOp_457_in0
	// controller for andOp_457.andOp_457_in1
	// Insensitive connections
	always @(*) begin
		andOp_457_in0 = valid ? andOp_453_out : andOp_453_out;
		andOp_457_in1 = valid ? notOp_456_out : notOp_456_out;
	end
	// controller for andOp_459.andOp_459_in0
	// controller for andOp_459.andOp_459_in1
	// Insensitive connections
	always @(*) begin
		andOp_459_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_459_in1 = valid ? notOp_458_out : notOp_458_out;
	end
	// controller for andOp_461.andOp_461_in0
	// controller for andOp_461.andOp_461_in1
	// Insensitive connections
	always @(*) begin
		andOp_461_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_461_in1 = valid ? notOp_460_out : notOp_460_out;
	end
	// controller for andOp_462.andOp_462_in0
	// controller for andOp_462.andOp_462_in1
	// Insensitive connections
	always @(*) begin
		andOp_462_in0 = valid ? 1'd0 : 1'd0;
		andOp_462_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_464.andOp_464_in0
	// controller for andOp_464.andOp_464_in1
	// Insensitive connections
	always @(*) begin
		andOp_464_in0 = valid ? andOp_462_out : andOp_462_out;
		andOp_464_in1 = valid ? eq_463_out : eq_463_out;
	end
	// controller for andOp_466.andOp_466_in0
	// controller for andOp_466.andOp_466_in1
	// Insensitive connections
	always @(*) begin
		andOp_466_in0 = valid ? andOp_462_out : andOp_462_out;
		andOp_466_in1 = valid ? notOp_465_out : notOp_465_out;
	end
	// controller for andOp_468.andOp_468_in0
	// controller for andOp_468.andOp_468_in1
	// Insensitive connections
	always @(*) begin
		andOp_468_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_468_in1 = valid ? notOp_467_out : notOp_467_out;
	end
	// controller for andOp_470.andOp_470_in0
	// controller for andOp_470.andOp_470_in1
	// Insensitive connections
	always @(*) begin
		andOp_470_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_470_in1 = valid ? notOp_469_out : notOp_469_out;
	end
	// controller for andOp_471.andOp_471_in0
	// controller for andOp_471.andOp_471_in1
	// Insensitive connections
	always @(*) begin
		andOp_471_in0 = valid ? 1'd0 : 1'd0;
		andOp_471_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_473.andOp_473_in0
	// controller for andOp_473.andOp_473_in1
	// Insensitive connections
	always @(*) begin
		andOp_473_in0 = valid ? andOp_471_out : andOp_471_out;
		andOp_473_in1 = valid ? eq_472_out : eq_472_out;
	end
	// controller for andOp_475.andOp_475_in0
	// controller for andOp_475.andOp_475_in1
	// Insensitive connections
	always @(*) begin
		andOp_475_in0 = valid ? andOp_471_out : andOp_471_out;
		andOp_475_in1 = valid ? notOp_474_out : notOp_474_out;
	end
	// controller for andOp_477.andOp_477_in0
	// controller for andOp_477.andOp_477_in1
	// Insensitive connections
	always @(*) begin
		andOp_477_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_477_in1 = valid ? notOp_476_out : notOp_476_out;
	end
	// controller for andOp_479.andOp_479_in0
	// controller for andOp_479.andOp_479_in1
	// Insensitive connections
	always @(*) begin
		andOp_479_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_479_in1 = valid ? notOp_478_out : notOp_478_out;
	end
	// controller for andOp_480.andOp_480_in0
	// controller for andOp_480.andOp_480_in1
	// Insensitive connections
	always @(*) begin
		andOp_480_in0 = valid ? 1'd0 : 1'd0;
		andOp_480_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_482.andOp_482_in0
	// controller for andOp_482.andOp_482_in1
	// Insensitive connections
	always @(*) begin
		andOp_482_in0 = valid ? andOp_480_out : andOp_480_out;
		andOp_482_in1 = valid ? eq_481_out : eq_481_out;
	end
	// controller for andOp_484.andOp_484_in0
	// controller for andOp_484.andOp_484_in1
	// Insensitive connections
	always @(*) begin
		andOp_484_in0 = valid ? andOp_480_out : andOp_480_out;
		andOp_484_in1 = valid ? notOp_483_out : notOp_483_out;
	end
	// controller for andOp_486.andOp_486_in0
	// controller for andOp_486.andOp_486_in1
	// Insensitive connections
	always @(*) begin
		andOp_486_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_486_in1 = valid ? notOp_485_out : notOp_485_out;
	end
	// controller for andOp_488.andOp_488_in0
	// controller for andOp_488.andOp_488_in1
	// Insensitive connections
	always @(*) begin
		andOp_488_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_488_in1 = valid ? notOp_487_out : notOp_487_out;
	end
	// controller for andOp_489.andOp_489_in0
	// controller for andOp_489.andOp_489_in1
	// Insensitive connections
	always @(*) begin
		andOp_489_in0 = valid ? 1'd0 : 1'd0;
		andOp_489_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_491.andOp_491_in0
	// controller for andOp_491.andOp_491_in1
	// Insensitive connections
	always @(*) begin
		andOp_491_in0 = valid ? andOp_489_out : andOp_489_out;
		andOp_491_in1 = valid ? eq_490_out : eq_490_out;
	end
	// controller for andOp_493.andOp_493_in0
	// controller for andOp_493.andOp_493_in1
	// Insensitive connections
	always @(*) begin
		andOp_493_in0 = valid ? andOp_489_out : andOp_489_out;
		andOp_493_in1 = valid ? notOp_492_out : notOp_492_out;
	end
	// controller for andOp_495.andOp_495_in0
	// controller for andOp_495.andOp_495_in1
	// Insensitive connections
	always @(*) begin
		andOp_495_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_495_in1 = valid ? notOp_494_out : notOp_494_out;
	end
	// controller for andOp_497.andOp_497_in0
	// controller for andOp_497.andOp_497_in1
	// Insensitive connections
	always @(*) begin
		andOp_497_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_497_in1 = valid ? notOp_496_out : notOp_496_out;
	end
	// controller for andOp_498.andOp_498_in0
	// controller for andOp_498.andOp_498_in1
	// Insensitive connections
	always @(*) begin
		andOp_498_in0 = valid ? 1'd0 : 1'd0;
		andOp_498_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_500.andOp_500_in0
	// controller for andOp_500.andOp_500_in1
	// Insensitive connections
	always @(*) begin
		andOp_500_in0 = valid ? andOp_498_out : andOp_498_out;
		andOp_500_in1 = valid ? eq_499_out : eq_499_out;
	end
	// controller for andOp_502.andOp_502_in0
	// controller for andOp_502.andOp_502_in1
	// Insensitive connections
	always @(*) begin
		andOp_502_in0 = valid ? andOp_498_out : andOp_498_out;
		andOp_502_in1 = valid ? notOp_501_out : notOp_501_out;
	end
	// controller for andOp_504.andOp_504_in0
	// controller for andOp_504.andOp_504_in1
	// Insensitive connections
	always @(*) begin
		andOp_504_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_504_in1 = valid ? notOp_503_out : notOp_503_out;
	end
	// controller for andOp_506.andOp_506_in0
	// controller for andOp_506.andOp_506_in1
	// Insensitive connections
	always @(*) begin
		andOp_506_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_506_in1 = valid ? notOp_505_out : notOp_505_out;
	end
	// controller for andOp_507.andOp_507_in0
	// controller for andOp_507.andOp_507_in1
	// Insensitive connections
	always @(*) begin
		andOp_507_in0 = valid ? 1'd0 : 1'd0;
		andOp_507_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_509.andOp_509_in0
	// controller for andOp_509.andOp_509_in1
	// Insensitive connections
	always @(*) begin
		andOp_509_in0 = valid ? andOp_507_out : andOp_507_out;
		andOp_509_in1 = valid ? eq_508_out : eq_508_out;
	end
	// controller for andOp_511.andOp_511_in0
	// controller for andOp_511.andOp_511_in1
	// Insensitive connections
	always @(*) begin
		andOp_511_in0 = valid ? andOp_507_out : andOp_507_out;
		andOp_511_in1 = valid ? notOp_510_out : notOp_510_out;
	end
	// controller for andOp_513.andOp_513_in0
	// controller for andOp_513.andOp_513_in1
	// Insensitive connections
	always @(*) begin
		andOp_513_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_513_in1 = valid ? notOp_512_out : notOp_512_out;
	end
	// controller for andOp_515.andOp_515_in0
	// controller for andOp_515.andOp_515_in1
	// Insensitive connections
	always @(*) begin
		andOp_515_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_515_in1 = valid ? notOp_514_out : notOp_514_out;
	end
	// controller for andOp_517.andOp_517_in0
	// controller for andOp_517.andOp_517_in1
	// Insensitive connections
	always @(*) begin
		andOp_517_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_517_in1 = valid ? eq_516_out : eq_516_out;
	end
	// controller for andOp_519.andOp_519_in0
	// controller for andOp_519.andOp_519_in1
	// Insensitive connections
	always @(*) begin
		andOp_519_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_519_in1 = valid ? eq_518_out : eq_518_out;
	end
	// controller for andOp_521.andOp_521_in0
	// controller for andOp_521.andOp_521_in1
	// Insensitive connections
	always @(*) begin
		andOp_521_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_521_in1 = valid ? eq_520_out : eq_520_out;
	end
	// controller for andOp_523.andOp_523_in0
	// controller for andOp_523.andOp_523_in1
	// Insensitive connections
	always @(*) begin
		andOp_523_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_523_in1 = valid ? eq_522_out : eq_522_out;
	end
	// controller for andOp_525.andOp_525_in0
	// controller for andOp_525.andOp_525_in1
	// Insensitive connections
	always @(*) begin
		andOp_525_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_525_in1 = valid ? eq_524_out : eq_524_out;
	end
	// controller for andOp_526.andOp_526_in0
	// controller for andOp_526.andOp_526_in1
	// Insensitive connections
	always @(*) begin
		andOp_526_in0 = valid ? 1'd0 : 1'd0;
		andOp_526_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_528.andOp_528_in0
	// controller for andOp_528.andOp_528_in1
	// Insensitive connections
	always @(*) begin
		andOp_528_in0 = valid ? andOp_526_out : andOp_526_out;
		andOp_528_in1 = valid ? eq_527_out : eq_527_out;
	end
	// controller for andOp_530.andOp_530_in0
	// controller for andOp_530.andOp_530_in1
	// Insensitive connections
	always @(*) begin
		andOp_530_in0 = valid ? andOp_526_out : andOp_526_out;
		andOp_530_in1 = valid ? notOp_529_out : notOp_529_out;
	end
	// controller for andOp_532.andOp_532_in0
	// controller for andOp_532.andOp_532_in1
	// Insensitive connections
	always @(*) begin
		andOp_532_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_532_in1 = valid ? notOp_531_out : notOp_531_out;
	end
	// controller for andOp_534.andOp_534_in0
	// controller for andOp_534.andOp_534_in1
	// Insensitive connections
	always @(*) begin
		andOp_534_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_534_in1 = valid ? notOp_533_out : notOp_533_out;
	end
	// controller for andOp_535.andOp_535_in0
	// controller for andOp_535.andOp_535_in1
	// Insensitive connections
	always @(*) begin
		andOp_535_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_535_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_537.andOp_537_in0
	// controller for andOp_537.andOp_537_in1
	// Insensitive connections
	always @(*) begin
		andOp_537_in0 = valid ? andOp_535_out : andOp_535_out;
		andOp_537_in1 = valid ? eq_536_out : eq_536_out;
	end
	// controller for andOp_539.andOp_539_in0
	// controller for andOp_539.andOp_539_in1
	// Insensitive connections
	always @(*) begin
		andOp_539_in0 = valid ? andOp_535_out : andOp_535_out;
		andOp_539_in1 = valid ? notOp_538_out : notOp_538_out;
	end
	// controller for andOp_541.andOp_541_in0
	// controller for andOp_541.andOp_541_in1
	// Insensitive connections
	always @(*) begin
		andOp_541_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_541_in1 = valid ? notOp_540_out : notOp_540_out;
	end
	// controller for andOp_543.andOp_543_in0
	// controller for andOp_543.andOp_543_in1
	// Insensitive connections
	always @(*) begin
		andOp_543_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_543_in1 = valid ? notOp_542_out : notOp_542_out;
	end
	// controller for andOp_544.andOp_544_in0
	// controller for andOp_544.andOp_544_in1
	// Insensitive connections
	always @(*) begin
		andOp_544_in0 = valid ? 1'd0 : 1'd0;
		andOp_544_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_546.andOp_546_in0
	// controller for andOp_546.andOp_546_in1
	// Insensitive connections
	always @(*) begin
		andOp_546_in0 = valid ? andOp_544_out : andOp_544_out;
		andOp_546_in1 = valid ? eq_545_out : eq_545_out;
	end
	// controller for andOp_548.andOp_548_in0
	// controller for andOp_548.andOp_548_in1
	// Insensitive connections
	always @(*) begin
		andOp_548_in0 = valid ? andOp_544_out : andOp_544_out;
		andOp_548_in1 = valid ? notOp_547_out : notOp_547_out;
	end
	// controller for andOp_550.andOp_550_in0
	// controller for andOp_550.andOp_550_in1
	// Insensitive connections
	always @(*) begin
		andOp_550_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_550_in1 = valid ? notOp_549_out : notOp_549_out;
	end
	// controller for andOp_552.andOp_552_in0
	// controller for andOp_552.andOp_552_in1
	// Insensitive connections
	always @(*) begin
		andOp_552_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_552_in1 = valid ? notOp_551_out : notOp_551_out;
	end
	// controller for andOp_553.andOp_553_in0
	// controller for andOp_553.andOp_553_in1
	// Insensitive connections
	always @(*) begin
		andOp_553_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_553_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_555.andOp_555_in0
	// controller for andOp_555.andOp_555_in1
	// Insensitive connections
	always @(*) begin
		andOp_555_in0 = valid ? andOp_553_out : andOp_553_out;
		andOp_555_in1 = valid ? eq_554_out : eq_554_out;
	end
	// controller for andOp_557.andOp_557_in0
	// controller for andOp_557.andOp_557_in1
	// Insensitive connections
	always @(*) begin
		andOp_557_in0 = valid ? andOp_553_out : andOp_553_out;
		andOp_557_in1 = valid ? notOp_556_out : notOp_556_out;
	end
	// controller for andOp_559.andOp_559_in0
	// controller for andOp_559.andOp_559_in1
	// Insensitive connections
	always @(*) begin
		andOp_559_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_559_in1 = valid ? notOp_558_out : notOp_558_out;
	end
	// controller for andOp_561.andOp_561_in0
	// controller for andOp_561.andOp_561_in1
	// Insensitive connections
	always @(*) begin
		andOp_561_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_561_in1 = valid ? notOp_560_out : notOp_560_out;
	end
	// controller for andOp_562.andOp_562_in0
	// controller for andOp_562.andOp_562_in1
	// Insensitive connections
	always @(*) begin
		andOp_562_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_562_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_564.andOp_564_in0
	// controller for andOp_564.andOp_564_in1
	// Insensitive connections
	always @(*) begin
		andOp_564_in0 = valid ? andOp_562_out : andOp_562_out;
		andOp_564_in1 = valid ? eq_563_out : eq_563_out;
	end
	// controller for andOp_566.andOp_566_in0
	// controller for andOp_566.andOp_566_in1
	// Insensitive connections
	always @(*) begin
		andOp_566_in0 = valid ? andOp_562_out : andOp_562_out;
		andOp_566_in1 = valid ? notOp_565_out : notOp_565_out;
	end
	// controller for andOp_568.andOp_568_in0
	// controller for andOp_568.andOp_568_in1
	// Insensitive connections
	always @(*) begin
		andOp_568_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_568_in1 = valid ? notOp_567_out : notOp_567_out;
	end
	// controller for andOp_570.andOp_570_in0
	// controller for andOp_570.andOp_570_in1
	// Insensitive connections
	always @(*) begin
		andOp_570_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_570_in1 = valid ? notOp_569_out : notOp_569_out;
	end
	// controller for andOp_571.andOp_571_in0
	// controller for andOp_571.andOp_571_in1
	// Insensitive connections
	always @(*) begin
		andOp_571_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_571_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_573.andOp_573_in0
	// controller for andOp_573.andOp_573_in1
	// Insensitive connections
	always @(*) begin
		andOp_573_in0 = valid ? andOp_571_out : andOp_571_out;
		andOp_573_in1 = valid ? eq_572_out : eq_572_out;
	end
	// controller for andOp_575.andOp_575_in0
	// controller for andOp_575.andOp_575_in1
	// Insensitive connections
	always @(*) begin
		andOp_575_in0 = valid ? andOp_571_out : andOp_571_out;
		andOp_575_in1 = valid ? notOp_574_out : notOp_574_out;
	end
	// controller for andOp_577.andOp_577_in0
	// controller for andOp_577.andOp_577_in1
	// Insensitive connections
	always @(*) begin
		andOp_577_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_577_in1 = valid ? notOp_576_out : notOp_576_out;
	end
	// controller for andOp_579.andOp_579_in0
	// controller for andOp_579.andOp_579_in1
	// Insensitive connections
	always @(*) begin
		andOp_579_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_579_in1 = valid ? notOp_578_out : notOp_578_out;
	end
	// controller for andOp_580.andOp_580_in0
	// controller for andOp_580.andOp_580_in1
	// Insensitive connections
	always @(*) begin
		andOp_580_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_580_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_582.andOp_582_in0
	// controller for andOp_582.andOp_582_in1
	// Insensitive connections
	always @(*) begin
		andOp_582_in0 = valid ? andOp_580_out : andOp_580_out;
		andOp_582_in1 = valid ? eq_581_out : eq_581_out;
	end
	// controller for andOp_584.andOp_584_in0
	// controller for andOp_584.andOp_584_in1
	// Insensitive connections
	always @(*) begin
		andOp_584_in0 = valid ? andOp_580_out : andOp_580_out;
		andOp_584_in1 = valid ? notOp_583_out : notOp_583_out;
	end
	// controller for andOp_586.andOp_586_in0
	// controller for andOp_586.andOp_586_in1
	// Insensitive connections
	always @(*) begin
		andOp_586_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_586_in1 = valid ? notOp_585_out : notOp_585_out;
	end
	// controller for andOp_588.andOp_588_in0
	// controller for andOp_588.andOp_588_in1
	// Insensitive connections
	always @(*) begin
		andOp_588_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_588_in1 = valid ? notOp_587_out : notOp_587_out;
	end
	// controller for andOp_589.andOp_589_in0
	// controller for andOp_589.andOp_589_in1
	// Insensitive connections
	always @(*) begin
		andOp_589_in0 = valid ? 1'd0 : 1'd0;
		andOp_589_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_591.andOp_591_in0
	// controller for andOp_591.andOp_591_in1
	// Insensitive connections
	always @(*) begin
		andOp_591_in0 = valid ? andOp_589_out : andOp_589_out;
		andOp_591_in1 = valid ? eq_590_out : eq_590_out;
	end
	// controller for andOp_593.andOp_593_in0
	// controller for andOp_593.andOp_593_in1
	// Insensitive connections
	always @(*) begin
		andOp_593_in0 = valid ? andOp_589_out : andOp_589_out;
		andOp_593_in1 = valid ? notOp_592_out : notOp_592_out;
	end
	// controller for andOp_595.andOp_595_in0
	// controller for andOp_595.andOp_595_in1
	// Insensitive connections
	always @(*) begin
		andOp_595_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_595_in1 = valid ? notOp_594_out : notOp_594_out;
	end
	// controller for andOp_597.andOp_597_in0
	// controller for andOp_597.andOp_597_in1
	// Insensitive connections
	always @(*) begin
		andOp_597_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_597_in1 = valid ? notOp_596_out : notOp_596_out;
	end
	// controller for andOp_598.andOp_598_in0
	// controller for andOp_598.andOp_598_in1
	// Insensitive connections
	always @(*) begin
		andOp_598_in0 = valid ? 1'd0 : 1'd0;
		andOp_598_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_600.andOp_600_in0
	// controller for andOp_600.andOp_600_in1
	// Insensitive connections
	always @(*) begin
		andOp_600_in0 = valid ? andOp_598_out : andOp_598_out;
		andOp_600_in1 = valid ? eq_599_out : eq_599_out;
	end
	// controller for andOp_602.andOp_602_in0
	// controller for andOp_602.andOp_602_in1
	// Insensitive connections
	always @(*) begin
		andOp_602_in0 = valid ? andOp_598_out : andOp_598_out;
		andOp_602_in1 = valid ? notOp_601_out : notOp_601_out;
	end
	// controller for andOp_604.andOp_604_in0
	// controller for andOp_604.andOp_604_in1
	// Insensitive connections
	always @(*) begin
		andOp_604_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_604_in1 = valid ? notOp_603_out : notOp_603_out;
	end
	// controller for andOp_606.andOp_606_in0
	// controller for andOp_606.andOp_606_in1
	// Insensitive connections
	always @(*) begin
		andOp_606_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_606_in1 = valid ? notOp_605_out : notOp_605_out;
	end
	// controller for andOp_608.andOp_608_in0
	// controller for andOp_608.andOp_608_in1
	// Insensitive connections
	always @(*) begin
		andOp_608_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_608_in1 = valid ? eq_607_out : eq_607_out;
	end
	// controller for andOp_610.andOp_610_in0
	// controller for andOp_610.andOp_610_in1
	// Insensitive connections
	always @(*) begin
		andOp_610_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_610_in1 = valid ? eq_609_out : eq_609_out;
	end
	// controller for andOp_612.andOp_612_in0
	// controller for andOp_612.andOp_612_in1
	// Insensitive connections
	always @(*) begin
		andOp_612_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_612_in1 = valid ? eq_611_out : eq_611_out;
	end
	// controller for andOp_614.andOp_614_in0
	// controller for andOp_614.andOp_614_in1
	// Insensitive connections
	always @(*) begin
		andOp_614_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_614_in1 = valid ? eq_613_out : eq_613_out;
	end
	// controller for andOp_616.andOp_616_in0
	// controller for andOp_616.andOp_616_in1
	// Insensitive connections
	always @(*) begin
		andOp_616_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_616_in1 = valid ? eq_615_out : eq_615_out;
	end
	// controller for andOp_617.andOp_617_in0
	// controller for andOp_617.andOp_617_in1
	// Insensitive connections
	always @(*) begin
		andOp_617_in0 = valid ? 1'd0 : 1'd0;
		andOp_617_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_619.andOp_619_in0
	// controller for andOp_619.andOp_619_in1
	// Insensitive connections
	always @(*) begin
		andOp_619_in0 = valid ? andOp_617_out : andOp_617_out;
		andOp_619_in1 = valid ? eq_618_out : eq_618_out;
	end
	// controller for andOp_621.andOp_621_in0
	// controller for andOp_621.andOp_621_in1
	// Insensitive connections
	always @(*) begin
		andOp_621_in0 = valid ? andOp_617_out : andOp_617_out;
		andOp_621_in1 = valid ? notOp_620_out : notOp_620_out;
	end
	// controller for andOp_623.andOp_623_in0
	// controller for andOp_623.andOp_623_in1
	// Insensitive connections
	always @(*) begin
		andOp_623_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_623_in1 = valid ? notOp_622_out : notOp_622_out;
	end
	// controller for andOp_625.andOp_625_in0
	// controller for andOp_625.andOp_625_in1
	// Insensitive connections
	always @(*) begin
		andOp_625_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_625_in1 = valid ? notOp_624_out : notOp_624_out;
	end
	// controller for andOp_626.andOp_626_in0
	// controller for andOp_626.andOp_626_in1
	// Insensitive connections
	always @(*) begin
		andOp_626_in0 = valid ? 1'd0 : 1'd0;
		andOp_626_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_628.andOp_628_in0
	// controller for andOp_628.andOp_628_in1
	// Insensitive connections
	always @(*) begin
		andOp_628_in0 = valid ? andOp_626_out : andOp_626_out;
		andOp_628_in1 = valid ? eq_627_out : eq_627_out;
	end
	// controller for andOp_630.andOp_630_in0
	// controller for andOp_630.andOp_630_in1
	// Insensitive connections
	always @(*) begin
		andOp_630_in0 = valid ? andOp_626_out : andOp_626_out;
		andOp_630_in1 = valid ? notOp_629_out : notOp_629_out;
	end
	// controller for andOp_632.andOp_632_in0
	// controller for andOp_632.andOp_632_in1
	// Insensitive connections
	always @(*) begin
		andOp_632_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_632_in1 = valid ? notOp_631_out : notOp_631_out;
	end
	// controller for andOp_634.andOp_634_in0
	// controller for andOp_634.andOp_634_in1
	// Insensitive connections
	always @(*) begin
		andOp_634_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_634_in1 = valid ? notOp_633_out : notOp_633_out;
	end
	// controller for andOp_635.andOp_635_in0
	// controller for andOp_635.andOp_635_in1
	// Insensitive connections
	always @(*) begin
		andOp_635_in0 = valid ? 1'd0 : 1'd0;
		andOp_635_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_637.andOp_637_in0
	// controller for andOp_637.andOp_637_in1
	// Insensitive connections
	always @(*) begin
		andOp_637_in0 = valid ? andOp_635_out : andOp_635_out;
		andOp_637_in1 = valid ? eq_636_out : eq_636_out;
	end
	// controller for andOp_639.andOp_639_in0
	// controller for andOp_639.andOp_639_in1
	// Insensitive connections
	always @(*) begin
		andOp_639_in0 = valid ? andOp_635_out : andOp_635_out;
		andOp_639_in1 = valid ? notOp_638_out : notOp_638_out;
	end
	// controller for andOp_641.andOp_641_in0
	// controller for andOp_641.andOp_641_in1
	// Insensitive connections
	always @(*) begin
		andOp_641_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_641_in1 = valid ? notOp_640_out : notOp_640_out;
	end
	// controller for andOp_643.andOp_643_in0
	// controller for andOp_643.andOp_643_in1
	// Insensitive connections
	always @(*) begin
		andOp_643_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_643_in1 = valid ? notOp_642_out : notOp_642_out;
	end
	// controller for andOp_644.andOp_644_in0
	// controller for andOp_644.andOp_644_in1
	// Insensitive connections
	always @(*) begin
		andOp_644_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_644_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_646.andOp_646_in0
	// controller for andOp_646.andOp_646_in1
	// Insensitive connections
	always @(*) begin
		andOp_646_in0 = valid ? andOp_644_out : andOp_644_out;
		andOp_646_in1 = valid ? eq_645_out : eq_645_out;
	end
	// controller for andOp_648.andOp_648_in0
	// controller for andOp_648.andOp_648_in1
	// Insensitive connections
	always @(*) begin
		andOp_648_in0 = valid ? andOp_644_out : andOp_644_out;
		andOp_648_in1 = valid ? notOp_647_out : notOp_647_out;
	end
	// controller for andOp_650.andOp_650_in0
	// controller for andOp_650.andOp_650_in1
	// Insensitive connections
	always @(*) begin
		andOp_650_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_650_in1 = valid ? notOp_649_out : notOp_649_out;
	end
	// controller for andOp_652.andOp_652_in0
	// controller for andOp_652.andOp_652_in1
	// Insensitive connections
	always @(*) begin
		andOp_652_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_652_in1 = valid ? notOp_651_out : notOp_651_out;
	end
	// controller for andOp_653.andOp_653_in0
	// controller for andOp_653.andOp_653_in1
	// Insensitive connections
	always @(*) begin
		andOp_653_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_653_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_655.andOp_655_in0
	// controller for andOp_655.andOp_655_in1
	// Insensitive connections
	always @(*) begin
		andOp_655_in0 = valid ? andOp_653_out : andOp_653_out;
		andOp_655_in1 = valid ? eq_654_out : eq_654_out;
	end
	// controller for andOp_657.andOp_657_in0
	// controller for andOp_657.andOp_657_in1
	// Insensitive connections
	always @(*) begin
		andOp_657_in0 = valid ? andOp_653_out : andOp_653_out;
		andOp_657_in1 = valid ? notOp_656_out : notOp_656_out;
	end
	// controller for andOp_659.andOp_659_in0
	// controller for andOp_659.andOp_659_in1
	// Insensitive connections
	always @(*) begin
		andOp_659_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_659_in1 = valid ? notOp_658_out : notOp_658_out;
	end
	// controller for andOp_661.andOp_661_in0
	// controller for andOp_661.andOp_661_in1
	// Insensitive connections
	always @(*) begin
		andOp_661_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_661_in1 = valid ? notOp_660_out : notOp_660_out;
	end
	// controller for andOp_662.andOp_662_in0
	// controller for andOp_662.andOp_662_in1
	// Insensitive connections
	always @(*) begin
		andOp_662_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_662_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_664.andOp_664_in0
	// controller for andOp_664.andOp_664_in1
	// Insensitive connections
	always @(*) begin
		andOp_664_in0 = valid ? andOp_662_out : andOp_662_out;
		andOp_664_in1 = valid ? eq_663_out : eq_663_out;
	end
	// controller for andOp_666.andOp_666_in0
	// controller for andOp_666.andOp_666_in1
	// Insensitive connections
	always @(*) begin
		andOp_666_in0 = valid ? andOp_662_out : andOp_662_out;
		andOp_666_in1 = valid ? notOp_665_out : notOp_665_out;
	end
	// controller for andOp_668.andOp_668_in0
	// controller for andOp_668.andOp_668_in1
	// Insensitive connections
	always @(*) begin
		andOp_668_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_668_in1 = valid ? notOp_667_out : notOp_667_out;
	end
	// controller for andOp_670.andOp_670_in0
	// controller for andOp_670.andOp_670_in1
	// Insensitive connections
	always @(*) begin
		andOp_670_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_670_in1 = valid ? notOp_669_out : notOp_669_out;
	end
	// controller for andOp_671.andOp_671_in0
	// controller for andOp_671.andOp_671_in1
	// Insensitive connections
	always @(*) begin
		andOp_671_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_671_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_673.andOp_673_in0
	// controller for andOp_673.andOp_673_in1
	// Insensitive connections
	always @(*) begin
		andOp_673_in0 = valid ? andOp_671_out : andOp_671_out;
		andOp_673_in1 = valid ? eq_672_out : eq_672_out;
	end
	// controller for andOp_675.andOp_675_in0
	// controller for andOp_675.andOp_675_in1
	// Insensitive connections
	always @(*) begin
		andOp_675_in0 = valid ? andOp_671_out : andOp_671_out;
		andOp_675_in1 = valid ? notOp_674_out : notOp_674_out;
	end
	// controller for andOp_677.andOp_677_in0
	// controller for andOp_677.andOp_677_in1
	// Insensitive connections
	always @(*) begin
		andOp_677_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_677_in1 = valid ? notOp_676_out : notOp_676_out;
	end
	// controller for andOp_679.andOp_679_in0
	// controller for andOp_679.andOp_679_in1
	// Insensitive connections
	always @(*) begin
		andOp_679_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_679_in1 = valid ? notOp_678_out : notOp_678_out;
	end
	// controller for andOp_680.andOp_680_in0
	// controller for andOp_680.andOp_680_in1
	// Insensitive connections
	always @(*) begin
		andOp_680_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_680_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_682.andOp_682_in0
	// controller for andOp_682.andOp_682_in1
	// Insensitive connections
	always @(*) begin
		andOp_682_in0 = valid ? andOp_680_out : andOp_680_out;
		andOp_682_in1 = valid ? eq_681_out : eq_681_out;
	end
	// controller for andOp_684.andOp_684_in0
	// controller for andOp_684.andOp_684_in1
	// Insensitive connections
	always @(*) begin
		andOp_684_in0 = valid ? andOp_680_out : andOp_680_out;
		andOp_684_in1 = valid ? notOp_683_out : notOp_683_out;
	end
	// controller for andOp_686.andOp_686_in0
	// controller for andOp_686.andOp_686_in1
	// Insensitive connections
	always @(*) begin
		andOp_686_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_686_in1 = valid ? notOp_685_out : notOp_685_out;
	end
	// controller for andOp_688.andOp_688_in0
	// controller for andOp_688.andOp_688_in1
	// Insensitive connections
	always @(*) begin
		andOp_688_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_688_in1 = valid ? notOp_687_out : notOp_687_out;
	end
	// controller for andOp_689.andOp_689_in0
	// controller for andOp_689.andOp_689_in1
	// Insensitive connections
	always @(*) begin
		andOp_689_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
		andOp_689_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_691.andOp_691_in0
	// controller for andOp_691.andOp_691_in1
	// Insensitive connections
	always @(*) begin
		andOp_691_in0 = valid ? andOp_689_out : andOp_689_out;
		andOp_691_in1 = valid ? eq_690_out : eq_690_out;
	end
	// controller for andOp_693.andOp_693_in0
	// controller for andOp_693.andOp_693_in1
	// Insensitive connections
	always @(*) begin
		andOp_693_in0 = valid ? andOp_689_out : andOp_689_out;
		andOp_693_in1 = valid ? notOp_692_out : notOp_692_out;
	end
	// controller for andOp_695.andOp_695_in0
	// controller for andOp_695.andOp_695_in1
	// Insensitive connections
	always @(*) begin
		andOp_695_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_695_in1 = valid ? notOp_694_out : notOp_694_out;
	end
	// controller for andOp_697.andOp_697_in0
	// controller for andOp_697.andOp_697_in1
	// Insensitive connections
	always @(*) begin
		andOp_697_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_697_in1 = valid ? notOp_696_out : notOp_696_out;
	end
	// controller for andOp_90.andOp_90_in0
	// controller for andOp_90.andOp_90_in1
	// Insensitive connections
	always @(*) begin
		andOp_90_in0 = valid ? bb_0_active_in_state_1_out_data : bb_0_active_in_state_1_out_data;
		andOp_90_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_91.andOp_91_in0
	// controller for andOp_91.andOp_91_in1
	// Insensitive connections
	always @(*) begin
		andOp_91_in0 = valid ? andOp_90_out : andOp_90_out;
		andOp_91_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_93.andOp_93_in0
	// controller for andOp_93.andOp_93_in1
	// Insensitive connections
	always @(*) begin
		andOp_93_in0 = valid ? bb_8_active_in_state_1_out_data : bb_8_active_in_state_1_out_data;
		andOp_93_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_94.andOp_94_in0
	// controller for andOp_94.andOp_94_in1
	// Insensitive connections
	always @(*) begin
		andOp_94_in0 = valid ? andOp_93_out : andOp_93_out;
		andOp_94_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_96.andOp_96_in0
	// controller for andOp_96.andOp_96_in1
	// Insensitive connections
	always @(*) begin
		andOp_96_in0 = valid ? bb_0_active_in_state_1_out_data : bb_0_active_in_state_1_out_data;
		andOp_96_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_97.andOp_97_in0
	// controller for andOp_97.andOp_97_in1
	// Insensitive connections
	always @(*) begin
		andOp_97_in0 = valid ? andOp_96_out : andOp_96_out;
		andOp_97_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_99.andOp_99_in0
	// controller for andOp_99.andOp_99_in1
	// Insensitive connections
	always @(*) begin
		andOp_99_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_99_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_141_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_active_in_state_1.bb_0_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_1_in_data = eq_144_out;
		end else begin
			bb_0_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_164_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_1.bb_0_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_168_out) begin 
			bb_0_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_2.bb_10_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_2_in_data = eq_149_out;
		end else begin
			bb_10_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_3.bb_10_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_3_in_data = eq_152_out;
		end else begin
			bb_10_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_2.bb_10_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_175_out) begin 
			bb_10_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_3.bb_10_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_179_out) begin 
			bb_10_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_4.bb_1_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_4_in_data = orOp_163_out;
		end else begin
			bb_1_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_4.bb_1_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_195_out) begin 
			bb_1_predecessor_in_state_4_in_data = 32'd4;
		end else if (eq_193_out) begin 
			bb_1_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_4.bb_2_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_4_in_data = orOp_161_out;
		end else begin
			bb_2_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_4.bb_2_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_192_out) begin 
			bb_2_predecessor_in_state_4_in_data = 32'd7;
		end else if (eq_190_out) begin 
			bb_2_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_1.bb_3_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_1_in_data = orOp_146_out;
		end else begin
			bb_3_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_1.bb_3_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_171_out) begin 
			bb_3_predecessor_in_state_1_in_data = 32'd0;
		end else if (eq_169_out) begin 
			bb_3_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_3.bb_4_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_3_in_data = orOp_151_out;
		end else begin
			bb_4_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_4.bb_4_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_4_in_data = eq_159_out;
		end else begin
			bb_4_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_3.bb_4_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_178_out) begin 
			bb_4_predecessor_in_state_3_in_data = 32'd10;
		end else if (eq_176_out) begin 
			bb_4_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_4.bb_4_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_189_out) begin 
			bb_4_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_5_active_in_state_4.bb_5_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_5_active_in_state_4_in_data = orOp_154_out;
		end else begin
			bb_5_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_5_predecessor_in_state_4.bb_5_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_182_out) begin 
			bb_5_predecessor_in_state_4_in_data = 32'd1;
		end else if (eq_180_out) begin 
			bb_5_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_5_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_6_active_in_state_4.bb_6_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_6_active_in_state_4_in_data = orOp_156_out;
		end else begin
			bb_6_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_6_predecessor_in_state_4.bb_6_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_185_out) begin 
			bb_6_predecessor_in_state_4_in_data = 32'd5;
		end else if (eq_183_out) begin 
			bb_6_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_6_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_7_active_in_state_4.bb_7_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_7_active_in_state_4_in_data = orOp_158_out;
		end else begin
			bb_7_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_7_predecessor_in_state_4.bb_7_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_188_out) begin 
			bb_7_predecessor_in_state_4_in_data = 32'd6;
		end else if (eq_186_out) begin 
			bb_7_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_7_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_8_active_in_state_1.bb_8_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_state_1_in_data = orOp_143_out;
		end else begin
			bb_8_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_8_predecessor_in_state_1.bb_8_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_167_out) begin 
			bb_8_predecessor_in_state_1_in_data = 32'd3;
		end else if (eq_165_out) begin 
			bb_8_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_8_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_9_active_in_state_1.bb_9_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_9_active_in_state_1_in_data = orOp_148_out;
		end else begin
			bb_9_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_9_predecessor_in_state_1.bb_9_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_174_out) begin 
			bb_9_predecessor_in_state_1_in_data = 32'd8;
		end else if (eq_172_out) begin 
			bb_9_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_9_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_91_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_92_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_1.br_0_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_97_out) begin 
			br_0_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_98_out) begin 
			br_0_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_2.br_10_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_109_out) begin 
			br_10_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_110_out) begin 
			br_10_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_3.br_10_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_118_out) begin 
			br_10_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_119_out) begin 
			br_10_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_1_happened_in_state_4.br_1_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_139_out) begin 
			br_1_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_140_out) begin 
			br_1_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_1_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_1.br_3_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_100_out) begin 
			br_3_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_101_out) begin 
			br_3_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_3.br_4_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_112_out) begin 
			br_4_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_113_out) begin 
			br_4_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_4.br_4_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_133_out) begin 
			br_4_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_134_out) begin 
			br_4_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_5_happened_in_state_4.br_5_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_121_out) begin 
			br_5_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_122_out) begin 
			br_5_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_5_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_6_happened_in_state_4.br_6_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_124_out) begin 
			br_6_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_125_out) begin 
			br_6_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_6_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_7_happened_in_state_4.br_7_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_130_out) begin 
			br_7_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_131_out) begin 
			br_7_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_7_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_8_happened_in_state_1.br_8_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_94_out) begin 
			br_8_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_95_out) begin 
			br_8_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_8_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_9_happened_in_state_1.br_9_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_103_out) begin 
			br_9_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_104_out) begin 
			br_9_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_9_happened_in_state_1_in_data = 0;
		end
	end
	// controller for concat_207.concat_207_in0
	// controller for concat_207.concat_207_in1
	// Insensitive connections
	always @(*) begin
		concat_207_in0 = valid ? data_in_1_29_out_data : data_in_1_29_out_data;
		concat_207_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for concat_208.concat_208_in0
	// controller for concat_208.concat_208_in1
	// Insensitive connections
	always @(*) begin
		concat_208_in0 = valid ? 32'd4 : 32'd4;
		concat_208_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for data_in_0_1.data_in_0_1_in_data
	always @(*) begin
		if (andOp_244_out) begin 
			data_in_0_1_in_data = data_store_0_0;
		end else if (andOp_246_out) begin 
			data_in_0_1_in_data = data_store_1_18;
		end else if (andOp_248_out) begin 
			data_in_0_1_in_data = data_store_2_36;
		end else if (andOp_250_out) begin 
			data_in_0_1_in_data = data_store_3_54;
		end else if (andOp_252_out) begin 
			data_in_0_1_in_data = data_store_4_72;
		end else begin
			data_in_0_1_in_data = 0;
		end
	end
	// controller for data_in_0_11.data_in_0_11_in_data
	always @(*) begin
		if (andOp_244_out) begin 
			data_in_0_11_in_data = data_store_0_10;
		end else if (andOp_246_out) begin 
			data_in_0_11_in_data = data_store_1_28;
		end else if (andOp_248_out) begin 
			data_in_0_11_in_data = data_store_2_46;
		end else if (andOp_250_out) begin 
			data_in_0_11_in_data = data_store_3_64;
		end else if (andOp_252_out) begin 
			data_in_0_11_in_data = data_store_4_82;
		end else begin
			data_in_0_11_in_data = 0;
		end
	end
	// controller for data_in_0_13.data_in_0_13_in_data
	always @(*) begin
		if (andOp_244_out) begin 
			data_in_0_13_in_data = data_store_0_12;
		end else if (andOp_246_out) begin 
			data_in_0_13_in_data = data_store_1_30;
		end else if (andOp_248_out) begin 
			data_in_0_13_in_data = data_store_2_48;
		end else if (andOp_250_out) begin 
			data_in_0_13_in_data = data_store_3_66;
		end else if (andOp_252_out) begin 
			data_in_0_13_in_data = data_store_4_84;
		end else begin
			data_in_0_13_in_data = 0;
		end
	end
	// controller for data_in_0_15.data_in_0_15_in_data
	always @(*) begin
		if (andOp_244_out) begin 
			data_in_0_15_in_data = data_store_0_14;
		end else if (andOp_246_out) begin 
			data_in_0_15_in_data = data_store_1_32;
		end else if (andOp_248_out) begin 
			data_in_0_15_in_data = data_store_2_50;
		end else if (andOp_250_out) begin 
			data_in_0_15_in_data = data_store_3_68;
		end else if (andOp_252_out) begin 
			data_in_0_15_in_data = data_store_4_86;
		end else begin
			data_in_0_15_in_data = 0;
		end
	end
	// controller for data_in_0_17.data_in_0_17_in_data
	always @(*) begin
		if (andOp_244_out) begin 
			data_in_0_17_in_data = data_store_0_16;
		end else if (andOp_246_out) begin 
			data_in_0_17_in_data = data_store_1_34;
		end else if (andOp_248_out) begin 
			data_in_0_17_in_data = data_store_2_52;
		end else if (andOp_250_out) begin 
			data_in_0_17_in_data = data_store_3_70;
		end else if (andOp_252_out) begin 
			data_in_0_17_in_data = data_store_4_88;
		end else begin
			data_in_0_17_in_data = 0;
		end
	end
	// controller for data_in_0_3.data_in_0_3_in_data
	always @(*) begin
		if (andOp_244_out) begin 
			data_in_0_3_in_data = data_store_0_2;
		end else if (andOp_246_out) begin 
			data_in_0_3_in_data = data_store_1_20;
		end else if (andOp_248_out) begin 
			data_in_0_3_in_data = data_store_2_38;
		end else if (andOp_250_out) begin 
			data_in_0_3_in_data = data_store_3_56;
		end else if (andOp_252_out) begin 
			data_in_0_3_in_data = data_store_4_74;
		end else begin
			data_in_0_3_in_data = 0;
		end
	end
	// controller for data_in_0_5.data_in_0_5_in_data
	always @(*) begin
		if (andOp_244_out) begin 
			data_in_0_5_in_data = data_store_0_4;
		end else if (andOp_246_out) begin 
			data_in_0_5_in_data = data_store_1_22;
		end else if (andOp_248_out) begin 
			data_in_0_5_in_data = data_store_2_40;
		end else if (andOp_250_out) begin 
			data_in_0_5_in_data = data_store_3_58;
		end else if (andOp_252_out) begin 
			data_in_0_5_in_data = data_store_4_76;
		end else begin
			data_in_0_5_in_data = 0;
		end
	end
	// controller for data_in_0_7.data_in_0_7_in_data
	always @(*) begin
		if (andOp_244_out) begin 
			data_in_0_7_in_data = data_store_0_6;
		end else if (andOp_246_out) begin 
			data_in_0_7_in_data = data_store_1_24;
		end else if (andOp_248_out) begin 
			data_in_0_7_in_data = data_store_2_42;
		end else if (andOp_250_out) begin 
			data_in_0_7_in_data = data_store_3_60;
		end else if (andOp_252_out) begin 
			data_in_0_7_in_data = data_store_4_78;
		end else begin
			data_in_0_7_in_data = 0;
		end
	end
	// controller for data_in_0_9.data_in_0_9_in_data
	always @(*) begin
		if (andOp_244_out) begin 
			data_in_0_9_in_data = data_store_0_8;
		end else if (andOp_246_out) begin 
			data_in_0_9_in_data = data_store_1_26;
		end else if (andOp_248_out) begin 
			data_in_0_9_in_data = data_store_2_44;
		end else if (andOp_250_out) begin 
			data_in_0_9_in_data = data_store_3_62;
		end else if (andOp_252_out) begin 
			data_in_0_9_in_data = data_store_4_80;
		end else begin
			data_in_0_9_in_data = 0;
		end
	end
	// controller for data_in_1_19.data_in_1_19_in_data
	always @(*) begin
		if (andOp_335_out) begin 
			data_in_1_19_in_data = data_store_0_0;
		end else if (andOp_337_out) begin 
			data_in_1_19_in_data = data_store_1_18;
		end else if (andOp_339_out) begin 
			data_in_1_19_in_data = data_store_2_36;
		end else if (andOp_341_out) begin 
			data_in_1_19_in_data = data_store_3_54;
		end else if (andOp_343_out) begin 
			data_in_1_19_in_data = data_store_4_72;
		end else begin
			data_in_1_19_in_data = 0;
		end
	end
	// controller for data_in_1_21.data_in_1_21_in_data
	always @(*) begin
		if (andOp_335_out) begin 
			data_in_1_21_in_data = data_store_0_2;
		end else if (andOp_337_out) begin 
			data_in_1_21_in_data = data_store_1_20;
		end else if (andOp_339_out) begin 
			data_in_1_21_in_data = data_store_2_38;
		end else if (andOp_341_out) begin 
			data_in_1_21_in_data = data_store_3_56;
		end else if (andOp_343_out) begin 
			data_in_1_21_in_data = data_store_4_74;
		end else begin
			data_in_1_21_in_data = 0;
		end
	end
	// controller for data_in_1_23.data_in_1_23_in_data
	always @(*) begin
		if (andOp_335_out) begin 
			data_in_1_23_in_data = data_store_0_4;
		end else if (andOp_337_out) begin 
			data_in_1_23_in_data = data_store_1_22;
		end else if (andOp_339_out) begin 
			data_in_1_23_in_data = data_store_2_40;
		end else if (andOp_341_out) begin 
			data_in_1_23_in_data = data_store_3_58;
		end else if (andOp_343_out) begin 
			data_in_1_23_in_data = data_store_4_76;
		end else begin
			data_in_1_23_in_data = 0;
		end
	end
	// controller for data_in_1_25.data_in_1_25_in_data
	always @(*) begin
		if (andOp_335_out) begin 
			data_in_1_25_in_data = data_store_0_6;
		end else if (andOp_337_out) begin 
			data_in_1_25_in_data = data_store_1_24;
		end else if (andOp_339_out) begin 
			data_in_1_25_in_data = data_store_2_42;
		end else if (andOp_341_out) begin 
			data_in_1_25_in_data = data_store_3_60;
		end else if (andOp_343_out) begin 
			data_in_1_25_in_data = data_store_4_78;
		end else begin
			data_in_1_25_in_data = 0;
		end
	end
	// controller for data_in_1_27.data_in_1_27_in_data
	always @(*) begin
		if (andOp_335_out) begin 
			data_in_1_27_in_data = data_store_0_8;
		end else if (andOp_337_out) begin 
			data_in_1_27_in_data = data_store_1_26;
		end else if (andOp_339_out) begin 
			data_in_1_27_in_data = data_store_2_44;
		end else if (andOp_341_out) begin 
			data_in_1_27_in_data = data_store_3_62;
		end else if (andOp_343_out) begin 
			data_in_1_27_in_data = data_store_4_80;
		end else begin
			data_in_1_27_in_data = 0;
		end
	end
	// controller for data_in_1_29.data_in_1_29_in_data
	always @(*) begin
		if (andOp_335_out) begin 
			data_in_1_29_in_data = data_store_0_10;
		end else if (andOp_337_out) begin 
			data_in_1_29_in_data = data_store_1_28;
		end else if (andOp_339_out) begin 
			data_in_1_29_in_data = data_store_2_46;
		end else if (andOp_341_out) begin 
			data_in_1_29_in_data = data_store_3_64;
		end else if (andOp_343_out) begin 
			data_in_1_29_in_data = data_store_4_82;
		end else begin
			data_in_1_29_in_data = 0;
		end
	end
	// controller for data_in_1_31.data_in_1_31_in_data
	always @(*) begin
		if (andOp_335_out) begin 
			data_in_1_31_in_data = data_store_0_12;
		end else if (andOp_337_out) begin 
			data_in_1_31_in_data = data_store_1_30;
		end else if (andOp_339_out) begin 
			data_in_1_31_in_data = data_store_2_48;
		end else if (andOp_341_out) begin 
			data_in_1_31_in_data = data_store_3_66;
		end else if (andOp_343_out) begin 
			data_in_1_31_in_data = data_store_4_84;
		end else begin
			data_in_1_31_in_data = 0;
		end
	end
	// controller for data_in_1_33.data_in_1_33_in_data
	always @(*) begin
		if (andOp_335_out) begin 
			data_in_1_33_in_data = data_store_0_14;
		end else if (andOp_337_out) begin 
			data_in_1_33_in_data = data_store_1_32;
		end else if (andOp_339_out) begin 
			data_in_1_33_in_data = data_store_2_50;
		end else if (andOp_341_out) begin 
			data_in_1_33_in_data = data_store_3_68;
		end else if (andOp_343_out) begin 
			data_in_1_33_in_data = data_store_4_86;
		end else begin
			data_in_1_33_in_data = 0;
		end
	end
	// controller for data_in_1_35.data_in_1_35_in_data
	always @(*) begin
		if (andOp_335_out) begin 
			data_in_1_35_in_data = data_store_0_16;
		end else if (andOp_337_out) begin 
			data_in_1_35_in_data = data_store_1_34;
		end else if (andOp_339_out) begin 
			data_in_1_35_in_data = data_store_2_52;
		end else if (andOp_341_out) begin 
			data_in_1_35_in_data = data_store_3_70;
		end else if (andOp_343_out) begin 
			data_in_1_35_in_data = data_store_4_88;
		end else begin
			data_in_1_35_in_data = 0;
		end
	end
	// controller for data_in_2_37.data_in_2_37_in_data
	always @(*) begin
		if (andOp_426_out) begin 
			data_in_2_37_in_data = data_store_0_0;
		end else if (andOp_428_out) begin 
			data_in_2_37_in_data = data_store_1_18;
		end else if (andOp_430_out) begin 
			data_in_2_37_in_data = data_store_2_36;
		end else if (andOp_432_out) begin 
			data_in_2_37_in_data = data_store_3_54;
		end else if (andOp_434_out) begin 
			data_in_2_37_in_data = data_store_4_72;
		end else begin
			data_in_2_37_in_data = 0;
		end
	end
	// controller for data_in_2_39.data_in_2_39_in_data
	always @(*) begin
		if (andOp_426_out) begin 
			data_in_2_39_in_data = data_store_0_2;
		end else if (andOp_428_out) begin 
			data_in_2_39_in_data = data_store_1_20;
		end else if (andOp_430_out) begin 
			data_in_2_39_in_data = data_store_2_38;
		end else if (andOp_432_out) begin 
			data_in_2_39_in_data = data_store_3_56;
		end else if (andOp_434_out) begin 
			data_in_2_39_in_data = data_store_4_74;
		end else begin
			data_in_2_39_in_data = 0;
		end
	end
	// controller for data_in_2_41.data_in_2_41_in_data
	always @(*) begin
		if (andOp_426_out) begin 
			data_in_2_41_in_data = data_store_0_4;
		end else if (andOp_428_out) begin 
			data_in_2_41_in_data = data_store_1_22;
		end else if (andOp_430_out) begin 
			data_in_2_41_in_data = data_store_2_40;
		end else if (andOp_432_out) begin 
			data_in_2_41_in_data = data_store_3_58;
		end else if (andOp_434_out) begin 
			data_in_2_41_in_data = data_store_4_76;
		end else begin
			data_in_2_41_in_data = 0;
		end
	end
	// controller for data_in_2_43.data_in_2_43_in_data
	always @(*) begin
		if (andOp_426_out) begin 
			data_in_2_43_in_data = data_store_0_6;
		end else if (andOp_428_out) begin 
			data_in_2_43_in_data = data_store_1_24;
		end else if (andOp_430_out) begin 
			data_in_2_43_in_data = data_store_2_42;
		end else if (andOp_432_out) begin 
			data_in_2_43_in_data = data_store_3_60;
		end else if (andOp_434_out) begin 
			data_in_2_43_in_data = data_store_4_78;
		end else begin
			data_in_2_43_in_data = 0;
		end
	end
	// controller for data_in_2_45.data_in_2_45_in_data
	always @(*) begin
		if (andOp_426_out) begin 
			data_in_2_45_in_data = data_store_0_8;
		end else if (andOp_428_out) begin 
			data_in_2_45_in_data = data_store_1_26;
		end else if (andOp_430_out) begin 
			data_in_2_45_in_data = data_store_2_44;
		end else if (andOp_432_out) begin 
			data_in_2_45_in_data = data_store_3_62;
		end else if (andOp_434_out) begin 
			data_in_2_45_in_data = data_store_4_80;
		end else begin
			data_in_2_45_in_data = 0;
		end
	end
	// controller for data_in_2_47.data_in_2_47_in_data
	always @(*) begin
		if (andOp_426_out) begin 
			data_in_2_47_in_data = data_store_0_10;
		end else if (andOp_428_out) begin 
			data_in_2_47_in_data = data_store_1_28;
		end else if (andOp_430_out) begin 
			data_in_2_47_in_data = data_store_2_46;
		end else if (andOp_432_out) begin 
			data_in_2_47_in_data = data_store_3_64;
		end else if (andOp_434_out) begin 
			data_in_2_47_in_data = data_store_4_82;
		end else begin
			data_in_2_47_in_data = 0;
		end
	end
	// controller for data_in_2_49.data_in_2_49_in_data
	always @(*) begin
		if (andOp_426_out) begin 
			data_in_2_49_in_data = data_store_0_12;
		end else if (andOp_428_out) begin 
			data_in_2_49_in_data = data_store_1_30;
		end else if (andOp_430_out) begin 
			data_in_2_49_in_data = data_store_2_48;
		end else if (andOp_432_out) begin 
			data_in_2_49_in_data = data_store_3_66;
		end else if (andOp_434_out) begin 
			data_in_2_49_in_data = data_store_4_84;
		end else begin
			data_in_2_49_in_data = 0;
		end
	end
	// controller for data_in_2_51.data_in_2_51_in_data
	always @(*) begin
		if (andOp_426_out) begin 
			data_in_2_51_in_data = data_store_0_14;
		end else if (andOp_428_out) begin 
			data_in_2_51_in_data = data_store_1_32;
		end else if (andOp_430_out) begin 
			data_in_2_51_in_data = data_store_2_50;
		end else if (andOp_432_out) begin 
			data_in_2_51_in_data = data_store_3_68;
		end else if (andOp_434_out) begin 
			data_in_2_51_in_data = data_store_4_86;
		end else begin
			data_in_2_51_in_data = 0;
		end
	end
	// controller for data_in_2_53.data_in_2_53_in_data
	always @(*) begin
		if (andOp_426_out) begin 
			data_in_2_53_in_data = data_store_0_16;
		end else if (andOp_428_out) begin 
			data_in_2_53_in_data = data_store_1_34;
		end else if (andOp_430_out) begin 
			data_in_2_53_in_data = data_store_2_52;
		end else if (andOp_432_out) begin 
			data_in_2_53_in_data = data_store_3_70;
		end else if (andOp_434_out) begin 
			data_in_2_53_in_data = data_store_4_88;
		end else begin
			data_in_2_53_in_data = 0;
		end
	end
	// controller for data_in_3_55.data_in_3_55_in_data
	always @(*) begin
		if (andOp_517_out) begin 
			data_in_3_55_in_data = data_store_0_0;
		end else if (andOp_519_out) begin 
			data_in_3_55_in_data = data_store_1_18;
		end else if (andOp_521_out) begin 
			data_in_3_55_in_data = data_store_2_36;
		end else if (andOp_523_out) begin 
			data_in_3_55_in_data = data_store_3_54;
		end else if (andOp_525_out) begin 
			data_in_3_55_in_data = data_store_4_72;
		end else begin
			data_in_3_55_in_data = 0;
		end
	end
	// controller for data_in_3_57.data_in_3_57_in_data
	always @(*) begin
		if (andOp_517_out) begin 
			data_in_3_57_in_data = data_store_0_2;
		end else if (andOp_519_out) begin 
			data_in_3_57_in_data = data_store_1_20;
		end else if (andOp_521_out) begin 
			data_in_3_57_in_data = data_store_2_38;
		end else if (andOp_523_out) begin 
			data_in_3_57_in_data = data_store_3_56;
		end else if (andOp_525_out) begin 
			data_in_3_57_in_data = data_store_4_74;
		end else begin
			data_in_3_57_in_data = 0;
		end
	end
	// controller for data_in_3_59.data_in_3_59_in_data
	always @(*) begin
		if (andOp_517_out) begin 
			data_in_3_59_in_data = data_store_0_4;
		end else if (andOp_519_out) begin 
			data_in_3_59_in_data = data_store_1_22;
		end else if (andOp_521_out) begin 
			data_in_3_59_in_data = data_store_2_40;
		end else if (andOp_523_out) begin 
			data_in_3_59_in_data = data_store_3_58;
		end else if (andOp_525_out) begin 
			data_in_3_59_in_data = data_store_4_76;
		end else begin
			data_in_3_59_in_data = 0;
		end
	end
	// controller for data_in_3_61.data_in_3_61_in_data
	always @(*) begin
		if (andOp_517_out) begin 
			data_in_3_61_in_data = data_store_0_6;
		end else if (andOp_519_out) begin 
			data_in_3_61_in_data = data_store_1_24;
		end else if (andOp_521_out) begin 
			data_in_3_61_in_data = data_store_2_42;
		end else if (andOp_523_out) begin 
			data_in_3_61_in_data = data_store_3_60;
		end else if (andOp_525_out) begin 
			data_in_3_61_in_data = data_store_4_78;
		end else begin
			data_in_3_61_in_data = 0;
		end
	end
	// controller for data_in_3_63.data_in_3_63_in_data
	always @(*) begin
		if (andOp_517_out) begin 
			data_in_3_63_in_data = data_store_0_8;
		end else if (andOp_519_out) begin 
			data_in_3_63_in_data = data_store_1_26;
		end else if (andOp_521_out) begin 
			data_in_3_63_in_data = data_store_2_44;
		end else if (andOp_523_out) begin 
			data_in_3_63_in_data = data_store_3_62;
		end else if (andOp_525_out) begin 
			data_in_3_63_in_data = data_store_4_80;
		end else begin
			data_in_3_63_in_data = 0;
		end
	end
	// controller for data_in_3_65.data_in_3_65_in_data
	always @(*) begin
		if (andOp_517_out) begin 
			data_in_3_65_in_data = data_store_0_10;
		end else if (andOp_519_out) begin 
			data_in_3_65_in_data = data_store_1_28;
		end else if (andOp_521_out) begin 
			data_in_3_65_in_data = data_store_2_46;
		end else if (andOp_523_out) begin 
			data_in_3_65_in_data = data_store_3_64;
		end else if (andOp_525_out) begin 
			data_in_3_65_in_data = data_store_4_82;
		end else begin
			data_in_3_65_in_data = 0;
		end
	end
	// controller for data_in_3_67.data_in_3_67_in_data
	always @(*) begin
		if (andOp_517_out) begin 
			data_in_3_67_in_data = data_store_0_12;
		end else if (andOp_519_out) begin 
			data_in_3_67_in_data = data_store_1_30;
		end else if (andOp_521_out) begin 
			data_in_3_67_in_data = data_store_2_48;
		end else if (andOp_523_out) begin 
			data_in_3_67_in_data = data_store_3_66;
		end else if (andOp_525_out) begin 
			data_in_3_67_in_data = data_store_4_84;
		end else begin
			data_in_3_67_in_data = 0;
		end
	end
	// controller for data_in_3_69.data_in_3_69_in_data
	always @(*) begin
		if (andOp_517_out) begin 
			data_in_3_69_in_data = data_store_0_14;
		end else if (andOp_519_out) begin 
			data_in_3_69_in_data = data_store_1_32;
		end else if (andOp_521_out) begin 
			data_in_3_69_in_data = data_store_2_50;
		end else if (andOp_523_out) begin 
			data_in_3_69_in_data = data_store_3_68;
		end else if (andOp_525_out) begin 
			data_in_3_69_in_data = data_store_4_86;
		end else begin
			data_in_3_69_in_data = 0;
		end
	end
	// controller for data_in_3_71.data_in_3_71_in_data
	always @(*) begin
		if (andOp_517_out) begin 
			data_in_3_71_in_data = data_store_0_16;
		end else if (andOp_519_out) begin 
			data_in_3_71_in_data = data_store_1_34;
		end else if (andOp_521_out) begin 
			data_in_3_71_in_data = data_store_2_52;
		end else if (andOp_523_out) begin 
			data_in_3_71_in_data = data_store_3_70;
		end else if (andOp_525_out) begin 
			data_in_3_71_in_data = data_store_4_88;
		end else begin
			data_in_3_71_in_data = 0;
		end
	end
	// controller for data_in_4_73.data_in_4_73_in_data
	always @(*) begin
		if (andOp_608_out) begin 
			data_in_4_73_in_data = data_store_0_0;
		end else if (andOp_610_out) begin 
			data_in_4_73_in_data = data_store_1_18;
		end else if (andOp_612_out) begin 
			data_in_4_73_in_data = data_store_2_36;
		end else if (andOp_614_out) begin 
			data_in_4_73_in_data = data_store_3_54;
		end else if (andOp_616_out) begin 
			data_in_4_73_in_data = data_store_4_72;
		end else begin
			data_in_4_73_in_data = 0;
		end
	end
	// controller for data_in_4_75.data_in_4_75_in_data
	always @(*) begin
		if (andOp_608_out) begin 
			data_in_4_75_in_data = data_store_0_2;
		end else if (andOp_610_out) begin 
			data_in_4_75_in_data = data_store_1_20;
		end else if (andOp_612_out) begin 
			data_in_4_75_in_data = data_store_2_38;
		end else if (andOp_614_out) begin 
			data_in_4_75_in_data = data_store_3_56;
		end else if (andOp_616_out) begin 
			data_in_4_75_in_data = data_store_4_74;
		end else begin
			data_in_4_75_in_data = 0;
		end
	end
	// controller for data_in_4_77.data_in_4_77_in_data
	always @(*) begin
		if (andOp_608_out) begin 
			data_in_4_77_in_data = data_store_0_4;
		end else if (andOp_610_out) begin 
			data_in_4_77_in_data = data_store_1_22;
		end else if (andOp_612_out) begin 
			data_in_4_77_in_data = data_store_2_40;
		end else if (andOp_614_out) begin 
			data_in_4_77_in_data = data_store_3_58;
		end else if (andOp_616_out) begin 
			data_in_4_77_in_data = data_store_4_76;
		end else begin
			data_in_4_77_in_data = 0;
		end
	end
	// controller for data_in_4_79.data_in_4_79_in_data
	always @(*) begin
		if (andOp_608_out) begin 
			data_in_4_79_in_data = data_store_0_6;
		end else if (andOp_610_out) begin 
			data_in_4_79_in_data = data_store_1_24;
		end else if (andOp_612_out) begin 
			data_in_4_79_in_data = data_store_2_42;
		end else if (andOp_614_out) begin 
			data_in_4_79_in_data = data_store_3_60;
		end else if (andOp_616_out) begin 
			data_in_4_79_in_data = data_store_4_78;
		end else begin
			data_in_4_79_in_data = 0;
		end
	end
	// controller for data_in_4_81.data_in_4_81_in_data
	always @(*) begin
		if (andOp_608_out) begin 
			data_in_4_81_in_data = data_store_0_8;
		end else if (andOp_610_out) begin 
			data_in_4_81_in_data = data_store_1_26;
		end else if (andOp_612_out) begin 
			data_in_4_81_in_data = data_store_2_44;
		end else if (andOp_614_out) begin 
			data_in_4_81_in_data = data_store_3_62;
		end else if (andOp_616_out) begin 
			data_in_4_81_in_data = data_store_4_80;
		end else begin
			data_in_4_81_in_data = 0;
		end
	end
	// controller for data_in_4_83.data_in_4_83_in_data
	always @(*) begin
		if (andOp_608_out) begin 
			data_in_4_83_in_data = data_store_0_10;
		end else if (andOp_610_out) begin 
			data_in_4_83_in_data = data_store_1_28;
		end else if (andOp_612_out) begin 
			data_in_4_83_in_data = data_store_2_46;
		end else if (andOp_614_out) begin 
			data_in_4_83_in_data = data_store_3_64;
		end else if (andOp_616_out) begin 
			data_in_4_83_in_data = data_store_4_82;
		end else begin
			data_in_4_83_in_data = 0;
		end
	end
	// controller for data_in_4_85.data_in_4_85_in_data
	always @(*) begin
		if (andOp_608_out) begin 
			data_in_4_85_in_data = data_store_0_12;
		end else if (andOp_610_out) begin 
			data_in_4_85_in_data = data_store_1_30;
		end else if (andOp_612_out) begin 
			data_in_4_85_in_data = data_store_2_48;
		end else if (andOp_614_out) begin 
			data_in_4_85_in_data = data_store_3_66;
		end else if (andOp_616_out) begin 
			data_in_4_85_in_data = data_store_4_84;
		end else begin
			data_in_4_85_in_data = 0;
		end
	end
	// controller for data_in_4_87.data_in_4_87_in_data
	always @(*) begin
		if (andOp_608_out) begin 
			data_in_4_87_in_data = data_store_0_14;
		end else if (andOp_610_out) begin 
			data_in_4_87_in_data = data_store_1_32;
		end else if (andOp_612_out) begin 
			data_in_4_87_in_data = data_store_2_50;
		end else if (andOp_614_out) begin 
			data_in_4_87_in_data = data_store_3_68;
		end else if (andOp_616_out) begin 
			data_in_4_87_in_data = data_store_4_86;
		end else begin
			data_in_4_87_in_data = 0;
		end
	end
	// controller for data_in_4_89.data_in_4_89_in_data
	always @(*) begin
		if (andOp_608_out) begin 
			data_in_4_89_in_data = data_store_0_16;
		end else if (andOp_610_out) begin 
			data_in_4_89_in_data = data_store_1_34;
		end else if (andOp_612_out) begin 
			data_in_4_89_in_data = data_store_2_52;
		end else if (andOp_614_out) begin 
			data_in_4_89_in_data = data_store_3_70;
		end else if (andOp_616_out) begin 
			data_in_4_89_in_data = data_store_4_88;
		end else begin
			data_in_4_89_in_data = 0;
		end
	end
	// controller for eq_141.eq_141_in0
	// controller for eq_141.eq_141_in1
	// Insensitive connections
	always @(*) begin
		eq_141_in0 = valid ? 32'd0 : 32'd0;
		eq_141_in1 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
	end
	// controller for eq_142.eq_142_in0
	// controller for eq_142.eq_142_in1
	// Insensitive connections
	always @(*) begin
		eq_142_in0 = valid ? 32'd8 : 32'd8;
		eq_142_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_144.eq_144_in0
	// controller for eq_144.eq_144_in1
	// Insensitive connections
	always @(*) begin
		eq_144_in0 = valid ? 32'd0 : 32'd0;
		eq_144_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_145.eq_145_in0
	// controller for eq_145.eq_145_in1
	// Insensitive connections
	always @(*) begin
		eq_145_in0 = valid ? 32'd3 : 32'd3;
		eq_145_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_147.eq_147_in0
	// controller for eq_147.eq_147_in1
	// Insensitive connections
	always @(*) begin
		eq_147_in0 = valid ? 32'd9 : 32'd9;
		eq_147_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_149.eq_149_in0
	// controller for eq_149.eq_149_in1
	// Insensitive connections
	always @(*) begin
		eq_149_in0 = valid ? 32'd10 : 32'd10;
		eq_149_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_150.eq_150_in0
	// controller for eq_150.eq_150_in1
	// Insensitive connections
	always @(*) begin
		eq_150_in0 = valid ? 32'd4 : 32'd4;
		eq_150_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_152.eq_152_in0
	// controller for eq_152.eq_152_in1
	// Insensitive connections
	always @(*) begin
		eq_152_in0 = valid ? 32'd10 : 32'd10;
		eq_152_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_153.eq_153_in0
	// controller for eq_153.eq_153_in1
	// Insensitive connections
	always @(*) begin
		eq_153_in0 = valid ? 32'd5 : 32'd5;
		eq_153_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_155.eq_155_in0
	// controller for eq_155.eq_155_in1
	// Insensitive connections
	always @(*) begin
		eq_155_in0 = valid ? 32'd6 : 32'd6;
		eq_155_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_157.eq_157_in0
	// controller for eq_157.eq_157_in1
	// Insensitive connections
	always @(*) begin
		eq_157_in0 = valid ? 32'd7 : 32'd7;
		eq_157_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_159.eq_159_in0
	// controller for eq_159.eq_159_in1
	// Insensitive connections
	always @(*) begin
		eq_159_in0 = valid ? 32'd4 : 32'd4;
		eq_159_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_160.eq_160_in0
	// controller for eq_160.eq_160_in1
	// Insensitive connections
	always @(*) begin
		eq_160_in0 = valid ? 32'd2 : 32'd2;
		eq_160_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_162.eq_162_in0
	// controller for eq_162.eq_162_in1
	// Insensitive connections
	always @(*) begin
		eq_162_in0 = valid ? 32'd1 : 32'd1;
		eq_162_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_164.eq_164_in0
	// controller for eq_164.eq_164_in1
	// Insensitive connections
	always @(*) begin
		eq_164_in0 = valid ? 32'd0 : 32'd0;
		eq_164_in1 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
	end
	// controller for eq_165.eq_165_in0
	// controller for eq_165.eq_165_in1
	// Insensitive connections
	always @(*) begin
		eq_165_in0 = valid ? 32'd8 : 32'd8;
		eq_165_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_168.eq_168_in0
	// controller for eq_168.eq_168_in1
	// Insensitive connections
	always @(*) begin
		eq_168_in0 = valid ? 32'd0 : 32'd0;
		eq_168_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_169.eq_169_in0
	// controller for eq_169.eq_169_in1
	// Insensitive connections
	always @(*) begin
		eq_169_in0 = valid ? 32'd3 : 32'd3;
		eq_169_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_172.eq_172_in0
	// controller for eq_172.eq_172_in1
	// Insensitive connections
	always @(*) begin
		eq_172_in0 = valid ? 32'd9 : 32'd9;
		eq_172_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_175.eq_175_in0
	// controller for eq_175.eq_175_in1
	// Insensitive connections
	always @(*) begin
		eq_175_in0 = valid ? 32'd10 : 32'd10;
		eq_175_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_176.eq_176_in0
	// controller for eq_176.eq_176_in1
	// Insensitive connections
	always @(*) begin
		eq_176_in0 = valid ? 32'd4 : 32'd4;
		eq_176_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_179.eq_179_in0
	// controller for eq_179.eq_179_in1
	// Insensitive connections
	always @(*) begin
		eq_179_in0 = valid ? 32'd10 : 32'd10;
		eq_179_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_180.eq_180_in0
	// controller for eq_180.eq_180_in1
	// Insensitive connections
	always @(*) begin
		eq_180_in0 = valid ? 32'd5 : 32'd5;
		eq_180_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_183.eq_183_in0
	// controller for eq_183.eq_183_in1
	// Insensitive connections
	always @(*) begin
		eq_183_in0 = valid ? 32'd6 : 32'd6;
		eq_183_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_186.eq_186_in0
	// controller for eq_186.eq_186_in1
	// Insensitive connections
	always @(*) begin
		eq_186_in0 = valid ? 32'd7 : 32'd7;
		eq_186_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_189.eq_189_in0
	// controller for eq_189.eq_189_in1
	// Insensitive connections
	always @(*) begin
		eq_189_in0 = valid ? 32'd4 : 32'd4;
		eq_189_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_190.eq_190_in0
	// controller for eq_190.eq_190_in1
	// Insensitive connections
	always @(*) begin
		eq_190_in0 = valid ? 32'd2 : 32'd2;
		eq_190_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_193.eq_193_in0
	// controller for eq_193.eq_193_in1
	// Insensitive connections
	always @(*) begin
		eq_193_in0 = valid ? 32'd1 : 32'd1;
		eq_193_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_211.eq_211_in0
	// controller for eq_211.eq_211_in1
	// Insensitive connections
	always @(*) begin
		eq_211_in0 = valid ? 32'd10 : 32'd10;
		eq_211_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_243.eq_243_in0
	// controller for eq_243.eq_243_in1
	// Insensitive connections
	always @(*) begin
		eq_243_in0 = valid ? 32'd0 : 32'd0;
		eq_243_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_245.eq_245_in0
	// controller for eq_245.eq_245_in1
	// Insensitive connections
	always @(*) begin
		eq_245_in0 = valid ? 32'd1 : 32'd1;
		eq_245_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_247.eq_247_in0
	// controller for eq_247.eq_247_in1
	// Insensitive connections
	always @(*) begin
		eq_247_in0 = valid ? 32'd2 : 32'd2;
		eq_247_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_249.eq_249_in0
	// controller for eq_249.eq_249_in1
	// Insensitive connections
	always @(*) begin
		eq_249_in0 = valid ? 32'd3 : 32'd3;
		eq_249_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_251.eq_251_in0
	// controller for eq_251.eq_251_in1
	// Insensitive connections
	always @(*) begin
		eq_251_in0 = valid ? 32'd4 : 32'd4;
		eq_251_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_254.eq_254_in0
	// controller for eq_254.eq_254_in1
	// Insensitive connections
	always @(*) begin
		eq_254_in0 = valid ? 32'd1 : 32'd1;
		eq_254_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_263.eq_263_in0
	// controller for eq_263.eq_263_in1
	// Insensitive connections
	always @(*) begin
		eq_263_in0 = valid ? 32'd3 : 32'd3;
		eq_263_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_272.eq_272_in0
	// controller for eq_272.eq_272_in1
	// Insensitive connections
	always @(*) begin
		eq_272_in0 = valid ? 32'd1 : 32'd1;
		eq_272_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_281.eq_281_in0
	// controller for eq_281.eq_281_in1
	// Insensitive connections
	always @(*) begin
		eq_281_in0 = valid ? 32'd3 : 32'd3;
		eq_281_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_290.eq_290_in0
	// controller for eq_290.eq_290_in1
	// Insensitive connections
	always @(*) begin
		eq_290_in0 = valid ? 32'd3 : 32'd3;
		eq_290_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_299.eq_299_in0
	// controller for eq_299.eq_299_in1
	// Insensitive connections
	always @(*) begin
		eq_299_in0 = valid ? 32'd3 : 32'd3;
		eq_299_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_308.eq_308_in0
	// controller for eq_308.eq_308_in1
	// Insensitive connections
	always @(*) begin
		eq_308_in0 = valid ? 32'd3 : 32'd3;
		eq_308_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_317.eq_317_in0
	// controller for eq_317.eq_317_in1
	// Insensitive connections
	always @(*) begin
		eq_317_in0 = valid ? 32'd4 : 32'd4;
		eq_317_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_326.eq_326_in0
	// controller for eq_326.eq_326_in1
	// Insensitive connections
	always @(*) begin
		eq_326_in0 = valid ? 32'd4 : 32'd4;
		eq_326_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_334.eq_334_in0
	// controller for eq_334.eq_334_in1
	// Insensitive connections
	always @(*) begin
		eq_334_in0 = valid ? 32'd0 : 32'd0;
		eq_334_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_336.eq_336_in0
	// controller for eq_336.eq_336_in1
	// Insensitive connections
	always @(*) begin
		eq_336_in0 = valid ? 32'd1 : 32'd1;
		eq_336_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_338.eq_338_in0
	// controller for eq_338.eq_338_in1
	// Insensitive connections
	always @(*) begin
		eq_338_in0 = valid ? 32'd2 : 32'd2;
		eq_338_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_340.eq_340_in0
	// controller for eq_340.eq_340_in1
	// Insensitive connections
	always @(*) begin
		eq_340_in0 = valid ? 32'd3 : 32'd3;
		eq_340_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_342.eq_342_in0
	// controller for eq_342.eq_342_in1
	// Insensitive connections
	always @(*) begin
		eq_342_in0 = valid ? 32'd4 : 32'd4;
		eq_342_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_345.eq_345_in0
	// controller for eq_345.eq_345_in1
	// Insensitive connections
	always @(*) begin
		eq_345_in0 = valid ? 32'd1 : 32'd1;
		eq_345_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_354.eq_354_in0
	// controller for eq_354.eq_354_in1
	// Insensitive connections
	always @(*) begin
		eq_354_in0 = valid ? 32'd3 : 32'd3;
		eq_354_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_363.eq_363_in0
	// controller for eq_363.eq_363_in1
	// Insensitive connections
	always @(*) begin
		eq_363_in0 = valid ? 32'd1 : 32'd1;
		eq_363_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_372.eq_372_in0
	// controller for eq_372.eq_372_in1
	// Insensitive connections
	always @(*) begin
		eq_372_in0 = valid ? 32'd3 : 32'd3;
		eq_372_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_381.eq_381_in0
	// controller for eq_381.eq_381_in1
	// Insensitive connections
	always @(*) begin
		eq_381_in0 = valid ? 32'd3 : 32'd3;
		eq_381_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_390.eq_390_in0
	// controller for eq_390.eq_390_in1
	// Insensitive connections
	always @(*) begin
		eq_390_in0 = valid ? 32'd3 : 32'd3;
		eq_390_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_399.eq_399_in0
	// controller for eq_399.eq_399_in1
	// Insensitive connections
	always @(*) begin
		eq_399_in0 = valid ? 32'd3 : 32'd3;
		eq_399_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_408.eq_408_in0
	// controller for eq_408.eq_408_in1
	// Insensitive connections
	always @(*) begin
		eq_408_in0 = valid ? 32'd4 : 32'd4;
		eq_408_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_417.eq_417_in0
	// controller for eq_417.eq_417_in1
	// Insensitive connections
	always @(*) begin
		eq_417_in0 = valid ? 32'd4 : 32'd4;
		eq_417_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_425.eq_425_in0
	// controller for eq_425.eq_425_in1
	// Insensitive connections
	always @(*) begin
		eq_425_in0 = valid ? 32'd0 : 32'd0;
		eq_425_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_427.eq_427_in0
	// controller for eq_427.eq_427_in1
	// Insensitive connections
	always @(*) begin
		eq_427_in0 = valid ? 32'd1 : 32'd1;
		eq_427_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_429.eq_429_in0
	// controller for eq_429.eq_429_in1
	// Insensitive connections
	always @(*) begin
		eq_429_in0 = valid ? 32'd2 : 32'd2;
		eq_429_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_431.eq_431_in0
	// controller for eq_431.eq_431_in1
	// Insensitive connections
	always @(*) begin
		eq_431_in0 = valid ? 32'd3 : 32'd3;
		eq_431_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_433.eq_433_in0
	// controller for eq_433.eq_433_in1
	// Insensitive connections
	always @(*) begin
		eq_433_in0 = valid ? 32'd4 : 32'd4;
		eq_433_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_436.eq_436_in0
	// controller for eq_436.eq_436_in1
	// Insensitive connections
	always @(*) begin
		eq_436_in0 = valid ? 32'd1 : 32'd1;
		eq_436_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_445.eq_445_in0
	// controller for eq_445.eq_445_in1
	// Insensitive connections
	always @(*) begin
		eq_445_in0 = valid ? 32'd3 : 32'd3;
		eq_445_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_454.eq_454_in0
	// controller for eq_454.eq_454_in1
	// Insensitive connections
	always @(*) begin
		eq_454_in0 = valid ? 32'd1 : 32'd1;
		eq_454_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_463.eq_463_in0
	// controller for eq_463.eq_463_in1
	// Insensitive connections
	always @(*) begin
		eq_463_in0 = valid ? 32'd3 : 32'd3;
		eq_463_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_472.eq_472_in0
	// controller for eq_472.eq_472_in1
	// Insensitive connections
	always @(*) begin
		eq_472_in0 = valid ? 32'd3 : 32'd3;
		eq_472_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_481.eq_481_in0
	// controller for eq_481.eq_481_in1
	// Insensitive connections
	always @(*) begin
		eq_481_in0 = valid ? 32'd3 : 32'd3;
		eq_481_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_490.eq_490_in0
	// controller for eq_490.eq_490_in1
	// Insensitive connections
	always @(*) begin
		eq_490_in0 = valid ? 32'd3 : 32'd3;
		eq_490_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_499.eq_499_in0
	// controller for eq_499.eq_499_in1
	// Insensitive connections
	always @(*) begin
		eq_499_in0 = valid ? 32'd4 : 32'd4;
		eq_499_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_508.eq_508_in0
	// controller for eq_508.eq_508_in1
	// Insensitive connections
	always @(*) begin
		eq_508_in0 = valid ? 32'd4 : 32'd4;
		eq_508_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_516.eq_516_in0
	// controller for eq_516.eq_516_in1
	// Insensitive connections
	always @(*) begin
		eq_516_in0 = valid ? 32'd0 : 32'd0;
		eq_516_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_518.eq_518_in0
	// controller for eq_518.eq_518_in1
	// Insensitive connections
	always @(*) begin
		eq_518_in0 = valid ? 32'd1 : 32'd1;
		eq_518_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_520.eq_520_in0
	// controller for eq_520.eq_520_in1
	// Insensitive connections
	always @(*) begin
		eq_520_in0 = valid ? 32'd2 : 32'd2;
		eq_520_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_522.eq_522_in0
	// controller for eq_522.eq_522_in1
	// Insensitive connections
	always @(*) begin
		eq_522_in0 = valid ? 32'd3 : 32'd3;
		eq_522_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_524.eq_524_in0
	// controller for eq_524.eq_524_in1
	// Insensitive connections
	always @(*) begin
		eq_524_in0 = valid ? 32'd4 : 32'd4;
		eq_524_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_527.eq_527_in0
	// controller for eq_527.eq_527_in1
	// Insensitive connections
	always @(*) begin
		eq_527_in0 = valid ? 32'd1 : 32'd1;
		eq_527_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_536.eq_536_in0
	// controller for eq_536.eq_536_in1
	// Insensitive connections
	always @(*) begin
		eq_536_in0 = valid ? 32'd3 : 32'd3;
		eq_536_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_545.eq_545_in0
	// controller for eq_545.eq_545_in1
	// Insensitive connections
	always @(*) begin
		eq_545_in0 = valid ? 32'd1 : 32'd1;
		eq_545_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_554.eq_554_in0
	// controller for eq_554.eq_554_in1
	// Insensitive connections
	always @(*) begin
		eq_554_in0 = valid ? 32'd3 : 32'd3;
		eq_554_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_563.eq_563_in0
	// controller for eq_563.eq_563_in1
	// Insensitive connections
	always @(*) begin
		eq_563_in0 = valid ? 32'd3 : 32'd3;
		eq_563_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_572.eq_572_in0
	// controller for eq_572.eq_572_in1
	// Insensitive connections
	always @(*) begin
		eq_572_in0 = valid ? 32'd3 : 32'd3;
		eq_572_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_581.eq_581_in0
	// controller for eq_581.eq_581_in1
	// Insensitive connections
	always @(*) begin
		eq_581_in0 = valid ? 32'd3 : 32'd3;
		eq_581_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_590.eq_590_in0
	// controller for eq_590.eq_590_in1
	// Insensitive connections
	always @(*) begin
		eq_590_in0 = valid ? 32'd4 : 32'd4;
		eq_590_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_599.eq_599_in0
	// controller for eq_599.eq_599_in1
	// Insensitive connections
	always @(*) begin
		eq_599_in0 = valid ? 32'd4 : 32'd4;
		eq_599_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_607.eq_607_in0
	// controller for eq_607.eq_607_in1
	// Insensitive connections
	always @(*) begin
		eq_607_in0 = valid ? 32'd0 : 32'd0;
		eq_607_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_609.eq_609_in0
	// controller for eq_609.eq_609_in1
	// Insensitive connections
	always @(*) begin
		eq_609_in0 = valid ? 32'd1 : 32'd1;
		eq_609_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_611.eq_611_in0
	// controller for eq_611.eq_611_in1
	// Insensitive connections
	always @(*) begin
		eq_611_in0 = valid ? 32'd2 : 32'd2;
		eq_611_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_613.eq_613_in0
	// controller for eq_613.eq_613_in1
	// Insensitive connections
	always @(*) begin
		eq_613_in0 = valid ? 32'd3 : 32'd3;
		eq_613_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_615.eq_615_in0
	// controller for eq_615.eq_615_in1
	// Insensitive connections
	always @(*) begin
		eq_615_in0 = valid ? 32'd4 : 32'd4;
		eq_615_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_618.eq_618_in0
	// controller for eq_618.eq_618_in1
	// Insensitive connections
	always @(*) begin
		eq_618_in0 = valid ? 32'd1 : 32'd1;
		eq_618_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_627.eq_627_in0
	// controller for eq_627.eq_627_in1
	// Insensitive connections
	always @(*) begin
		eq_627_in0 = valid ? 32'd3 : 32'd3;
		eq_627_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_636.eq_636_in0
	// controller for eq_636.eq_636_in1
	// Insensitive connections
	always @(*) begin
		eq_636_in0 = valid ? 32'd1 : 32'd1;
		eq_636_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_645.eq_645_in0
	// controller for eq_645.eq_645_in1
	// Insensitive connections
	always @(*) begin
		eq_645_in0 = valid ? 32'd3 : 32'd3;
		eq_645_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_654.eq_654_in0
	// controller for eq_654.eq_654_in1
	// Insensitive connections
	always @(*) begin
		eq_654_in0 = valid ? 32'd3 : 32'd3;
		eq_654_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_663.eq_663_in0
	// controller for eq_663.eq_663_in1
	// Insensitive connections
	always @(*) begin
		eq_663_in0 = valid ? 32'd3 : 32'd3;
		eq_663_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_672.eq_672_in0
	// controller for eq_672.eq_672_in1
	// Insensitive connections
	always @(*) begin
		eq_672_in0 = valid ? 32'd3 : 32'd3;
		eq_672_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_681.eq_681_in0
	// controller for eq_681.eq_681_in1
	// Insensitive connections
	always @(*) begin
		eq_681_in0 = valid ? 32'd4 : 32'd4;
		eq_681_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_690.eq_690_in0
	// controller for eq_690.eq_690_in1
	// Insensitive connections
	always @(*) begin
		eq_690_in0 = valid ? 32'd4 : 32'd4;
		eq_690_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for icmp_17.cmp_in0_icmp_17
	// controller for icmp_17.cmp_in1_icmp_17
	// Insensitive connections
	always @(*) begin
		cmp_in0_icmp_17 = valid ? add_out_add_16 : add_out_add_16;
		cmp_in1_icmp_17 = valid ? 32'd4 : 32'd4;
	end
	// controller for in.in_read_valid_reg
	always @(*) begin
		if (andOp_204_out) begin 
			in_read_valid_reg = -(1'd1);
		end else begin
			in_read_valid_reg = 0;
		end
	end
	// controller for notOp_101.notOp_101_in0
	// Insensitive connections
	always @(*) begin
		notOp_101_in0 = valid ? andOp_100_out : andOp_100_out;
	end
	// controller for notOp_104.notOp_104_in0
	// Insensitive connections
	always @(*) begin
		notOp_104_in0 = valid ? andOp_103_out : andOp_103_out;
	end
	// controller for notOp_106.notOp_106_in0
	// Insensitive connections
	always @(*) begin
		notOp_106_in0 = valid ? in_read_ready : in_read_ready;
	end
	// controller for notOp_110.notOp_110_in0
	// Insensitive connections
	always @(*) begin
		notOp_110_in0 = valid ? andOp_109_out : andOp_109_out;
	end
	// controller for notOp_113.notOp_113_in0
	// Insensitive connections
	always @(*) begin
		notOp_113_in0 = valid ? andOp_112_out : andOp_112_out;
	end
	// controller for notOp_115.notOp_115_in0
	// Insensitive connections
	always @(*) begin
		notOp_115_in0 = valid ? data_in_4_85_out_data : data_in_4_85_out_data;
	end
	// controller for notOp_119.notOp_119_in0
	// Insensitive connections
	always @(*) begin
		notOp_119_in0 = valid ? andOp_118_out : andOp_118_out;
	end
	// controller for notOp_122.notOp_122_in0
	// Insensitive connections
	always @(*) begin
		notOp_122_in0 = valid ? andOp_121_out : andOp_121_out;
	end
	// controller for notOp_125.notOp_125_in0
	// Insensitive connections
	always @(*) begin
		notOp_125_in0 = valid ? andOp_124_out : andOp_124_out;
	end
	// controller for notOp_127.notOp_127_in0
	// Insensitive connections
	always @(*) begin
		notOp_127_in0 = valid ? out_write_ready : out_write_ready;
	end
	// controller for notOp_131.notOp_131_in0
	// Insensitive connections
	always @(*) begin
		notOp_131_in0 = valid ? andOp_130_out : andOp_130_out;
	end
	// controller for notOp_134.notOp_134_in0
	// Insensitive connections
	always @(*) begin
		notOp_134_in0 = valid ? andOp_133_out : andOp_133_out;
	end
	// controller for notOp_136.notOp_136_in0
	// Insensitive connections
	always @(*) begin
		notOp_136_in0 = valid ? data_in_4_85_out_data : data_in_4_85_out_data;
	end
	// controller for notOp_140.notOp_140_in0
	// Insensitive connections
	always @(*) begin
		notOp_140_in0 = valid ? andOp_139_out : andOp_139_out;
	end
	// controller for notOp_166.notOp_166_in0
	// Insensitive connections
	always @(*) begin
		notOp_166_in0 = valid ? eq_165_out : eq_165_out;
	end
	// controller for notOp_170.notOp_170_in0
	// Insensitive connections
	always @(*) begin
		notOp_170_in0 = valid ? eq_169_out : eq_169_out;
	end
	// controller for notOp_173.notOp_173_in0
	// Insensitive connections
	always @(*) begin
		notOp_173_in0 = valid ? eq_172_out : eq_172_out;
	end
	// controller for notOp_177.notOp_177_in0
	// Insensitive connections
	always @(*) begin
		notOp_177_in0 = valid ? eq_176_out : eq_176_out;
	end
	// controller for notOp_181.notOp_181_in0
	// Insensitive connections
	always @(*) begin
		notOp_181_in0 = valid ? eq_180_out : eq_180_out;
	end
	// controller for notOp_184.notOp_184_in0
	// Insensitive connections
	always @(*) begin
		notOp_184_in0 = valid ? eq_183_out : eq_183_out;
	end
	// controller for notOp_187.notOp_187_in0
	// Insensitive connections
	always @(*) begin
		notOp_187_in0 = valid ? eq_186_out : eq_186_out;
	end
	// controller for notOp_191.notOp_191_in0
	// Insensitive connections
	always @(*) begin
		notOp_191_in0 = valid ? eq_190_out : eq_190_out;
	end
	// controller for notOp_194.notOp_194_in0
	// Insensitive connections
	always @(*) begin
		notOp_194_in0 = valid ? eq_193_out : eq_193_out;
	end
	// controller for notOp_223.notOp_223_in0
	// Insensitive connections
	always @(*) begin
		notOp_223_in0 = valid ? andOp_107_out : andOp_107_out;
	end
	// controller for notOp_225.notOp_225_in0
	// Insensitive connections
	always @(*) begin
		notOp_225_in0 = valid ? andOp_116_out : andOp_116_out;
	end
	// controller for notOp_227.notOp_227_in0
	// Insensitive connections
	always @(*) begin
		notOp_227_in0 = valid ? andOp_219_out : andOp_219_out;
	end
	// controller for notOp_229.notOp_229_in0
	// Insensitive connections
	always @(*) begin
		notOp_229_in0 = valid ? andOp_105_out : andOp_105_out;
	end
	// controller for notOp_231.notOp_231_in0
	// Insensitive connections
	always @(*) begin
		notOp_231_in0 = valid ? andOp_220_out : andOp_220_out;
	end
	// controller for notOp_233.notOp_233_in0
	// Insensitive connections
	always @(*) begin
		notOp_233_in0 = valid ? andOp_128_out : andOp_128_out;
	end
	// controller for notOp_235.notOp_235_in0
	// Insensitive connections
	always @(*) begin
		notOp_235_in0 = valid ? andOp_221_out : andOp_221_out;
	end
	// controller for notOp_237.notOp_237_in0
	// Insensitive connections
	always @(*) begin
		notOp_237_in0 = valid ? andOp_222_out : andOp_222_out;
	end
	// controller for notOp_256.notOp_256_in0
	// Insensitive connections
	always @(*) begin
		notOp_256_in0 = valid ? eq_254_out : eq_254_out;
	end
	// controller for notOp_258.notOp_258_in0
	// Insensitive connections
	always @(*) begin
		notOp_258_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_260.notOp_260_in0
	// Insensitive connections
	always @(*) begin
		notOp_260_in0 = valid ? andOp_255_out : andOp_255_out;
	end
	// controller for notOp_265.notOp_265_in0
	// Insensitive connections
	always @(*) begin
		notOp_265_in0 = valid ? eq_263_out : eq_263_out;
	end
	// controller for notOp_267.notOp_267_in0
	// Insensitive connections
	always @(*) begin
		notOp_267_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_269.notOp_269_in0
	// Insensitive connections
	always @(*) begin
		notOp_269_in0 = valid ? andOp_264_out : andOp_264_out;
	end
	// controller for notOp_274.notOp_274_in0
	// Insensitive connections
	always @(*) begin
		notOp_274_in0 = valid ? eq_272_out : eq_272_out;
	end
	// controller for notOp_276.notOp_276_in0
	// Insensitive connections
	always @(*) begin
		notOp_276_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_278.notOp_278_in0
	// Insensitive connections
	always @(*) begin
		notOp_278_in0 = valid ? andOp_273_out : andOp_273_out;
	end
	// controller for notOp_283.notOp_283_in0
	// Insensitive connections
	always @(*) begin
		notOp_283_in0 = valid ? eq_281_out : eq_281_out;
	end
	// controller for notOp_285.notOp_285_in0
	// Insensitive connections
	always @(*) begin
		notOp_285_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_287.notOp_287_in0
	// Insensitive connections
	always @(*) begin
		notOp_287_in0 = valid ? andOp_282_out : andOp_282_out;
	end
	// controller for notOp_292.notOp_292_in0
	// Insensitive connections
	always @(*) begin
		notOp_292_in0 = valid ? eq_290_out : eq_290_out;
	end
	// controller for notOp_294.notOp_294_in0
	// Insensitive connections
	always @(*) begin
		notOp_294_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_296.notOp_296_in0
	// Insensitive connections
	always @(*) begin
		notOp_296_in0 = valid ? andOp_291_out : andOp_291_out;
	end
	// controller for notOp_301.notOp_301_in0
	// Insensitive connections
	always @(*) begin
		notOp_301_in0 = valid ? eq_299_out : eq_299_out;
	end
	// controller for notOp_303.notOp_303_in0
	// Insensitive connections
	always @(*) begin
		notOp_303_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_305.notOp_305_in0
	// Insensitive connections
	always @(*) begin
		notOp_305_in0 = valid ? andOp_300_out : andOp_300_out;
	end
	// controller for notOp_310.notOp_310_in0
	// Insensitive connections
	always @(*) begin
		notOp_310_in0 = valid ? eq_308_out : eq_308_out;
	end
	// controller for notOp_312.notOp_312_in0
	// Insensitive connections
	always @(*) begin
		notOp_312_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_314.notOp_314_in0
	// Insensitive connections
	always @(*) begin
		notOp_314_in0 = valid ? andOp_309_out : andOp_309_out;
	end
	// controller for notOp_319.notOp_319_in0
	// Insensitive connections
	always @(*) begin
		notOp_319_in0 = valid ? eq_317_out : eq_317_out;
	end
	// controller for notOp_321.notOp_321_in0
	// Insensitive connections
	always @(*) begin
		notOp_321_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_323.notOp_323_in0
	// Insensitive connections
	always @(*) begin
		notOp_323_in0 = valid ? andOp_318_out : andOp_318_out;
	end
	// controller for notOp_328.notOp_328_in0
	// Insensitive connections
	always @(*) begin
		notOp_328_in0 = valid ? eq_326_out : eq_326_out;
	end
	// controller for notOp_330.notOp_330_in0
	// Insensitive connections
	always @(*) begin
		notOp_330_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_332.notOp_332_in0
	// Insensitive connections
	always @(*) begin
		notOp_332_in0 = valid ? andOp_327_out : andOp_327_out;
	end
	// controller for notOp_347.notOp_347_in0
	// Insensitive connections
	always @(*) begin
		notOp_347_in0 = valid ? eq_345_out : eq_345_out;
	end
	// controller for notOp_349.notOp_349_in0
	// Insensitive connections
	always @(*) begin
		notOp_349_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
	end
	// controller for notOp_351.notOp_351_in0
	// Insensitive connections
	always @(*) begin
		notOp_351_in0 = valid ? andOp_346_out : andOp_346_out;
	end
	// controller for notOp_356.notOp_356_in0
	// Insensitive connections
	always @(*) begin
		notOp_356_in0 = valid ? eq_354_out : eq_354_out;
	end
	// controller for notOp_358.notOp_358_in0
	// Insensitive connections
	always @(*) begin
		notOp_358_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_360.notOp_360_in0
	// Insensitive connections
	always @(*) begin
		notOp_360_in0 = valid ? andOp_355_out : andOp_355_out;
	end
	// controller for notOp_365.notOp_365_in0
	// Insensitive connections
	always @(*) begin
		notOp_365_in0 = valid ? eq_363_out : eq_363_out;
	end
	// controller for notOp_367.notOp_367_in0
	// Insensitive connections
	always @(*) begin
		notOp_367_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
	end
	// controller for notOp_369.notOp_369_in0
	// Insensitive connections
	always @(*) begin
		notOp_369_in0 = valid ? andOp_364_out : andOp_364_out;
	end
	// controller for notOp_374.notOp_374_in0
	// Insensitive connections
	always @(*) begin
		notOp_374_in0 = valid ? eq_372_out : eq_372_out;
	end
	// controller for notOp_376.notOp_376_in0
	// Insensitive connections
	always @(*) begin
		notOp_376_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_378.notOp_378_in0
	// Insensitive connections
	always @(*) begin
		notOp_378_in0 = valid ? andOp_373_out : andOp_373_out;
	end
	// controller for notOp_383.notOp_383_in0
	// Insensitive connections
	always @(*) begin
		notOp_383_in0 = valid ? eq_381_out : eq_381_out;
	end
	// controller for notOp_385.notOp_385_in0
	// Insensitive connections
	always @(*) begin
		notOp_385_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_387.notOp_387_in0
	// Insensitive connections
	always @(*) begin
		notOp_387_in0 = valid ? andOp_382_out : andOp_382_out;
	end
	// controller for notOp_392.notOp_392_in0
	// Insensitive connections
	always @(*) begin
		notOp_392_in0 = valid ? eq_390_out : eq_390_out;
	end
	// controller for notOp_394.notOp_394_in0
	// Insensitive connections
	always @(*) begin
		notOp_394_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_396.notOp_396_in0
	// Insensitive connections
	always @(*) begin
		notOp_396_in0 = valid ? andOp_391_out : andOp_391_out;
	end
	// controller for notOp_401.notOp_401_in0
	// Insensitive connections
	always @(*) begin
		notOp_401_in0 = valid ? eq_399_out : eq_399_out;
	end
	// controller for notOp_403.notOp_403_in0
	// Insensitive connections
	always @(*) begin
		notOp_403_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_405.notOp_405_in0
	// Insensitive connections
	always @(*) begin
		notOp_405_in0 = valid ? andOp_400_out : andOp_400_out;
	end
	// controller for notOp_410.notOp_410_in0
	// Insensitive connections
	always @(*) begin
		notOp_410_in0 = valid ? eq_408_out : eq_408_out;
	end
	// controller for notOp_412.notOp_412_in0
	// Insensitive connections
	always @(*) begin
		notOp_412_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_414.notOp_414_in0
	// Insensitive connections
	always @(*) begin
		notOp_414_in0 = valid ? andOp_409_out : andOp_409_out;
	end
	// controller for notOp_419.notOp_419_in0
	// Insensitive connections
	always @(*) begin
		notOp_419_in0 = valid ? eq_417_out : eq_417_out;
	end
	// controller for notOp_421.notOp_421_in0
	// Insensitive connections
	always @(*) begin
		notOp_421_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_423.notOp_423_in0
	// Insensitive connections
	always @(*) begin
		notOp_423_in0 = valid ? andOp_418_out : andOp_418_out;
	end
	// controller for notOp_438.notOp_438_in0
	// Insensitive connections
	always @(*) begin
		notOp_438_in0 = valid ? eq_436_out : eq_436_out;
	end
	// controller for notOp_440.notOp_440_in0
	// Insensitive connections
	always @(*) begin
		notOp_440_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_442.notOp_442_in0
	// Insensitive connections
	always @(*) begin
		notOp_442_in0 = valid ? andOp_437_out : andOp_437_out;
	end
	// controller for notOp_447.notOp_447_in0
	// Insensitive connections
	always @(*) begin
		notOp_447_in0 = valid ? eq_445_out : eq_445_out;
	end
	// controller for notOp_449.notOp_449_in0
	// Insensitive connections
	always @(*) begin
		notOp_449_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
	end
	// controller for notOp_451.notOp_451_in0
	// Insensitive connections
	always @(*) begin
		notOp_451_in0 = valid ? andOp_446_out : andOp_446_out;
	end
	// controller for notOp_456.notOp_456_in0
	// Insensitive connections
	always @(*) begin
		notOp_456_in0 = valid ? eq_454_out : eq_454_out;
	end
	// controller for notOp_458.notOp_458_in0
	// Insensitive connections
	always @(*) begin
		notOp_458_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_460.notOp_460_in0
	// Insensitive connections
	always @(*) begin
		notOp_460_in0 = valid ? andOp_455_out : andOp_455_out;
	end
	// controller for notOp_465.notOp_465_in0
	// Insensitive connections
	always @(*) begin
		notOp_465_in0 = valid ? eq_463_out : eq_463_out;
	end
	// controller for notOp_467.notOp_467_in0
	// Insensitive connections
	always @(*) begin
		notOp_467_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_469.notOp_469_in0
	// Insensitive connections
	always @(*) begin
		notOp_469_in0 = valid ? andOp_464_out : andOp_464_out;
	end
	// controller for notOp_474.notOp_474_in0
	// Insensitive connections
	always @(*) begin
		notOp_474_in0 = valid ? eq_472_out : eq_472_out;
	end
	// controller for notOp_476.notOp_476_in0
	// Insensitive connections
	always @(*) begin
		notOp_476_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_478.notOp_478_in0
	// Insensitive connections
	always @(*) begin
		notOp_478_in0 = valid ? andOp_473_out : andOp_473_out;
	end
	// controller for notOp_483.notOp_483_in0
	// Insensitive connections
	always @(*) begin
		notOp_483_in0 = valid ? eq_481_out : eq_481_out;
	end
	// controller for notOp_485.notOp_485_in0
	// Insensitive connections
	always @(*) begin
		notOp_485_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_487.notOp_487_in0
	// Insensitive connections
	always @(*) begin
		notOp_487_in0 = valid ? andOp_482_out : andOp_482_out;
	end
	// controller for notOp_492.notOp_492_in0
	// Insensitive connections
	always @(*) begin
		notOp_492_in0 = valid ? eq_490_out : eq_490_out;
	end
	// controller for notOp_494.notOp_494_in0
	// Insensitive connections
	always @(*) begin
		notOp_494_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_496.notOp_496_in0
	// Insensitive connections
	always @(*) begin
		notOp_496_in0 = valid ? andOp_491_out : andOp_491_out;
	end
	// controller for notOp_501.notOp_501_in0
	// Insensitive connections
	always @(*) begin
		notOp_501_in0 = valid ? eq_499_out : eq_499_out;
	end
	// controller for notOp_503.notOp_503_in0
	// Insensitive connections
	always @(*) begin
		notOp_503_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_505.notOp_505_in0
	// Insensitive connections
	always @(*) begin
		notOp_505_in0 = valid ? andOp_500_out : andOp_500_out;
	end
	// controller for notOp_510.notOp_510_in0
	// Insensitive connections
	always @(*) begin
		notOp_510_in0 = valid ? eq_508_out : eq_508_out;
	end
	// controller for notOp_512.notOp_512_in0
	// Insensitive connections
	always @(*) begin
		notOp_512_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_514.notOp_514_in0
	// Insensitive connections
	always @(*) begin
		notOp_514_in0 = valid ? andOp_509_out : andOp_509_out;
	end
	// controller for notOp_529.notOp_529_in0
	// Insensitive connections
	always @(*) begin
		notOp_529_in0 = valid ? eq_527_out : eq_527_out;
	end
	// controller for notOp_531.notOp_531_in0
	// Insensitive connections
	always @(*) begin
		notOp_531_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_533.notOp_533_in0
	// Insensitive connections
	always @(*) begin
		notOp_533_in0 = valid ? andOp_528_out : andOp_528_out;
	end
	// controller for notOp_538.notOp_538_in0
	// Insensitive connections
	always @(*) begin
		notOp_538_in0 = valid ? eq_536_out : eq_536_out;
	end
	// controller for notOp_540.notOp_540_in0
	// Insensitive connections
	always @(*) begin
		notOp_540_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
	end
	// controller for notOp_542.notOp_542_in0
	// Insensitive connections
	always @(*) begin
		notOp_542_in0 = valid ? andOp_537_out : andOp_537_out;
	end
	// controller for notOp_547.notOp_547_in0
	// Insensitive connections
	always @(*) begin
		notOp_547_in0 = valid ? eq_545_out : eq_545_out;
	end
	// controller for notOp_549.notOp_549_in0
	// Insensitive connections
	always @(*) begin
		notOp_549_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_551.notOp_551_in0
	// Insensitive connections
	always @(*) begin
		notOp_551_in0 = valid ? andOp_546_out : andOp_546_out;
	end
	// controller for notOp_556.notOp_556_in0
	// Insensitive connections
	always @(*) begin
		notOp_556_in0 = valid ? eq_554_out : eq_554_out;
	end
	// controller for notOp_558.notOp_558_in0
	// Insensitive connections
	always @(*) begin
		notOp_558_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
	end
	// controller for notOp_560.notOp_560_in0
	// Insensitive connections
	always @(*) begin
		notOp_560_in0 = valid ? andOp_555_out : andOp_555_out;
	end
	// controller for notOp_565.notOp_565_in0
	// Insensitive connections
	always @(*) begin
		notOp_565_in0 = valid ? eq_563_out : eq_563_out;
	end
	// controller for notOp_567.notOp_567_in0
	// Insensitive connections
	always @(*) begin
		notOp_567_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
	end
	// controller for notOp_569.notOp_569_in0
	// Insensitive connections
	always @(*) begin
		notOp_569_in0 = valid ? andOp_564_out : andOp_564_out;
	end
	// controller for notOp_574.notOp_574_in0
	// Insensitive connections
	always @(*) begin
		notOp_574_in0 = valid ? eq_572_out : eq_572_out;
	end
	// controller for notOp_576.notOp_576_in0
	// Insensitive connections
	always @(*) begin
		notOp_576_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
	end
	// controller for notOp_578.notOp_578_in0
	// Insensitive connections
	always @(*) begin
		notOp_578_in0 = valid ? andOp_573_out : andOp_573_out;
	end
	// controller for notOp_583.notOp_583_in0
	// Insensitive connections
	always @(*) begin
		notOp_583_in0 = valid ? eq_581_out : eq_581_out;
	end
	// controller for notOp_585.notOp_585_in0
	// Insensitive connections
	always @(*) begin
		notOp_585_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
	end
	// controller for notOp_587.notOp_587_in0
	// Insensitive connections
	always @(*) begin
		notOp_587_in0 = valid ? andOp_582_out : andOp_582_out;
	end
	// controller for notOp_592.notOp_592_in0
	// Insensitive connections
	always @(*) begin
		notOp_592_in0 = valid ? eq_590_out : eq_590_out;
	end
	// controller for notOp_594.notOp_594_in0
	// Insensitive connections
	always @(*) begin
		notOp_594_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_596.notOp_596_in0
	// Insensitive connections
	always @(*) begin
		notOp_596_in0 = valid ? andOp_591_out : andOp_591_out;
	end
	// controller for notOp_601.notOp_601_in0
	// Insensitive connections
	always @(*) begin
		notOp_601_in0 = valid ? eq_599_out : eq_599_out;
	end
	// controller for notOp_603.notOp_603_in0
	// Insensitive connections
	always @(*) begin
		notOp_603_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_605.notOp_605_in0
	// Insensitive connections
	always @(*) begin
		notOp_605_in0 = valid ? andOp_600_out : andOp_600_out;
	end
	// controller for notOp_620.notOp_620_in0
	// Insensitive connections
	always @(*) begin
		notOp_620_in0 = valid ? eq_618_out : eq_618_out;
	end
	// controller for notOp_622.notOp_622_in0
	// Insensitive connections
	always @(*) begin
		notOp_622_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_624.notOp_624_in0
	// Insensitive connections
	always @(*) begin
		notOp_624_in0 = valid ? andOp_619_out : andOp_619_out;
	end
	// controller for notOp_629.notOp_629_in0
	// Insensitive connections
	always @(*) begin
		notOp_629_in0 = valid ? eq_627_out : eq_627_out;
	end
	// controller for notOp_631.notOp_631_in0
	// Insensitive connections
	always @(*) begin
		notOp_631_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_633.notOp_633_in0
	// Insensitive connections
	always @(*) begin
		notOp_633_in0 = valid ? andOp_628_out : andOp_628_out;
	end
	// controller for notOp_638.notOp_638_in0
	// Insensitive connections
	always @(*) begin
		notOp_638_in0 = valid ? eq_636_out : eq_636_out;
	end
	// controller for notOp_640.notOp_640_in0
	// Insensitive connections
	always @(*) begin
		notOp_640_in0 = valid ? 1'd0 : 1'd0;
	end
	// controller for notOp_642.notOp_642_in0
	// Insensitive connections
	always @(*) begin
		notOp_642_in0 = valid ? andOp_637_out : andOp_637_out;
	end
	// controller for notOp_647.notOp_647_in0
	// Insensitive connections
	always @(*) begin
		notOp_647_in0 = valid ? eq_645_out : eq_645_out;
	end
	// controller for notOp_649.notOp_649_in0
	// Insensitive connections
	always @(*) begin
		notOp_649_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
	end
	// controller for notOp_651.notOp_651_in0
	// Insensitive connections
	always @(*) begin
		notOp_651_in0 = valid ? andOp_646_out : andOp_646_out;
	end
	// controller for notOp_656.notOp_656_in0
	// Insensitive connections
	always @(*) begin
		notOp_656_in0 = valid ? eq_654_out : eq_654_out;
	end
	// controller for notOp_658.notOp_658_in0
	// Insensitive connections
	always @(*) begin
		notOp_658_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
	end
	// controller for notOp_660.notOp_660_in0
	// Insensitive connections
	always @(*) begin
		notOp_660_in0 = valid ? andOp_655_out : andOp_655_out;
	end
	// controller for notOp_665.notOp_665_in0
	// Insensitive connections
	always @(*) begin
		notOp_665_in0 = valid ? eq_663_out : eq_663_out;
	end
	// controller for notOp_667.notOp_667_in0
	// Insensitive connections
	always @(*) begin
		notOp_667_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
	end
	// controller for notOp_669.notOp_669_in0
	// Insensitive connections
	always @(*) begin
		notOp_669_in0 = valid ? andOp_664_out : andOp_664_out;
	end
	// controller for notOp_674.notOp_674_in0
	// Insensitive connections
	always @(*) begin
		notOp_674_in0 = valid ? eq_672_out : eq_672_out;
	end
	// controller for notOp_676.notOp_676_in0
	// Insensitive connections
	always @(*) begin
		notOp_676_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
	end
	// controller for notOp_678.notOp_678_in0
	// Insensitive connections
	always @(*) begin
		notOp_678_in0 = valid ? andOp_673_out : andOp_673_out;
	end
	// controller for notOp_683.notOp_683_in0
	// Insensitive connections
	always @(*) begin
		notOp_683_in0 = valid ? eq_681_out : eq_681_out;
	end
	// controller for notOp_685.notOp_685_in0
	// Insensitive connections
	always @(*) begin
		notOp_685_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
	end
	// controller for notOp_687.notOp_687_in0
	// Insensitive connections
	always @(*) begin
		notOp_687_in0 = valid ? andOp_682_out : andOp_682_out;
	end
	// controller for notOp_692.notOp_692_in0
	// Insensitive connections
	always @(*) begin
		notOp_692_in0 = valid ? eq_690_out : eq_690_out;
	end
	// controller for notOp_694.notOp_694_in0
	// Insensitive connections
	always @(*) begin
		notOp_694_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
	end
	// controller for notOp_696.notOp_696_in0
	// Insensitive connections
	always @(*) begin
		notOp_696_in0 = valid ? andOp_691_out : andOp_691_out;
	end
	// controller for notOp_92.notOp_92_in0
	// Insensitive connections
	always @(*) begin
		notOp_92_in0 = valid ? andOp_91_out : andOp_91_out;
	end
	// controller for notOp_95.notOp_95_in0
	// Insensitive connections
	always @(*) begin
		notOp_95_in0 = valid ? andOp_94_out : andOp_94_out;
	end
	// controller for notOp_98.notOp_98_in0
	// Insensitive connections
	always @(*) begin
		notOp_98_in0 = valid ? andOp_97_out : andOp_97_out;
	end
	// controller for orOp_143.orOp_143_in0
	// controller for orOp_143.orOp_143_in1
	// Insensitive connections
	always @(*) begin
		orOp_143_in0 = valid ? eq_142_out : eq_142_out;
		orOp_143_in1 = valid ? andOp_100_out : andOp_100_out;
	end
	// controller for orOp_146.orOp_146_in0
	// controller for orOp_146.orOp_146_in1
	// Insensitive connections
	always @(*) begin
		orOp_146_in0 = valid ? eq_145_out : eq_145_out;
		orOp_146_in1 = valid ? andOp_91_out : andOp_91_out;
	end
	// controller for orOp_148.orOp_148_in0
	// controller for orOp_148.orOp_148_in1
	// Insensitive connections
	always @(*) begin
		orOp_148_in0 = valid ? eq_147_out : eq_147_out;
		orOp_148_in1 = valid ? andOp_94_out : andOp_94_out;
	end
	// controller for orOp_151.orOp_151_in0
	// controller for orOp_151.orOp_151_in1
	// Insensitive connections
	always @(*) begin
		orOp_151_in0 = valid ? eq_150_out : eq_150_out;
		orOp_151_in1 = valid ? andOp_109_out : andOp_109_out;
	end
	// controller for orOp_154.orOp_154_in0
	// controller for orOp_154.orOp_154_in1
	// Insensitive connections
	always @(*) begin
		orOp_154_in0 = valid ? eq_153_out : eq_153_out;
		orOp_154_in1 = valid ? andOp_139_out : andOp_139_out;
	end
	// controller for orOp_156.orOp_156_in0
	// controller for orOp_156.orOp_156_in1
	// Insensitive connections
	always @(*) begin
		orOp_156_in0 = valid ? eq_155_out : eq_155_out;
		orOp_156_in1 = valid ? andOp_121_out : andOp_121_out;
	end
	// controller for orOp_158.orOp_158_in0
	// controller for orOp_158.orOp_158_in1
	// Insensitive connections
	always @(*) begin
		orOp_158_in0 = valid ? eq_157_out : eq_157_out;
		orOp_158_in1 = valid ? andOp_126_out : andOp_126_out;
	end
	// controller for orOp_161.orOp_161_in0
	// controller for orOp_161.orOp_161_in1
	// Insensitive connections
	always @(*) begin
		orOp_161_in0 = valid ? eq_160_out : eq_160_out;
		orOp_161_in1 = valid ? andOp_130_out : andOp_130_out;
	end
	// controller for orOp_163.orOp_163_in0
	// controller for orOp_163.orOp_163_in1
	// Insensitive connections
	always @(*) begin
		orOp_163_in0 = valid ? eq_162_out : eq_162_out;
		orOp_163_in1 = valid ? andOp_114_out : andOp_114_out;
	end
	// controller for out.out_in_data_reg
	always @(*) begin
		if (andOp_215_out) begin 
			out_in_data_reg = rdata_ram_0;
		end else begin
			out_in_data_reg = 0;
		end
	end
	// controller for out.out_write_valid_reg
	always @(*) begin
		if (andOp_214_out) begin 
			out_write_valid_reg = -(1'd1);
		end else begin
			out_write_valid_reg = 0;
		end
	end
	// controller for phi_7.phi_in_phi_7
	// controller for phi_7.phi_last_block_phi_7
	// controller for phi_7.phi_s_phi_7
	// Insensitive connections
	always @(*) begin
		phi_in_phi_7 = valid ? concat_207_out : concat_207_out;
		phi_last_block_phi_7 = valid ? bb_3_predecessor_in_state_1_out_data : bb_3_predecessor_in_state_1_out_data;
		phi_s_phi_7 = valid ? concat_208_out : concat_208_out;
	end
	// controller for ram_0.raddr_ram_0_reg
	always @(*) begin
		if (andOp_200_out) begin 
			raddr_ram_0_reg = 32'd0;
		end else if (andOp_202_out) begin 
			raddr_ram_0_reg = 32'd0;
		end else begin
			raddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.waddr_ram_0_reg
	always @(*) begin
		if (andOp_199_out) begin 
			waddr_ram_0_reg = 32'd0;
		end else if (andOp_201_out) begin 
			waddr_ram_0_reg = 32'd0;
		end else begin
			waddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wdata_ram_0_reg
	always @(*) begin
		if (andOp_199_out) begin 
			wdata_ram_0_reg = 32'd0;
		end else if (andOp_201_out) begin 
			wdata_ram_0_reg = add_out_add_14;
		end else begin
			wdata_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wen_ram_0_reg
	always @(*) begin
		if (andOp_199_out) begin 
			wen_ram_0_reg = 1'd1;
		end else if (andOp_201_out) begin 
			wen_ram_0_reg = 1'd1;
		end else begin
			wen_ram_0_reg = 0;
		end
	end
	// controller for ret_23.valid_reg
	always @(*) begin
		if (andOp_218_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// controller for tmp_output_210.tmp_output_210_in_data
	always @(*) begin
		if (eq_211_out) begin 
			tmp_output_210_in_data = in_out_data;
		end else begin
			tmp_output_210_in_data = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			add_tmp_5 <= 0;
		end else begin
			if (andOp_241_out) begin
				add_tmp_5 <= add_out_add_16;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			call_tmp_2 <= 0;
		end else begin
			if (andOp_240_out) begin
				call_tmp_2 <= in_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_0 <= 0;
		end else begin
			if (andOp_255_out) begin
				data_store_0_0 <= in_read_ready;
			end
			if (andOp_261_out) begin
				data_store_0_0 <= data_in_0_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_10 <= 0;
		end else begin
			if (andOp_300_out) begin
				data_store_0_10 <= add_out_add_16;
			end
			if (andOp_306_out) begin
				data_store_0_10 <= data_in_0_11_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_12 <= 0;
		end else begin
			if (andOp_309_out) begin
				data_store_0_12 <= cmp_out_icmp_17;
			end
			if (andOp_315_out) begin
				data_store_0_12 <= data_in_0_13_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_14 <= 0;
		end else begin
			if (andOp_318_out) begin
				data_store_0_14 <= rdata_ram_0;
			end
			if (andOp_324_out) begin
				data_store_0_14 <= data_in_0_15_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_16 <= 0;
		end else begin
			if (andOp_327_out) begin
				data_store_0_16 <= out_write_ready;
			end
			if (andOp_333_out) begin
				data_store_0_16 <= data_in_0_17_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_2 <= 0;
		end else begin
			if (andOp_264_out) begin
				data_store_0_2 <= in_out_data;
			end
			if (andOp_270_out) begin
				data_store_0_2 <= data_in_0_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_4 <= 0;
		end else begin
			if (andOp_273_out) begin
				data_store_0_4 <= phi_out_phi_7;
			end
			if (andOp_279_out) begin
				data_store_0_4 <= data_in_0_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_6 <= 0;
		end else begin
			if (andOp_282_out) begin
				data_store_0_6 <= rdata_ram_0;
			end
			if (andOp_288_out) begin
				data_store_0_6 <= data_in_0_7_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_8 <= 0;
		end else begin
			if (andOp_291_out) begin
				data_store_0_8 <= add_out_add_14;
			end
			if (andOp_297_out) begin
				data_store_0_8 <= data_in_0_9_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_18 <= 0;
		end else begin
			if (andOp_346_out) begin
				data_store_1_18 <= in_read_ready;
			end
			if (andOp_352_out) begin
				data_store_1_18 <= data_in_1_19_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_20 <= 0;
		end else begin
			if (andOp_355_out) begin
				data_store_1_20 <= in_out_data;
			end
			if (andOp_361_out) begin
				data_store_1_20 <= data_in_1_21_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_22 <= 0;
		end else begin
			if (andOp_364_out) begin
				data_store_1_22 <= phi_out_phi_7;
			end
			if (andOp_370_out) begin
				data_store_1_22 <= data_in_1_23_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_24 <= 0;
		end else begin
			if (andOp_373_out) begin
				data_store_1_24 <= rdata_ram_0;
			end
			if (andOp_379_out) begin
				data_store_1_24 <= data_in_1_25_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_26 <= 0;
		end else begin
			if (andOp_382_out) begin
				data_store_1_26 <= add_out_add_14;
			end
			if (andOp_388_out) begin
				data_store_1_26 <= data_in_1_27_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_28 <= 0;
		end else begin
			if (andOp_391_out) begin
				data_store_1_28 <= add_out_add_16;
			end
			if (andOp_397_out) begin
				data_store_1_28 <= data_in_1_29_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_30 <= 0;
		end else begin
			if (andOp_400_out) begin
				data_store_1_30 <= cmp_out_icmp_17;
			end
			if (andOp_406_out) begin
				data_store_1_30 <= data_in_1_31_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_32 <= 0;
		end else begin
			if (andOp_409_out) begin
				data_store_1_32 <= rdata_ram_0;
			end
			if (andOp_415_out) begin
				data_store_1_32 <= data_in_1_33_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_34 <= 0;
		end else begin
			if (andOp_418_out) begin
				data_store_1_34 <= out_write_ready;
			end
			if (andOp_424_out) begin
				data_store_1_34 <= data_in_1_35_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_36 <= 0;
		end else begin
			if (andOp_437_out) begin
				data_store_2_36 <= in_read_ready;
			end
			if (andOp_443_out) begin
				data_store_2_36 <= data_in_2_37_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_38 <= 0;
		end else begin
			if (andOp_446_out) begin
				data_store_2_38 <= in_out_data;
			end
			if (andOp_452_out) begin
				data_store_2_38 <= data_in_2_39_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_40 <= 0;
		end else begin
			if (andOp_455_out) begin
				data_store_2_40 <= phi_out_phi_7;
			end
			if (andOp_461_out) begin
				data_store_2_40 <= data_in_2_41_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_42 <= 0;
		end else begin
			if (andOp_464_out) begin
				data_store_2_42 <= rdata_ram_0;
			end
			if (andOp_470_out) begin
				data_store_2_42 <= data_in_2_43_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_44 <= 0;
		end else begin
			if (andOp_473_out) begin
				data_store_2_44 <= add_out_add_14;
			end
			if (andOp_479_out) begin
				data_store_2_44 <= data_in_2_45_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_46 <= 0;
		end else begin
			if (andOp_482_out) begin
				data_store_2_46 <= add_out_add_16;
			end
			if (andOp_488_out) begin
				data_store_2_46 <= data_in_2_47_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_48 <= 0;
		end else begin
			if (andOp_491_out) begin
				data_store_2_48 <= cmp_out_icmp_17;
			end
			if (andOp_497_out) begin
				data_store_2_48 <= data_in_2_49_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_50 <= 0;
		end else begin
			if (andOp_500_out) begin
				data_store_2_50 <= rdata_ram_0;
			end
			if (andOp_506_out) begin
				data_store_2_50 <= data_in_2_51_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_52 <= 0;
		end else begin
			if (andOp_509_out) begin
				data_store_2_52 <= out_write_ready;
			end
			if (andOp_515_out) begin
				data_store_2_52 <= data_in_2_53_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_54 <= 0;
		end else begin
			if (andOp_528_out) begin
				data_store_3_54 <= in_read_ready;
			end
			if (andOp_534_out) begin
				data_store_3_54 <= data_in_3_55_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_56 <= 0;
		end else begin
			if (andOp_537_out) begin
				data_store_3_56 <= in_out_data;
			end
			if (andOp_543_out) begin
				data_store_3_56 <= data_in_3_57_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_58 <= 0;
		end else begin
			if (andOp_546_out) begin
				data_store_3_58 <= phi_out_phi_7;
			end
			if (andOp_552_out) begin
				data_store_3_58 <= data_in_3_59_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_60 <= 0;
		end else begin
			if (andOp_555_out) begin
				data_store_3_60 <= rdata_ram_0;
			end
			if (andOp_561_out) begin
				data_store_3_60 <= data_in_3_61_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_62 <= 0;
		end else begin
			if (andOp_564_out) begin
				data_store_3_62 <= add_out_add_14;
			end
			if (andOp_570_out) begin
				data_store_3_62 <= data_in_3_63_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_64 <= 0;
		end else begin
			if (andOp_573_out) begin
				data_store_3_64 <= add_out_add_16;
			end
			if (andOp_579_out) begin
				data_store_3_64 <= data_in_3_65_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_66 <= 0;
		end else begin
			if (andOp_582_out) begin
				data_store_3_66 <= cmp_out_icmp_17;
			end
			if (andOp_588_out) begin
				data_store_3_66 <= data_in_3_67_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_68 <= 0;
		end else begin
			if (andOp_591_out) begin
				data_store_3_68 <= rdata_ram_0;
			end
			if (andOp_597_out) begin
				data_store_3_68 <= data_in_3_69_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_70 <= 0;
		end else begin
			if (andOp_600_out) begin
				data_store_3_70 <= out_write_ready;
			end
			if (andOp_606_out) begin
				data_store_3_70 <= data_in_3_71_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_72 <= 0;
		end else begin
			if (andOp_619_out) begin
				data_store_4_72 <= in_read_ready;
			end
			if (andOp_625_out) begin
				data_store_4_72 <= data_in_4_73_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_74 <= 0;
		end else begin
			if (andOp_628_out) begin
				data_store_4_74 <= in_out_data;
			end
			if (andOp_634_out) begin
				data_store_4_74 <= data_in_4_75_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_76 <= 0;
		end else begin
			if (andOp_637_out) begin
				data_store_4_76 <= phi_out_phi_7;
			end
			if (andOp_643_out) begin
				data_store_4_76 <= data_in_4_77_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_78 <= 0;
		end else begin
			if (andOp_646_out) begin
				data_store_4_78 <= rdata_ram_0;
			end
			if (andOp_652_out) begin
				data_store_4_78 <= data_in_4_79_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_80 <= 0;
		end else begin
			if (andOp_655_out) begin
				data_store_4_80 <= add_out_add_14;
			end
			if (andOp_661_out) begin
				data_store_4_80 <= data_in_4_81_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_82 <= 0;
		end else begin
			if (andOp_664_out) begin
				data_store_4_82 <= add_out_add_16;
			end
			if (andOp_670_out) begin
				data_store_4_82 <= data_in_4_83_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_84 <= 0;
		end else begin
			if (andOp_673_out) begin
				data_store_4_84 <= cmp_out_icmp_17;
			end
			if (andOp_679_out) begin
				data_store_4_84 <= data_in_4_85_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_86 <= 0;
		end else begin
			if (andOp_682_out) begin
				data_store_4_86 <= rdata_ram_0;
			end
			if (andOp_688_out) begin
				data_store_4_86 <= data_in_4_87_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_88 <= 0;
		end else begin
			if (andOp_691_out) begin
				data_store_4_88 <= out_write_ready;
			end
			if (andOp_697_out) begin
				data_store_4_88 <= data_in_4_89_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_105_out) begin
				global_state <= 32'd2;
			end
			if (andOp_107_out) begin
				global_state <= 32'd1;
			end
			if (andOp_116_out) begin
				global_state <= 32'd1;
			end
			if (andOp_128_out) begin
				global_state <= 32'd4;
			end
			if (andOp_219_out) begin
				global_state <= 32'd1;
			end
			if (andOp_220_out) begin
				global_state <= 32'd3;
			end
			if (andOp_221_out) begin
				global_state <= 32'd4;
			end
			if (andOp_222_out) begin
				global_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			icmp_tmp_6 <= 0;
		end else begin
			if (andOp_242_out) begin
				icmp_tmp_6 <= cmp_out_icmp_17;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			phi_tmp_1 <= 0;
		end else begin
			if (andOp_239_out) begin
				phi_tmp_1 <= phi_out_phi_7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (1'd1) begin
				state_0_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_107_out) begin
				state_1_entry_BB_reg <= 32'd9;
			end
			if (andOp_116_out) begin
				state_1_entry_BB_reg <= 32'd3;
			end
			if (andOp_219_out) begin
				state_1_entry_BB_reg <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_107_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_116_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_219_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_228_out) begin
				state_1_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_107_out) begin
				state_1_last_BB_reg <= 32'd9;
			end
			if (andOp_116_out) begin
				state_1_last_BB_reg <= 32'd4;
			end
			if (andOp_219_out) begin
				state_1_last_BB_reg <= bb_0_predecessor_in_state_0_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_107_out) begin
				state_1_last_state <= 32'd1;
			end
			if (andOp_116_out) begin
				state_1_last_state <= 32'd4;
			end
			if (andOp_219_out) begin
				state_1_last_state <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_105_out) begin
				state_2_entry_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_105_out) begin
				state_2_is_active <= 1'd1;
			end
			if (andOp_230_out) begin
				state_2_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_105_out) begin
				state_2_last_BB_reg <= 32'd9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_105_out) begin
				state_2_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_220_out) begin
				state_3_entry_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_220_out) begin
				state_3_is_active <= 1'd1;
			end
			if (andOp_232_out) begin
				state_3_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_220_out) begin
				state_3_last_BB_reg <= bb_10_predecessor_in_state_2_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_state <= 0;
		end else begin
			if (andOp_220_out) begin
				state_3_last_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_128_out) begin
				state_4_entry_BB_reg <= 32'd6;
			end
			if (andOp_221_out) begin
				state_4_entry_BB_reg <= 32'd4;
			end
			if (andOp_222_out) begin
				state_4_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_128_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_221_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_222_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_238_out) begin
				state_4_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_128_out) begin
				state_4_last_BB_reg <= 32'd6;
			end
			if (andOp_221_out) begin
				state_4_last_BB_reg <= bb_4_predecessor_in_state_3_out_data;
			end
			if (andOp_222_out) begin
				state_4_last_BB_reg <= bb_2_predecessor_in_state_4_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_state <= 0;
		end else begin
			if (andOp_128_out) begin
				state_4_last_state <= 32'd4;
			end
			if (andOp_221_out) begin
				state_4_last_state <= 32'd3;
			end
			if (andOp_222_out) begin
				state_4_last_state <= 32'd4;
			end
		end
	end

endmodule

