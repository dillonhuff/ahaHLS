module channel_reduce_4(input [0:0] clk, input [0:0] rst, output [0:0] valid, output [31:0] out_in_data, output [0:0] out_read_valid, output [0:0] out_rst, output [0:0] out_write_valid, input [31:0] out_out_data, input [0:0] out_read_ready, input [0:0] out_write_ready, output [31:0] in_in_data, output [0:0] in_read_valid, output [0:0] in_rst, output [0:0] in_write_valid, input [31:0] in_out_data, input [0:0] in_read_ready, input [0:0] in_write_ready);

	reg [0:0] valid_reg;
	reg [31:0] out_in_data_reg;
	reg [0:0] out_read_valid_reg;
	reg [0:0] out_rst_reg;
	reg [0:0] out_write_valid_reg;
	reg [31:0] in_in_data_reg;
	reg [0:0] in_read_valid_reg;
	reg [0:0] in_rst_reg;
	reg [0:0] in_write_valid_reg;

	assign valid = valid_reg;
	assign out_in_data = out_in_data_reg;
	assign out_read_valid = out_read_valid_reg;
	assign out_rst = out_rst_reg;
	assign out_write_valid = out_write_valid_reg;
	assign in_in_data = in_in_data_reg;
	assign in_read_valid = in_read_valid_reg;
	assign in_rst = in_rst_reg;
	assign in_write_valid = in_write_valid_reg;

	// Start debug wires and ports

	initial begin
	end





	// End debug wires and ports

	// Start Functional Units
	add call_0();

	reg [31:0] raddr_ram_0_reg;
	reg [31:0] waddr_ram_0_reg;
	reg [31:0] wdata_ram_0_reg;
	reg [0:0] wen_ram_0_reg;
	wire [31:0] rdata_ram_0;
	register #(.WIDTH(32)) ram_0(.clk(clk), .raddr(raddr_ram_0_reg), .rdata(rdata_ram_0), .rst(rst), .waddr(waddr_ram_0_reg), .wdata(wdata_ram_0_reg), .wen(wen_ram_0_reg));

	br_dummy br_unit();

	add call_18();

	reg [63:0] phi_in_phi_6;
	reg [31:0] phi_last_block_phi_6;
	reg [63:0] phi_s_phi_6;
	wire [31:0] phi_out_phi_6;
	phi #(.NB_PAIR(2), .WIDTH(32)) phi_6(.in(phi_in_phi_6), .last_block(phi_last_block_phi_6), .out(phi_out_phi_6), .s(phi_s_phi_6));

	reg [31:0] add_in0_add_12;
	reg [31:0] add_in1_add_12;
	wire [31:0] add_out_add_12;
	add #(.WIDTH(32)) add_add_12(.in0(add_in0_add_12), .in1(add_in1_add_12), .out(add_out_add_12));

	reg [31:0] add_in0_add_14;
	reg [31:0] add_in1_add_14;
	wire [31:0] add_out_add_14;
	add #(.WIDTH(32)) add_add_14(.in0(add_in0_add_14), .in1(add_in1_add_14), .out(add_out_add_14));

	reg [31:0] cmp_in0_icmp_15;
	reg [31:0] cmp_in1_icmp_15;
	wire [0:0] cmp_out_icmp_15;
	eq #(.WIDTH(32)) icmp_15(.in0(cmp_in0_icmp_15), .in1(cmp_in1_icmp_15), .out(cmp_out_icmp_15));

	add alloca_2();

	add bitcast_3();

	reg [31:0] data_in_0_1_in_data;
	wire [31:0] data_in_0_1_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_1(.in_data(data_in_0_1_in_data), .out_data(data_in_0_1_out_data));

	reg [31:0] data_in_0_3_in_data;
	wire [31:0] data_in_0_3_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_3(.in_data(data_in_0_3_in_data), .out_data(data_in_0_3_out_data));

	reg [31:0] data_in_0_5_in_data;
	wire [31:0] data_in_0_5_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_5(.in_data(data_in_0_5_in_data), .out_data(data_in_0_5_out_data));

	reg [31:0] data_in_0_7_in_data;
	wire [31:0] data_in_0_7_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_7(.in_data(data_in_0_7_in_data), .out_data(data_in_0_7_out_data));

	reg [0:0] data_in_0_9_in_data;
	wire [0:0] data_in_0_9_out_data;
	hls_wire #(.WIDTH(1)) data_in_0_9(.in_data(data_in_0_9_in_data), .out_data(data_in_0_9_out_data));

	reg [0:0] data_in_0_11_in_data;
	wire [0:0] data_in_0_11_out_data;
	hls_wire #(.WIDTH(1)) data_in_0_11(.in_data(data_in_0_11_in_data), .out_data(data_in_0_11_out_data));

	reg [31:0] data_in_0_13_in_data;
	wire [31:0] data_in_0_13_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_13(.in_data(data_in_0_13_in_data), .out_data(data_in_0_13_out_data));

	reg [0:0] data_in_0_15_in_data;
	wire [0:0] data_in_0_15_out_data;
	hls_wire #(.WIDTH(1)) data_in_0_15(.in_data(data_in_0_15_in_data), .out_data(data_in_0_15_out_data));

	reg [31:0] data_in_0_17_in_data;
	wire [31:0] data_in_0_17_out_data;
	hls_wire #(.WIDTH(32)) data_in_0_17(.in_data(data_in_0_17_in_data), .out_data(data_in_0_17_out_data));

	reg [31:0] data_in_1_19_in_data;
	wire [31:0] data_in_1_19_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_19(.in_data(data_in_1_19_in_data), .out_data(data_in_1_19_out_data));

	reg [31:0] data_in_1_21_in_data;
	wire [31:0] data_in_1_21_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_21(.in_data(data_in_1_21_in_data), .out_data(data_in_1_21_out_data));

	reg [31:0] data_in_1_23_in_data;
	wire [31:0] data_in_1_23_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_23(.in_data(data_in_1_23_in_data), .out_data(data_in_1_23_out_data));

	reg [31:0] data_in_1_25_in_data;
	wire [31:0] data_in_1_25_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_25(.in_data(data_in_1_25_in_data), .out_data(data_in_1_25_out_data));

	reg [0:0] data_in_1_27_in_data;
	wire [0:0] data_in_1_27_out_data;
	hls_wire #(.WIDTH(1)) data_in_1_27(.in_data(data_in_1_27_in_data), .out_data(data_in_1_27_out_data));

	reg [0:0] data_in_1_29_in_data;
	wire [0:0] data_in_1_29_out_data;
	hls_wire #(.WIDTH(1)) data_in_1_29(.in_data(data_in_1_29_in_data), .out_data(data_in_1_29_out_data));

	reg [31:0] data_in_1_31_in_data;
	wire [31:0] data_in_1_31_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_31(.in_data(data_in_1_31_in_data), .out_data(data_in_1_31_out_data));

	reg [0:0] data_in_1_33_in_data;
	wire [0:0] data_in_1_33_out_data;
	hls_wire #(.WIDTH(1)) data_in_1_33(.in_data(data_in_1_33_in_data), .out_data(data_in_1_33_out_data));

	reg [31:0] data_in_1_35_in_data;
	wire [31:0] data_in_1_35_out_data;
	hls_wire #(.WIDTH(32)) data_in_1_35(.in_data(data_in_1_35_in_data), .out_data(data_in_1_35_out_data));

	reg [31:0] data_in_2_37_in_data;
	wire [31:0] data_in_2_37_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_37(.in_data(data_in_2_37_in_data), .out_data(data_in_2_37_out_data));

	reg [31:0] data_in_2_39_in_data;
	wire [31:0] data_in_2_39_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_39(.in_data(data_in_2_39_in_data), .out_data(data_in_2_39_out_data));

	reg [31:0] data_in_2_41_in_data;
	wire [31:0] data_in_2_41_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_41(.in_data(data_in_2_41_in_data), .out_data(data_in_2_41_out_data));

	reg [31:0] data_in_2_43_in_data;
	wire [31:0] data_in_2_43_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_43(.in_data(data_in_2_43_in_data), .out_data(data_in_2_43_out_data));

	reg [0:0] data_in_2_45_in_data;
	wire [0:0] data_in_2_45_out_data;
	hls_wire #(.WIDTH(1)) data_in_2_45(.in_data(data_in_2_45_in_data), .out_data(data_in_2_45_out_data));

	reg [0:0] data_in_2_47_in_data;
	wire [0:0] data_in_2_47_out_data;
	hls_wire #(.WIDTH(1)) data_in_2_47(.in_data(data_in_2_47_in_data), .out_data(data_in_2_47_out_data));

	reg [31:0] data_in_2_49_in_data;
	wire [31:0] data_in_2_49_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_49(.in_data(data_in_2_49_in_data), .out_data(data_in_2_49_out_data));

	reg [0:0] data_in_2_51_in_data;
	wire [0:0] data_in_2_51_out_data;
	hls_wire #(.WIDTH(1)) data_in_2_51(.in_data(data_in_2_51_in_data), .out_data(data_in_2_51_out_data));

	reg [31:0] data_in_2_53_in_data;
	wire [31:0] data_in_2_53_out_data;
	hls_wire #(.WIDTH(32)) data_in_2_53(.in_data(data_in_2_53_in_data), .out_data(data_in_2_53_out_data));

	reg [31:0] data_in_3_55_in_data;
	wire [31:0] data_in_3_55_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_55(.in_data(data_in_3_55_in_data), .out_data(data_in_3_55_out_data));

	reg [31:0] data_in_3_57_in_data;
	wire [31:0] data_in_3_57_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_57(.in_data(data_in_3_57_in_data), .out_data(data_in_3_57_out_data));

	reg [31:0] data_in_3_59_in_data;
	wire [31:0] data_in_3_59_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_59(.in_data(data_in_3_59_in_data), .out_data(data_in_3_59_out_data));

	reg [31:0] data_in_3_61_in_data;
	wire [31:0] data_in_3_61_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_61(.in_data(data_in_3_61_in_data), .out_data(data_in_3_61_out_data));

	reg [0:0] data_in_3_63_in_data;
	wire [0:0] data_in_3_63_out_data;
	hls_wire #(.WIDTH(1)) data_in_3_63(.in_data(data_in_3_63_in_data), .out_data(data_in_3_63_out_data));

	reg [0:0] data_in_3_65_in_data;
	wire [0:0] data_in_3_65_out_data;
	hls_wire #(.WIDTH(1)) data_in_3_65(.in_data(data_in_3_65_in_data), .out_data(data_in_3_65_out_data));

	reg [31:0] data_in_3_67_in_data;
	wire [31:0] data_in_3_67_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_67(.in_data(data_in_3_67_in_data), .out_data(data_in_3_67_out_data));

	reg [0:0] data_in_3_69_in_data;
	wire [0:0] data_in_3_69_out_data;
	hls_wire #(.WIDTH(1)) data_in_3_69(.in_data(data_in_3_69_in_data), .out_data(data_in_3_69_out_data));

	reg [31:0] data_in_3_71_in_data;
	wire [31:0] data_in_3_71_out_data;
	hls_wire #(.WIDTH(32)) data_in_3_71(.in_data(data_in_3_71_in_data), .out_data(data_in_3_71_out_data));

	reg [31:0] data_in_4_73_in_data;
	wire [31:0] data_in_4_73_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_73(.in_data(data_in_4_73_in_data), .out_data(data_in_4_73_out_data));

	reg [31:0] data_in_4_75_in_data;
	wire [31:0] data_in_4_75_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_75(.in_data(data_in_4_75_in_data), .out_data(data_in_4_75_out_data));

	reg [31:0] data_in_4_77_in_data;
	wire [31:0] data_in_4_77_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_77(.in_data(data_in_4_77_in_data), .out_data(data_in_4_77_out_data));

	reg [31:0] data_in_4_79_in_data;
	wire [31:0] data_in_4_79_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_79(.in_data(data_in_4_79_in_data), .out_data(data_in_4_79_out_data));

	reg [0:0] data_in_4_81_in_data;
	wire [0:0] data_in_4_81_out_data;
	hls_wire #(.WIDTH(1)) data_in_4_81(.in_data(data_in_4_81_in_data), .out_data(data_in_4_81_out_data));

	reg [0:0] data_in_4_83_in_data;
	wire [0:0] data_in_4_83_out_data;
	hls_wire #(.WIDTH(1)) data_in_4_83(.in_data(data_in_4_83_in_data), .out_data(data_in_4_83_out_data));

	reg [31:0] data_in_4_85_in_data;
	wire [31:0] data_in_4_85_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_85(.in_data(data_in_4_85_in_data), .out_data(data_in_4_85_out_data));

	reg [0:0] data_in_4_87_in_data;
	wire [0:0] data_in_4_87_out_data;
	hls_wire #(.WIDTH(1)) data_in_4_87(.in_data(data_in_4_87_in_data), .out_data(data_in_4_87_out_data));

	reg [31:0] data_in_4_89_in_data;
	wire [31:0] data_in_4_89_out_data;
	hls_wire #(.WIDTH(32)) data_in_4_89(.in_data(data_in_4_89_in_data), .out_data(data_in_4_89_out_data));

	reg [0:0] bb_0_active_in_state_0_in_data;
	wire [0:0] bb_0_active_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_0(.in_data(bb_0_active_in_state_0_in_data), .out_data(bb_0_active_in_state_0_out_data));

	reg [31:0] bb_0_predecessor_in_state_0_in_data;
	wire [31:0] bb_0_predecessor_in_state_0_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_0(.in_data(bb_0_predecessor_in_state_0_in_data), .out_data(bb_0_predecessor_in_state_0_out_data));

	reg [0:0] bb_3_active_in_state_1_in_data;
	wire [0:0] bb_3_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_3_active_in_state_1(.in_data(bb_3_active_in_state_1_in_data), .out_data(bb_3_active_in_state_1_out_data));

	reg [31:0] bb_3_predecessor_in_state_1_in_data;
	wire [31:0] bb_3_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_3_predecessor_in_state_1(.in_data(bb_3_predecessor_in_state_1_in_data), .out_data(bb_3_predecessor_in_state_1_out_data));

	reg [0:0] bb_8_active_in_state_1_in_data;
	wire [0:0] bb_8_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_8_active_in_state_1(.in_data(bb_8_active_in_state_1_in_data), .out_data(bb_8_active_in_state_1_out_data));

	reg [31:0] bb_8_predecessor_in_state_1_in_data;
	wire [31:0] bb_8_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_8_predecessor_in_state_1(.in_data(bb_8_predecessor_in_state_1_in_data), .out_data(bb_8_predecessor_in_state_1_out_data));

	reg [0:0] bb_9_active_in_state_1_in_data;
	wire [0:0] bb_9_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_9_active_in_state_1(.in_data(bb_9_active_in_state_1_in_data), .out_data(bb_9_active_in_state_1_out_data));

	reg [31:0] bb_9_predecessor_in_state_1_in_data;
	wire [31:0] bb_9_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_9_predecessor_in_state_1(.in_data(bb_9_predecessor_in_state_1_in_data), .out_data(bb_9_predecessor_in_state_1_out_data));

	reg [0:0] bb_0_active_in_state_1_in_data;
	wire [0:0] bb_0_active_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) bb_0_active_in_state_1(.in_data(bb_0_active_in_state_1_in_data), .out_data(bb_0_active_in_state_1_out_data));

	reg [31:0] bb_0_predecessor_in_state_1_in_data;
	wire [31:0] bb_0_predecessor_in_state_1_out_data;
	hls_wire #(.WIDTH(32)) bb_0_predecessor_in_state_1(.in_data(bb_0_predecessor_in_state_1_in_data), .out_data(bb_0_predecessor_in_state_1_out_data));

	reg [0:0] bb_10_active_in_state_2_in_data;
	wire [0:0] bb_10_active_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_2(.in_data(bb_10_active_in_state_2_in_data), .out_data(bb_10_active_in_state_2_out_data));

	reg [31:0] bb_10_predecessor_in_state_2_in_data;
	wire [31:0] bb_10_predecessor_in_state_2_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_2(.in_data(bb_10_predecessor_in_state_2_in_data), .out_data(bb_10_predecessor_in_state_2_out_data));

	reg [0:0] bb_10_active_in_state_3_in_data;
	wire [0:0] bb_10_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_10_active_in_state_3(.in_data(bb_10_active_in_state_3_in_data), .out_data(bb_10_active_in_state_3_out_data));

	reg [31:0] bb_10_predecessor_in_state_3_in_data;
	wire [31:0] bb_10_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_10_predecessor_in_state_3(.in_data(bb_10_predecessor_in_state_3_in_data), .out_data(bb_10_predecessor_in_state_3_out_data));

	reg [0:0] bb_4_active_in_state_3_in_data;
	wire [0:0] bb_4_active_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_3(.in_data(bb_4_active_in_state_3_in_data), .out_data(bb_4_active_in_state_3_out_data));

	reg [31:0] bb_4_predecessor_in_state_3_in_data;
	wire [31:0] bb_4_predecessor_in_state_3_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_3(.in_data(bb_4_predecessor_in_state_3_in_data), .out_data(bb_4_predecessor_in_state_3_out_data));

	reg [0:0] bb_1_active_in_state_4_in_data;
	wire [0:0] bb_1_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_1_active_in_state_4(.in_data(bb_1_active_in_state_4_in_data), .out_data(bb_1_active_in_state_4_out_data));

	reg [31:0] bb_1_predecessor_in_state_4_in_data;
	wire [31:0] bb_1_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_1_predecessor_in_state_4(.in_data(bb_1_predecessor_in_state_4_in_data), .out_data(bb_1_predecessor_in_state_4_out_data));

	reg [0:0] bb_5_active_in_state_4_in_data;
	wire [0:0] bb_5_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_5_active_in_state_4(.in_data(bb_5_active_in_state_4_in_data), .out_data(bb_5_active_in_state_4_out_data));

	reg [31:0] bb_5_predecessor_in_state_4_in_data;
	wire [31:0] bb_5_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_5_predecessor_in_state_4(.in_data(bb_5_predecessor_in_state_4_in_data), .out_data(bb_5_predecessor_in_state_4_out_data));

	reg [0:0] bb_6_active_in_state_4_in_data;
	wire [0:0] bb_6_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_6_active_in_state_4(.in_data(bb_6_active_in_state_4_in_data), .out_data(bb_6_active_in_state_4_out_data));

	reg [31:0] bb_6_predecessor_in_state_4_in_data;
	wire [31:0] bb_6_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_6_predecessor_in_state_4(.in_data(bb_6_predecessor_in_state_4_in_data), .out_data(bb_6_predecessor_in_state_4_out_data));

	reg [0:0] bb_7_active_in_state_4_in_data;
	wire [0:0] bb_7_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_7_active_in_state_4(.in_data(bb_7_active_in_state_4_in_data), .out_data(bb_7_active_in_state_4_out_data));

	reg [31:0] bb_7_predecessor_in_state_4_in_data;
	wire [31:0] bb_7_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_7_predecessor_in_state_4(.in_data(bb_7_predecessor_in_state_4_in_data), .out_data(bb_7_predecessor_in_state_4_out_data));

	reg [0:0] bb_4_active_in_state_4_in_data;
	wire [0:0] bb_4_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_4_active_in_state_4(.in_data(bb_4_active_in_state_4_in_data), .out_data(bb_4_active_in_state_4_out_data));

	reg [31:0] bb_4_predecessor_in_state_4_in_data;
	wire [31:0] bb_4_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_4_predecessor_in_state_4(.in_data(bb_4_predecessor_in_state_4_in_data), .out_data(bb_4_predecessor_in_state_4_out_data));

	reg [0:0] bb_2_active_in_state_4_in_data;
	wire [0:0] bb_2_active_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) bb_2_active_in_state_4(.in_data(bb_2_active_in_state_4_in_data), .out_data(bb_2_active_in_state_4_out_data));

	reg [31:0] bb_2_predecessor_in_state_4_in_data;
	wire [31:0] bb_2_predecessor_in_state_4_out_data;
	hls_wire #(.WIDTH(32)) bb_2_predecessor_in_state_4(.in_data(bb_2_predecessor_in_state_4_in_data), .out_data(bb_2_predecessor_in_state_4_out_data));

	reg [0:0] andOp_90_in0;
	reg [0:0] andOp_90_in1;
	wire [0:0] andOp_90_out;
	andOp #(.WIDTH(1)) andOp_90(.in0(andOp_90_in0), .in1(andOp_90_in1), .out(andOp_90_out));

	reg [0:0] andOp_91_in0;
	reg [0:0] andOp_91_in1;
	wire [0:0] andOp_91_out;
	andOp #(.WIDTH(1)) andOp_91(.in0(andOp_91_in0), .in1(andOp_91_in1), .out(andOp_91_out));

	reg [0:0] br_0_happened_in_state_0_in_data;
	wire [0:0] br_0_happened_in_state_0_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_0(.in_data(br_0_happened_in_state_0_in_data), .out_data(br_0_happened_in_state_0_out_data));

	reg [0:0] notOp_92_in0;
	wire [0:0] notOp_92_out;
	notOp #(.WIDTH(1)) notOp_92(.in(notOp_92_in0), .out(notOp_92_out));

	reg [0:0] andOp_93_in0;
	reg [0:0] andOp_93_in1;
	wire [0:0] andOp_93_out;
	andOp #(.WIDTH(1)) andOp_93(.in0(andOp_93_in0), .in1(andOp_93_in1), .out(andOp_93_out));

	reg [0:0] andOp_94_in0;
	reg [0:0] andOp_94_in1;
	wire [0:0] andOp_94_out;
	andOp #(.WIDTH(1)) andOp_94(.in0(andOp_94_in0), .in1(andOp_94_in1), .out(andOp_94_out));

	reg [0:0] br_3_happened_in_state_1_in_data;
	wire [0:0] br_3_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_3_happened_in_state_1(.in_data(br_3_happened_in_state_1_in_data), .out_data(br_3_happened_in_state_1_out_data));

	reg [0:0] notOp_95_in0;
	wire [0:0] notOp_95_out;
	notOp #(.WIDTH(1)) notOp_95(.in(notOp_95_in0), .out(notOp_95_out));

	reg [0:0] andOp_96_in0;
	reg [0:0] andOp_96_in1;
	wire [0:0] andOp_96_out;
	andOp #(.WIDTH(1)) andOp_96(.in0(andOp_96_in0), .in1(andOp_96_in1), .out(andOp_96_out));

	reg [0:0] andOp_97_in0;
	reg [0:0] andOp_97_in1;
	wire [0:0] andOp_97_out;
	andOp #(.WIDTH(1)) andOp_97(.in0(andOp_97_in0), .in1(andOp_97_in1), .out(andOp_97_out));

	reg [0:0] br_8_happened_in_state_1_in_data;
	wire [0:0] br_8_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_8_happened_in_state_1(.in_data(br_8_happened_in_state_1_in_data), .out_data(br_8_happened_in_state_1_out_data));

	reg [0:0] notOp_98_in0;
	wire [0:0] notOp_98_out;
	notOp #(.WIDTH(1)) notOp_98(.in(notOp_98_in0), .out(notOp_98_out));

	reg [0:0] andOp_99_in0;
	reg [0:0] andOp_99_in1;
	wire [0:0] andOp_99_out;
	andOp #(.WIDTH(1)) andOp_99(.in0(andOp_99_in0), .in1(andOp_99_in1), .out(andOp_99_out));

	reg [0:0] andOp_100_in0;
	reg [0:0] andOp_100_in1;
	wire [0:0] andOp_100_out;
	andOp #(.WIDTH(1)) andOp_100(.in0(andOp_100_in0), .in1(andOp_100_in1), .out(andOp_100_out));

	reg [0:0] br_9_happened_in_state_1_in_data;
	wire [0:0] br_9_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_9_happened_in_state_1(.in_data(br_9_happened_in_state_1_in_data), .out_data(br_9_happened_in_state_1_out_data));

	reg [0:0] notOp_101_in0;
	wire [0:0] notOp_101_out;
	notOp #(.WIDTH(1)) notOp_101(.in(notOp_101_in0), .out(notOp_101_out));

	reg [0:0] andOp_102_in0;
	reg [0:0] andOp_102_in1;
	wire [0:0] andOp_102_out;
	andOp #(.WIDTH(1)) andOp_102(.in0(andOp_102_in0), .in1(andOp_102_in1), .out(andOp_102_out));

	reg [0:0] notOp_103_in0;
	wire [0:0] notOp_103_out;
	notOp #(.WIDTH(1)) notOp_103(.in(notOp_103_in0), .out(notOp_103_out));

	reg [0:0] andOp_104_in0;
	reg [0:0] andOp_104_in1;
	wire [0:0] andOp_104_out;
	andOp #(.WIDTH(1)) andOp_104(.in0(andOp_104_in0), .in1(andOp_104_in1), .out(andOp_104_out));

	reg [0:0] andOp_105_in0;
	reg [0:0] andOp_105_in1;
	wire [0:0] andOp_105_out;
	andOp #(.WIDTH(1)) andOp_105(.in0(andOp_105_in0), .in1(andOp_105_in1), .out(andOp_105_out));

	reg [0:0] andOp_106_in0;
	reg [0:0] andOp_106_in1;
	wire [0:0] andOp_106_out;
	andOp #(.WIDTH(1)) andOp_106(.in0(andOp_106_in0), .in1(andOp_106_in1), .out(andOp_106_out));

	reg [0:0] br_0_happened_in_state_1_in_data;
	wire [0:0] br_0_happened_in_state_1_out_data;
	hls_wire #(.WIDTH(1)) br_0_happened_in_state_1(.in_data(br_0_happened_in_state_1_in_data), .out_data(br_0_happened_in_state_1_out_data));

	reg [0:0] notOp_107_in0;
	wire [0:0] notOp_107_out;
	notOp #(.WIDTH(1)) notOp_107(.in(notOp_107_in0), .out(notOp_107_out));

	reg [0:0] andOp_108_in0;
	reg [0:0] andOp_108_in1;
	wire [0:0] andOp_108_out;
	andOp #(.WIDTH(1)) andOp_108(.in0(andOp_108_in0), .in1(andOp_108_in1), .out(andOp_108_out));

	reg [0:0] andOp_109_in0;
	reg [0:0] andOp_109_in1;
	wire [0:0] andOp_109_out;
	andOp #(.WIDTH(1)) andOp_109(.in0(andOp_109_in0), .in1(andOp_109_in1), .out(andOp_109_out));

	reg [0:0] br_10_happened_in_state_2_in_data;
	wire [0:0] br_10_happened_in_state_2_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_2(.in_data(br_10_happened_in_state_2_in_data), .out_data(br_10_happened_in_state_2_out_data));

	reg [0:0] notOp_110_in0;
	wire [0:0] notOp_110_out;
	notOp #(.WIDTH(1)) notOp_110(.in(notOp_110_in0), .out(notOp_110_out));

	reg [0:0] andOp_111_in0;
	reg [0:0] andOp_111_in1;
	wire [0:0] andOp_111_out;
	andOp #(.WIDTH(1)) andOp_111(.in0(andOp_111_in0), .in1(andOp_111_in1), .out(andOp_111_out));

	reg [0:0] andOp_112_in0;
	reg [0:0] andOp_112_in1;
	wire [0:0] andOp_112_out;
	andOp #(.WIDTH(1)) andOp_112(.in0(andOp_112_in0), .in1(andOp_112_in1), .out(andOp_112_out));

	reg [0:0] br_10_happened_in_state_3_in_data;
	wire [0:0] br_10_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_10_happened_in_state_3(.in_data(br_10_happened_in_state_3_in_data), .out_data(br_10_happened_in_state_3_out_data));

	reg [0:0] notOp_113_in0;
	wire [0:0] notOp_113_out;
	notOp #(.WIDTH(1)) notOp_113(.in(notOp_113_in0), .out(notOp_113_out));

	reg [0:0] andOp_114_in0;
	reg [0:0] andOp_114_in1;
	wire [0:0] andOp_114_out;
	andOp #(.WIDTH(1)) andOp_114(.in0(andOp_114_in0), .in1(andOp_114_in1), .out(andOp_114_out));

	reg [0:0] andOp_115_in0;
	reg [0:0] andOp_115_in1;
	wire [0:0] andOp_115_out;
	andOp #(.WIDTH(1)) andOp_115(.in0(andOp_115_in0), .in1(andOp_115_in1), .out(andOp_115_out));

	reg [0:0] br_4_happened_in_state_3_in_data;
	wire [0:0] br_4_happened_in_state_3_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_3(.in_data(br_4_happened_in_state_3_in_data), .out_data(br_4_happened_in_state_3_out_data));

	reg [0:0] notOp_116_in0;
	wire [0:0] notOp_116_out;
	notOp #(.WIDTH(1)) notOp_116(.in(notOp_116_in0), .out(notOp_116_out));

	reg [0:0] andOp_117_in0;
	reg [0:0] andOp_117_in1;
	wire [0:0] andOp_117_out;
	andOp #(.WIDTH(1)) andOp_117(.in0(andOp_117_in0), .in1(andOp_117_in1), .out(andOp_117_out));

	reg [0:0] notOp_118_in0;
	wire [0:0] notOp_118_out;
	notOp #(.WIDTH(1)) notOp_118(.in(notOp_118_in0), .out(notOp_118_out));

	reg [0:0] andOp_119_in0;
	reg [0:0] andOp_119_in1;
	wire [0:0] andOp_119_out;
	andOp #(.WIDTH(1)) andOp_119(.in0(andOp_119_in0), .in1(andOp_119_in1), .out(andOp_119_out));

	reg [0:0] andOp_120_in0;
	reg [0:0] andOp_120_in1;
	wire [0:0] andOp_120_out;
	andOp #(.WIDTH(1)) andOp_120(.in0(andOp_120_in0), .in1(andOp_120_in1), .out(andOp_120_out));

	reg [0:0] andOp_121_in0;
	reg [0:0] andOp_121_in1;
	wire [0:0] andOp_121_out;
	andOp #(.WIDTH(1)) andOp_121(.in0(andOp_121_in0), .in1(andOp_121_in1), .out(andOp_121_out));

	reg [0:0] br_1_happened_in_state_4_in_data;
	wire [0:0] br_1_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_1_happened_in_state_4(.in_data(br_1_happened_in_state_4_in_data), .out_data(br_1_happened_in_state_4_out_data));

	reg [0:0] notOp_122_in0;
	wire [0:0] notOp_122_out;
	notOp #(.WIDTH(1)) notOp_122(.in(notOp_122_in0), .out(notOp_122_out));

	reg [0:0] andOp_123_in0;
	reg [0:0] andOp_123_in1;
	wire [0:0] andOp_123_out;
	andOp #(.WIDTH(1)) andOp_123(.in0(andOp_123_in0), .in1(andOp_123_in1), .out(andOp_123_out));

	reg [0:0] andOp_124_in0;
	reg [0:0] andOp_124_in1;
	wire [0:0] andOp_124_out;
	andOp #(.WIDTH(1)) andOp_124(.in0(andOp_124_in0), .in1(andOp_124_in1), .out(andOp_124_out));

	reg [0:0] br_5_happened_in_state_4_in_data;
	wire [0:0] br_5_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_5_happened_in_state_4(.in_data(br_5_happened_in_state_4_in_data), .out_data(br_5_happened_in_state_4_out_data));

	reg [0:0] notOp_125_in0;
	wire [0:0] notOp_125_out;
	notOp #(.WIDTH(1)) notOp_125(.in(notOp_125_in0), .out(notOp_125_out));

	reg [0:0] andOp_126_in0;
	reg [0:0] andOp_126_in1;
	wire [0:0] andOp_126_out;
	andOp #(.WIDTH(1)) andOp_126(.in0(andOp_126_in0), .in1(andOp_126_in1), .out(andOp_126_out));

	reg [0:0] andOp_127_in0;
	reg [0:0] andOp_127_in1;
	wire [0:0] andOp_127_out;
	andOp #(.WIDTH(1)) andOp_127(.in0(andOp_127_in0), .in1(andOp_127_in1), .out(andOp_127_out));

	reg [0:0] br_6_happened_in_state_4_in_data;
	wire [0:0] br_6_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_6_happened_in_state_4(.in_data(br_6_happened_in_state_4_in_data), .out_data(br_6_happened_in_state_4_out_data));

	reg [0:0] notOp_128_in0;
	wire [0:0] notOp_128_out;
	notOp #(.WIDTH(1)) notOp_128(.in(notOp_128_in0), .out(notOp_128_out));

	reg [0:0] andOp_129_in0;
	reg [0:0] andOp_129_in1;
	wire [0:0] andOp_129_out;
	andOp #(.WIDTH(1)) andOp_129(.in0(andOp_129_in0), .in1(andOp_129_in1), .out(andOp_129_out));

	reg [0:0] notOp_130_in0;
	wire [0:0] notOp_130_out;
	notOp #(.WIDTH(1)) notOp_130(.in(notOp_130_in0), .out(notOp_130_out));

	reg [0:0] andOp_131_in0;
	reg [0:0] andOp_131_in1;
	wire [0:0] andOp_131_out;
	andOp #(.WIDTH(1)) andOp_131(.in0(andOp_131_in0), .in1(andOp_131_in1), .out(andOp_131_out));

	reg [0:0] andOp_132_in0;
	reg [0:0] andOp_132_in1;
	wire [0:0] andOp_132_out;
	andOp #(.WIDTH(1)) andOp_132(.in0(andOp_132_in0), .in1(andOp_132_in1), .out(andOp_132_out));

	reg [0:0] andOp_133_in0;
	reg [0:0] andOp_133_in1;
	wire [0:0] andOp_133_out;
	andOp #(.WIDTH(1)) andOp_133(.in0(andOp_133_in0), .in1(andOp_133_in1), .out(andOp_133_out));

	reg [0:0] br_7_happened_in_state_4_in_data;
	wire [0:0] br_7_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_7_happened_in_state_4(.in_data(br_7_happened_in_state_4_in_data), .out_data(br_7_happened_in_state_4_out_data));

	reg [0:0] notOp_134_in0;
	wire [0:0] notOp_134_out;
	notOp #(.WIDTH(1)) notOp_134(.in(notOp_134_in0), .out(notOp_134_out));

	reg [0:0] andOp_135_in0;
	reg [0:0] andOp_135_in1;
	wire [0:0] andOp_135_out;
	andOp #(.WIDTH(1)) andOp_135(.in0(andOp_135_in0), .in1(andOp_135_in1), .out(andOp_135_out));

	reg [0:0] andOp_136_in0;
	reg [0:0] andOp_136_in1;
	wire [0:0] andOp_136_out;
	andOp #(.WIDTH(1)) andOp_136(.in0(andOp_136_in0), .in1(andOp_136_in1), .out(andOp_136_out));

	reg [0:0] br_4_happened_in_state_4_in_data;
	wire [0:0] br_4_happened_in_state_4_out_data;
	hls_wire #(.WIDTH(1)) br_4_happened_in_state_4(.in_data(br_4_happened_in_state_4_in_data), .out_data(br_4_happened_in_state_4_out_data));

	reg [0:0] notOp_137_in0;
	wire [0:0] notOp_137_out;
	notOp #(.WIDTH(1)) notOp_137(.in(notOp_137_in0), .out(notOp_137_out));

	reg [0:0] andOp_138_in0;
	reg [0:0] andOp_138_in1;
	wire [0:0] andOp_138_out;
	andOp #(.WIDTH(1)) andOp_138(.in0(andOp_138_in0), .in1(andOp_138_in1), .out(andOp_138_out));

	reg [0:0] notOp_139_in0;
	wire [0:0] notOp_139_out;
	notOp #(.WIDTH(1)) notOp_139(.in(notOp_139_in0), .out(notOp_139_out));

	reg [0:0] andOp_140_in0;
	reg [0:0] andOp_140_in1;
	wire [0:0] andOp_140_out;
	andOp #(.WIDTH(1)) andOp_140(.in0(andOp_140_in0), .in1(andOp_140_in1), .out(andOp_140_out));

	reg [31:0] eq_141_in0;
	reg [31:0] eq_141_in1;
	wire [0:0] eq_141_out;
	eq #(.WIDTH(32)) eq_141(.in0(eq_141_in0), .in1(eq_141_in1), .out(eq_141_out));

	reg [31:0] eq_142_in0;
	reg [31:0] eq_142_in1;
	wire [0:0] eq_142_out;
	eq #(.WIDTH(32)) eq_142(.in0(eq_142_in0), .in1(eq_142_in1), .out(eq_142_out));

	reg [0:0] orOp_143_in0;
	reg [0:0] orOp_143_in1;
	wire [0:0] orOp_143_out;
	orOp #(.WIDTH(1)) orOp_143(.in0(orOp_143_in0), .in1(orOp_143_in1), .out(orOp_143_out));

	reg [31:0] eq_144_in0;
	reg [31:0] eq_144_in1;
	wire [0:0] eq_144_out;
	eq #(.WIDTH(32)) eq_144(.in0(eq_144_in0), .in1(eq_144_in1), .out(eq_144_out));

	reg [0:0] orOp_145_in0;
	reg [0:0] orOp_145_in1;
	wire [0:0] orOp_145_out;
	orOp #(.WIDTH(1)) orOp_145(.in0(orOp_145_in0), .in1(orOp_145_in1), .out(orOp_145_out));

	reg [31:0] eq_146_in0;
	reg [31:0] eq_146_in1;
	wire [0:0] eq_146_out;
	eq #(.WIDTH(32)) eq_146(.in0(eq_146_in0), .in1(eq_146_in1), .out(eq_146_out));

	reg [0:0] orOp_147_in0;
	reg [0:0] orOp_147_in1;
	wire [0:0] orOp_147_out;
	orOp #(.WIDTH(1)) orOp_147(.in0(orOp_147_in0), .in1(orOp_147_in1), .out(orOp_147_out));

	reg [31:0] eq_148_in0;
	reg [31:0] eq_148_in1;
	wire [0:0] eq_148_out;
	eq #(.WIDTH(32)) eq_148(.in0(eq_148_in0), .in1(eq_148_in1), .out(eq_148_out));

	reg [31:0] eq_149_in0;
	reg [31:0] eq_149_in1;
	wire [0:0] eq_149_out;
	eq #(.WIDTH(32)) eq_149(.in0(eq_149_in0), .in1(eq_149_in1), .out(eq_149_out));

	reg [31:0] eq_150_in0;
	reg [31:0] eq_150_in1;
	wire [0:0] eq_150_out;
	eq #(.WIDTH(32)) eq_150(.in0(eq_150_in0), .in1(eq_150_in1), .out(eq_150_out));

	reg [31:0] eq_151_in0;
	reg [31:0] eq_151_in1;
	wire [0:0] eq_151_out;
	eq #(.WIDTH(32)) eq_151(.in0(eq_151_in0), .in1(eq_151_in1), .out(eq_151_out));

	reg [0:0] orOp_152_in0;
	reg [0:0] orOp_152_in1;
	wire [0:0] orOp_152_out;
	orOp #(.WIDTH(1)) orOp_152(.in0(orOp_152_in0), .in1(orOp_152_in1), .out(orOp_152_out));

	reg [31:0] eq_153_in0;
	reg [31:0] eq_153_in1;
	wire [0:0] eq_153_out;
	eq #(.WIDTH(32)) eq_153(.in0(eq_153_in0), .in1(eq_153_in1), .out(eq_153_out));

	reg [0:0] orOp_154_in0;
	reg [0:0] orOp_154_in1;
	wire [0:0] orOp_154_out;
	orOp #(.WIDTH(1)) orOp_154(.in0(orOp_154_in0), .in1(orOp_154_in1), .out(orOp_154_out));

	reg [31:0] eq_155_in0;
	reg [31:0] eq_155_in1;
	wire [0:0] eq_155_out;
	eq #(.WIDTH(32)) eq_155(.in0(eq_155_in0), .in1(eq_155_in1), .out(eq_155_out));

	reg [0:0] orOp_156_in0;
	reg [0:0] orOp_156_in1;
	wire [0:0] orOp_156_out;
	orOp #(.WIDTH(1)) orOp_156(.in0(orOp_156_in0), .in1(orOp_156_in1), .out(orOp_156_out));

	reg [31:0] eq_157_in0;
	reg [31:0] eq_157_in1;
	wire [0:0] eq_157_out;
	eq #(.WIDTH(32)) eq_157(.in0(eq_157_in0), .in1(eq_157_in1), .out(eq_157_out));

	reg [0:0] orOp_158_in0;
	reg [0:0] orOp_158_in1;
	wire [0:0] orOp_158_out;
	orOp #(.WIDTH(1)) orOp_158(.in0(orOp_158_in0), .in1(orOp_158_in1), .out(orOp_158_out));

	reg [31:0] eq_159_in0;
	reg [31:0] eq_159_in1;
	wire [0:0] eq_159_out;
	eq #(.WIDTH(32)) eq_159(.in0(eq_159_in0), .in1(eq_159_in1), .out(eq_159_out));

	reg [0:0] orOp_160_in0;
	reg [0:0] orOp_160_in1;
	wire [0:0] orOp_160_out;
	orOp #(.WIDTH(1)) orOp_160(.in0(orOp_160_in0), .in1(orOp_160_in1), .out(orOp_160_out));

	reg [31:0] eq_161_in0;
	reg [31:0] eq_161_in1;
	wire [0:0] eq_161_out;
	eq #(.WIDTH(32)) eq_161(.in0(eq_161_in0), .in1(eq_161_in1), .out(eq_161_out));

	reg [31:0] eq_162_in0;
	reg [31:0] eq_162_in1;
	wire [0:0] eq_162_out;
	eq #(.WIDTH(32)) eq_162(.in0(eq_162_in0), .in1(eq_162_in1), .out(eq_162_out));

	reg [0:0] orOp_163_in0;
	reg [0:0] orOp_163_in1;
	wire [0:0] orOp_163_out;
	orOp #(.WIDTH(1)) orOp_163(.in0(orOp_163_in0), .in1(orOp_163_in1), .out(orOp_163_out));

	reg [31:0] eq_164_in0;
	reg [31:0] eq_164_in1;
	wire [0:0] eq_164_out;
	eq #(.WIDTH(32)) eq_164(.in0(eq_164_in0), .in1(eq_164_in1), .out(eq_164_out));

	reg [31:0] eq_165_in0;
	reg [31:0] eq_165_in1;
	wire [0:0] eq_165_out;
	eq #(.WIDTH(32)) eq_165(.in0(eq_165_in0), .in1(eq_165_in1), .out(eq_165_out));

	reg [0:0] notOp_166_in0;
	wire [0:0] notOp_166_out;
	notOp #(.WIDTH(1)) notOp_166(.in(notOp_166_in0), .out(notOp_166_out));

	reg [0:0] andOp_167_in0;
	reg [0:0] andOp_167_in1;
	wire [0:0] andOp_167_out;
	andOp #(.WIDTH(1)) andOp_167(.in0(andOp_167_in0), .in1(andOp_167_in1), .out(andOp_167_out));

	reg [31:0] eq_168_in0;
	reg [31:0] eq_168_in1;
	wire [0:0] eq_168_out;
	eq #(.WIDTH(32)) eq_168(.in0(eq_168_in0), .in1(eq_168_in1), .out(eq_168_out));

	reg [0:0] notOp_169_in0;
	wire [0:0] notOp_169_out;
	notOp #(.WIDTH(1)) notOp_169(.in(notOp_169_in0), .out(notOp_169_out));

	reg [0:0] andOp_170_in0;
	reg [0:0] andOp_170_in1;
	wire [0:0] andOp_170_out;
	andOp #(.WIDTH(1)) andOp_170(.in0(andOp_170_in0), .in1(andOp_170_in1), .out(andOp_170_out));

	reg [31:0] eq_171_in0;
	reg [31:0] eq_171_in1;
	wire [0:0] eq_171_out;
	eq #(.WIDTH(32)) eq_171(.in0(eq_171_in0), .in1(eq_171_in1), .out(eq_171_out));

	reg [0:0] notOp_172_in0;
	wire [0:0] notOp_172_out;
	notOp #(.WIDTH(1)) notOp_172(.in(notOp_172_in0), .out(notOp_172_out));

	reg [0:0] andOp_173_in0;
	reg [0:0] andOp_173_in1;
	wire [0:0] andOp_173_out;
	andOp #(.WIDTH(1)) andOp_173(.in0(andOp_173_in0), .in1(andOp_173_in1), .out(andOp_173_out));

	reg [31:0] eq_174_in0;
	reg [31:0] eq_174_in1;
	wire [0:0] eq_174_out;
	eq #(.WIDTH(32)) eq_174(.in0(eq_174_in0), .in1(eq_174_in1), .out(eq_174_out));

	reg [31:0] eq_175_in0;
	reg [31:0] eq_175_in1;
	wire [0:0] eq_175_out;
	eq #(.WIDTH(32)) eq_175(.in0(eq_175_in0), .in1(eq_175_in1), .out(eq_175_out));

	reg [31:0] eq_176_in0;
	reg [31:0] eq_176_in1;
	wire [0:0] eq_176_out;
	eq #(.WIDTH(32)) eq_176(.in0(eq_176_in0), .in1(eq_176_in1), .out(eq_176_out));

	reg [31:0] eq_177_in0;
	reg [31:0] eq_177_in1;
	wire [0:0] eq_177_out;
	eq #(.WIDTH(32)) eq_177(.in0(eq_177_in0), .in1(eq_177_in1), .out(eq_177_out));

	reg [0:0] notOp_178_in0;
	wire [0:0] notOp_178_out;
	notOp #(.WIDTH(1)) notOp_178(.in(notOp_178_in0), .out(notOp_178_out));

	reg [0:0] andOp_179_in0;
	reg [0:0] andOp_179_in1;
	wire [0:0] andOp_179_out;
	andOp #(.WIDTH(1)) andOp_179(.in0(andOp_179_in0), .in1(andOp_179_in1), .out(andOp_179_out));

	reg [31:0] eq_180_in0;
	reg [31:0] eq_180_in1;
	wire [0:0] eq_180_out;
	eq #(.WIDTH(32)) eq_180(.in0(eq_180_in0), .in1(eq_180_in1), .out(eq_180_out));

	reg [0:0] notOp_181_in0;
	wire [0:0] notOp_181_out;
	notOp #(.WIDTH(1)) notOp_181(.in(notOp_181_in0), .out(notOp_181_out));

	reg [0:0] andOp_182_in0;
	reg [0:0] andOp_182_in1;
	wire [0:0] andOp_182_out;
	andOp #(.WIDTH(1)) andOp_182(.in0(andOp_182_in0), .in1(andOp_182_in1), .out(andOp_182_out));

	reg [31:0] eq_183_in0;
	reg [31:0] eq_183_in1;
	wire [0:0] eq_183_out;
	eq #(.WIDTH(32)) eq_183(.in0(eq_183_in0), .in1(eq_183_in1), .out(eq_183_out));

	reg [0:0] notOp_184_in0;
	wire [0:0] notOp_184_out;
	notOp #(.WIDTH(1)) notOp_184(.in(notOp_184_in0), .out(notOp_184_out));

	reg [0:0] andOp_185_in0;
	reg [0:0] andOp_185_in1;
	wire [0:0] andOp_185_out;
	andOp #(.WIDTH(1)) andOp_185(.in0(andOp_185_in0), .in1(andOp_185_in1), .out(andOp_185_out));

	reg [31:0] eq_186_in0;
	reg [31:0] eq_186_in1;
	wire [0:0] eq_186_out;
	eq #(.WIDTH(32)) eq_186(.in0(eq_186_in0), .in1(eq_186_in1), .out(eq_186_out));

	reg [0:0] notOp_187_in0;
	wire [0:0] notOp_187_out;
	notOp #(.WIDTH(1)) notOp_187(.in(notOp_187_in0), .out(notOp_187_out));

	reg [0:0] andOp_188_in0;
	reg [0:0] andOp_188_in1;
	wire [0:0] andOp_188_out;
	andOp #(.WIDTH(1)) andOp_188(.in0(andOp_188_in0), .in1(andOp_188_in1), .out(andOp_188_out));

	reg [31:0] eq_189_in0;
	reg [31:0] eq_189_in1;
	wire [0:0] eq_189_out;
	eq #(.WIDTH(32)) eq_189(.in0(eq_189_in0), .in1(eq_189_in1), .out(eq_189_out));

	reg [0:0] notOp_190_in0;
	wire [0:0] notOp_190_out;
	notOp #(.WIDTH(1)) notOp_190(.in(notOp_190_in0), .out(notOp_190_out));

	reg [0:0] andOp_191_in0;
	reg [0:0] andOp_191_in1;
	wire [0:0] andOp_191_out;
	andOp #(.WIDTH(1)) andOp_191(.in0(andOp_191_in0), .in1(andOp_191_in1), .out(andOp_191_out));

	reg [31:0] eq_192_in0;
	reg [31:0] eq_192_in1;
	wire [0:0] eq_192_out;
	eq #(.WIDTH(32)) eq_192(.in0(eq_192_in0), .in1(eq_192_in1), .out(eq_192_out));

	reg [31:0] eq_193_in0;
	reg [31:0] eq_193_in1;
	wire [0:0] eq_193_out;
	eq #(.WIDTH(32)) eq_193(.in0(eq_193_in0), .in1(eq_193_in1), .out(eq_193_out));

	reg [0:0] notOp_194_in0;
	wire [0:0] notOp_194_out;
	notOp #(.WIDTH(1)) notOp_194(.in(notOp_194_in0), .out(notOp_194_out));

	reg [0:0] andOp_195_in0;
	reg [0:0] andOp_195_in1;
	wire [0:0] andOp_195_out;
	andOp #(.WIDTH(1)) andOp_195(.in0(andOp_195_in0), .in1(andOp_195_in1), .out(andOp_195_out));

	reg [0:0] andOp_196_in0;
	reg [0:0] andOp_196_in1;
	wire [0:0] andOp_196_out;
	andOp #(.WIDTH(1)) andOp_196(.in0(andOp_196_in0), .in1(andOp_196_in1), .out(andOp_196_out));

	reg [0:0] andOp_197_in0;
	reg [0:0] andOp_197_in1;
	wire [0:0] andOp_197_out;
	andOp #(.WIDTH(1)) andOp_197(.in0(andOp_197_in0), .in1(andOp_197_in1), .out(andOp_197_out));

	reg [0:0] andOp_198_in0;
	reg [0:0] andOp_198_in1;
	wire [0:0] andOp_198_out;
	andOp #(.WIDTH(1)) andOp_198(.in0(andOp_198_in0), .in1(andOp_198_in1), .out(andOp_198_out));

	reg [0:0] andOp_199_in0;
	reg [0:0] andOp_199_in1;
	wire [0:0] andOp_199_out;
	andOp #(.WIDTH(1)) andOp_199(.in0(andOp_199_in0), .in1(andOp_199_in1), .out(andOp_199_out));

	reg [0:0] andOp_200_in0;
	reg [0:0] andOp_200_in1;
	wire [0:0] andOp_200_out;
	andOp #(.WIDTH(1)) andOp_200(.in0(andOp_200_in0), .in1(andOp_200_in1), .out(andOp_200_out));

	reg [0:0] andOp_201_in0;
	reg [0:0] andOp_201_in1;
	wire [0:0] andOp_201_out;
	andOp #(.WIDTH(1)) andOp_201(.in0(andOp_201_in0), .in1(andOp_201_in1), .out(andOp_201_out));

	reg [0:0] andOp_202_in0;
	reg [0:0] andOp_202_in1;
	wire [0:0] andOp_202_out;
	andOp #(.WIDTH(1)) andOp_202(.in0(andOp_202_in0), .in1(andOp_202_in1), .out(andOp_202_out));

	reg [0:0] andOp_203_in0;
	reg [0:0] andOp_203_in1;
	wire [0:0] andOp_203_out;
	andOp #(.WIDTH(1)) andOp_203(.in0(andOp_203_in0), .in1(andOp_203_in1), .out(andOp_203_out));

	reg [31:0] concat_204_in0;
	reg [31:0] concat_204_in1;
	wire [63:0] concat_204_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_204(.in0(concat_204_in0), .in1(concat_204_in1), .out(concat_204_out));

	reg [31:0] concat_205_in0;
	reg [31:0] concat_205_in1;
	wire [63:0] concat_205_out;
	concat #(.IN0_WIDTH(32), .IN1_WIDTH(32)) concat_205(.in0(concat_205_in0), .in1(concat_205_in1), .out(concat_205_out));

	reg [0:0] andOp_206_in0;
	reg [0:0] andOp_206_in1;
	wire [0:0] andOp_206_out;
	andOp #(.WIDTH(1)) andOp_206(.in0(andOp_206_in0), .in1(andOp_206_in1), .out(andOp_206_out));

	reg [0:0] andOp_207_in0;
	reg [0:0] andOp_207_in1;
	wire [0:0] andOp_207_out;
	andOp #(.WIDTH(1)) andOp_207(.in0(andOp_207_in0), .in1(andOp_207_in1), .out(andOp_207_out));

	reg [0:0] andOp_208_in0;
	reg [0:0] andOp_208_in1;
	wire [0:0] andOp_208_out;
	andOp #(.WIDTH(1)) andOp_208(.in0(andOp_208_in0), .in1(andOp_208_in1), .out(andOp_208_out));

	reg [0:0] andOp_209_in0;
	reg [0:0] andOp_209_in1;
	wire [0:0] andOp_209_out;
	andOp #(.WIDTH(1)) andOp_209(.in0(andOp_209_in0), .in1(andOp_209_in1), .out(andOp_209_out));

	reg [31:0] tmp_output_210_in_data;
	wire [31:0] tmp_output_210_out_data;
	hls_wire #(.WIDTH(32)) tmp_output_210(.in_data(tmp_output_210_in_data), .out_data(tmp_output_210_out_data));

	reg [31:0] eq_211_in0;
	reg [31:0] eq_211_in1;
	wire [0:0] eq_211_out;
	eq #(.WIDTH(32)) eq_211(.in0(eq_211_in0), .in1(eq_211_in1), .out(eq_211_out));

	reg [0:0] andOp_212_in0;
	reg [0:0] andOp_212_in1;
	wire [0:0] andOp_212_out;
	andOp #(.WIDTH(1)) andOp_212(.in0(andOp_212_in0), .in1(andOp_212_in1), .out(andOp_212_out));

	reg [0:0] andOp_213_in0;
	reg [0:0] andOp_213_in1;
	wire [0:0] andOp_213_out;
	andOp #(.WIDTH(1)) andOp_213(.in0(andOp_213_in0), .in1(andOp_213_in1), .out(andOp_213_out));

	reg [0:0] andOp_214_in0;
	reg [0:0] andOp_214_in1;
	wire [0:0] andOp_214_out;
	andOp #(.WIDTH(1)) andOp_214(.in0(andOp_214_in0), .in1(andOp_214_in1), .out(andOp_214_out));

	reg [0:0] andOp_215_in0;
	reg [0:0] andOp_215_in1;
	wire [0:0] andOp_215_out;
	andOp #(.WIDTH(1)) andOp_215(.in0(andOp_215_in0), .in1(andOp_215_in1), .out(andOp_215_out));

	reg [0:0] andOp_216_in0;
	reg [0:0] andOp_216_in1;
	wire [0:0] andOp_216_out;
	andOp #(.WIDTH(1)) andOp_216(.in0(andOp_216_in0), .in1(andOp_216_in1), .out(andOp_216_out));

	reg [0:0] andOp_217_in0;
	reg [0:0] andOp_217_in1;
	wire [0:0] andOp_217_out;
	andOp #(.WIDTH(1)) andOp_217(.in0(andOp_217_in0), .in1(andOp_217_in1), .out(andOp_217_out));

	reg [0:0] andOp_218_in0;
	reg [0:0] andOp_218_in1;
	wire [0:0] andOp_218_out;
	andOp #(.WIDTH(1)) andOp_218(.in0(andOp_218_in0), .in1(andOp_218_in1), .out(andOp_218_out));

	reg [0:0] andOp_219_in0;
	reg [0:0] andOp_219_in1;
	wire [0:0] andOp_219_out;
	andOp #(.WIDTH(1)) andOp_219(.in0(andOp_219_in0), .in1(andOp_219_in1), .out(andOp_219_out));

	reg [0:0] andOp_220_in0;
	reg [0:0] andOp_220_in1;
	wire [0:0] andOp_220_out;
	andOp #(.WIDTH(1)) andOp_220(.in0(andOp_220_in0), .in1(andOp_220_in1), .out(andOp_220_out));

	reg [0:0] andOp_221_in0;
	reg [0:0] andOp_221_in1;
	wire [0:0] andOp_221_out;
	andOp #(.WIDTH(1)) andOp_221(.in0(andOp_221_in0), .in1(andOp_221_in1), .out(andOp_221_out));

	reg [0:0] andOp_222_in0;
	reg [0:0] andOp_222_in1;
	wire [0:0] andOp_222_out;
	andOp #(.WIDTH(1)) andOp_222(.in0(andOp_222_in0), .in1(andOp_222_in1), .out(andOp_222_out));

	reg [0:0] notOp_223_in0;
	wire [0:0] notOp_223_out;
	notOp #(.WIDTH(1)) notOp_223(.in(notOp_223_in0), .out(notOp_223_out));

	reg [0:0] andOp_224_in0;
	reg [0:0] andOp_224_in1;
	wire [0:0] andOp_224_out;
	andOp #(.WIDTH(1)) andOp_224(.in0(andOp_224_in0), .in1(andOp_224_in1), .out(andOp_224_out));

	reg [0:0] notOp_225_in0;
	wire [0:0] notOp_225_out;
	notOp #(.WIDTH(1)) notOp_225(.in(notOp_225_in0), .out(notOp_225_out));

	reg [0:0] andOp_226_in0;
	reg [0:0] andOp_226_in1;
	wire [0:0] andOp_226_out;
	andOp #(.WIDTH(1)) andOp_226(.in0(andOp_226_in0), .in1(andOp_226_in1), .out(andOp_226_out));

	reg [0:0] notOp_227_in0;
	wire [0:0] notOp_227_out;
	notOp #(.WIDTH(1)) notOp_227(.in(notOp_227_in0), .out(notOp_227_out));

	reg [0:0] andOp_228_in0;
	reg [0:0] andOp_228_in1;
	wire [0:0] andOp_228_out;
	andOp #(.WIDTH(1)) andOp_228(.in0(andOp_228_in0), .in1(andOp_228_in1), .out(andOp_228_out));

	reg [0:0] notOp_229_in0;
	wire [0:0] notOp_229_out;
	notOp #(.WIDTH(1)) notOp_229(.in(notOp_229_in0), .out(notOp_229_out));

	reg [0:0] andOp_230_in0;
	reg [0:0] andOp_230_in1;
	wire [0:0] andOp_230_out;
	andOp #(.WIDTH(1)) andOp_230(.in0(andOp_230_in0), .in1(andOp_230_in1), .out(andOp_230_out));

	reg [0:0] notOp_231_in0;
	wire [0:0] notOp_231_out;
	notOp #(.WIDTH(1)) notOp_231(.in(notOp_231_in0), .out(notOp_231_out));

	reg [0:0] andOp_232_in0;
	reg [0:0] andOp_232_in1;
	wire [0:0] andOp_232_out;
	andOp #(.WIDTH(1)) andOp_232(.in0(andOp_232_in0), .in1(andOp_232_in1), .out(andOp_232_out));

	reg [0:0] notOp_233_in0;
	wire [0:0] notOp_233_out;
	notOp #(.WIDTH(1)) notOp_233(.in(notOp_233_in0), .out(notOp_233_out));

	reg [0:0] andOp_234_in0;
	reg [0:0] andOp_234_in1;
	wire [0:0] andOp_234_out;
	andOp #(.WIDTH(1)) andOp_234(.in0(andOp_234_in0), .in1(andOp_234_in1), .out(andOp_234_out));

	reg [0:0] notOp_235_in0;
	wire [0:0] notOp_235_out;
	notOp #(.WIDTH(1)) notOp_235(.in(notOp_235_in0), .out(notOp_235_out));

	reg [0:0] andOp_236_in0;
	reg [0:0] andOp_236_in1;
	wire [0:0] andOp_236_out;
	andOp #(.WIDTH(1)) andOp_236(.in0(andOp_236_in0), .in1(andOp_236_in1), .out(andOp_236_out));

	reg [0:0] notOp_237_in0;
	wire [0:0] notOp_237_out;
	notOp #(.WIDTH(1)) notOp_237(.in(notOp_237_in0), .out(notOp_237_out));

	reg [0:0] andOp_238_in0;
	reg [0:0] andOp_238_in1;
	wire [0:0] andOp_238_out;
	andOp #(.WIDTH(1)) andOp_238(.in0(andOp_238_in0), .in1(andOp_238_in1), .out(andOp_238_out));

	reg [0:0] andOp_239_in0;
	reg [0:0] andOp_239_in1;
	wire [0:0] andOp_239_out;
	andOp #(.WIDTH(1)) andOp_239(.in0(andOp_239_in0), .in1(andOp_239_in1), .out(andOp_239_out));

	reg [0:0] andOp_240_in0;
	reg [0:0] andOp_240_in1;
	wire [0:0] andOp_240_out;
	andOp #(.WIDTH(1)) andOp_240(.in0(andOp_240_in0), .in1(andOp_240_in1), .out(andOp_240_out));

	reg [0:0] andOp_241_in0;
	reg [0:0] andOp_241_in1;
	wire [0:0] andOp_241_out;
	andOp #(.WIDTH(1)) andOp_241(.in0(andOp_241_in0), .in1(andOp_241_in1), .out(andOp_241_out));

	reg [0:0] andOp_242_in0;
	reg [0:0] andOp_242_in1;
	wire [0:0] andOp_242_out;
	andOp #(.WIDTH(1)) andOp_242(.in0(andOp_242_in0), .in1(andOp_242_in1), .out(andOp_242_out));

	reg [31:0] eq_243_in0;
	reg [31:0] eq_243_in1;
	wire [0:0] eq_243_out;
	eq #(.WIDTH(32)) eq_243(.in0(eq_243_in0), .in1(eq_243_in1), .out(eq_243_out));

	reg [0:0] andOp_244_in0;
	reg [0:0] andOp_244_in1;
	wire [0:0] andOp_244_out;
	andOp #(.WIDTH(1)) andOp_244(.in0(andOp_244_in0), .in1(andOp_244_in1), .out(andOp_244_out));

	reg [31:0] eq_245_in0;
	reg [31:0] eq_245_in1;
	wire [0:0] eq_245_out;
	eq #(.WIDTH(32)) eq_245(.in0(eq_245_in0), .in1(eq_245_in1), .out(eq_245_out));

	reg [0:0] andOp_246_in0;
	reg [0:0] andOp_246_in1;
	wire [0:0] andOp_246_out;
	andOp #(.WIDTH(1)) andOp_246(.in0(andOp_246_in0), .in1(andOp_246_in1), .out(andOp_246_out));

	reg [31:0] eq_247_in0;
	reg [31:0] eq_247_in1;
	wire [0:0] eq_247_out;
	eq #(.WIDTH(32)) eq_247(.in0(eq_247_in0), .in1(eq_247_in1), .out(eq_247_out));

	reg [0:0] andOp_248_in0;
	reg [0:0] andOp_248_in1;
	wire [0:0] andOp_248_out;
	andOp #(.WIDTH(1)) andOp_248(.in0(andOp_248_in0), .in1(andOp_248_in1), .out(andOp_248_out));

	reg [31:0] eq_249_in0;
	reg [31:0] eq_249_in1;
	wire [0:0] eq_249_out;
	eq #(.WIDTH(32)) eq_249(.in0(eq_249_in0), .in1(eq_249_in1), .out(eq_249_out));

	reg [0:0] andOp_250_in0;
	reg [0:0] andOp_250_in1;
	wire [0:0] andOp_250_out;
	andOp #(.WIDTH(1)) andOp_250(.in0(andOp_250_in0), .in1(andOp_250_in1), .out(andOp_250_out));

	reg [31:0] eq_251_in0;
	reg [31:0] eq_251_in1;
	wire [0:0] eq_251_out;
	eq #(.WIDTH(32)) eq_251(.in0(eq_251_in0), .in1(eq_251_in1), .out(eq_251_out));

	reg [0:0] andOp_252_in0;
	reg [0:0] andOp_252_in1;
	wire [0:0] andOp_252_out;
	andOp #(.WIDTH(1)) andOp_252(.in0(andOp_252_in0), .in1(andOp_252_in1), .out(andOp_252_out));

	reg [0:0] andOp_253_in0;
	reg [0:0] andOp_253_in1;
	wire [0:0] andOp_253_out;
	andOp #(.WIDTH(1)) andOp_253(.in0(andOp_253_in0), .in1(andOp_253_in1), .out(andOp_253_out));

	reg [31:0] eq_254_in0;
	reg [31:0] eq_254_in1;
	wire [0:0] eq_254_out;
	eq #(.WIDTH(32)) eq_254(.in0(eq_254_in0), .in1(eq_254_in1), .out(eq_254_out));

	reg [0:0] andOp_255_in0;
	reg [0:0] andOp_255_in1;
	wire [0:0] andOp_255_out;
	andOp #(.WIDTH(1)) andOp_255(.in0(andOp_255_in0), .in1(andOp_255_in1), .out(andOp_255_out));

	reg [0:0] notOp_256_in0;
	wire [0:0] notOp_256_out;
	notOp #(.WIDTH(1)) notOp_256(.in(notOp_256_in0), .out(notOp_256_out));

	reg [0:0] andOp_257_in0;
	reg [0:0] andOp_257_in1;
	wire [0:0] andOp_257_out;
	andOp #(.WIDTH(1)) andOp_257(.in0(andOp_257_in0), .in1(andOp_257_in1), .out(andOp_257_out));

	reg [0:0] andOp_258_in0;
	reg [0:0] andOp_258_in1;
	wire [0:0] andOp_258_out;
	andOp #(.WIDTH(1)) andOp_258(.in0(andOp_258_in0), .in1(andOp_258_in1), .out(andOp_258_out));

	reg [31:0] eq_259_in0;
	reg [31:0] eq_259_in1;
	wire [0:0] eq_259_out;
	eq #(.WIDTH(32)) eq_259(.in0(eq_259_in0), .in1(eq_259_in1), .out(eq_259_out));

	reg [0:0] andOp_260_in0;
	reg [0:0] andOp_260_in1;
	wire [0:0] andOp_260_out;
	andOp #(.WIDTH(1)) andOp_260(.in0(andOp_260_in0), .in1(andOp_260_in1), .out(andOp_260_out));

	reg [0:0] notOp_261_in0;
	wire [0:0] notOp_261_out;
	notOp #(.WIDTH(1)) notOp_261(.in(notOp_261_in0), .out(notOp_261_out));

	reg [0:0] andOp_262_in0;
	reg [0:0] andOp_262_in1;
	wire [0:0] andOp_262_out;
	andOp #(.WIDTH(1)) andOp_262(.in0(andOp_262_in0), .in1(andOp_262_in1), .out(andOp_262_out));

	reg [0:0] andOp_263_in0;
	reg [0:0] andOp_263_in1;
	wire [0:0] andOp_263_out;
	andOp #(.WIDTH(1)) andOp_263(.in0(andOp_263_in0), .in1(andOp_263_in1), .out(andOp_263_out));

	reg [31:0] eq_264_in0;
	reg [31:0] eq_264_in1;
	wire [0:0] eq_264_out;
	eq #(.WIDTH(32)) eq_264(.in0(eq_264_in0), .in1(eq_264_in1), .out(eq_264_out));

	reg [0:0] andOp_265_in0;
	reg [0:0] andOp_265_in1;
	wire [0:0] andOp_265_out;
	andOp #(.WIDTH(1)) andOp_265(.in0(andOp_265_in0), .in1(andOp_265_in1), .out(andOp_265_out));

	reg [0:0] notOp_266_in0;
	wire [0:0] notOp_266_out;
	notOp #(.WIDTH(1)) notOp_266(.in(notOp_266_in0), .out(notOp_266_out));

	reg [0:0] andOp_267_in0;
	reg [0:0] andOp_267_in1;
	wire [0:0] andOp_267_out;
	andOp #(.WIDTH(1)) andOp_267(.in0(andOp_267_in0), .in1(andOp_267_in1), .out(andOp_267_out));

	reg [0:0] andOp_268_in0;
	reg [0:0] andOp_268_in1;
	wire [0:0] andOp_268_out;
	andOp #(.WIDTH(1)) andOp_268(.in0(andOp_268_in0), .in1(andOp_268_in1), .out(andOp_268_out));

	reg [31:0] eq_269_in0;
	reg [31:0] eq_269_in1;
	wire [0:0] eq_269_out;
	eq #(.WIDTH(32)) eq_269(.in0(eq_269_in0), .in1(eq_269_in1), .out(eq_269_out));

	reg [0:0] andOp_270_in0;
	reg [0:0] andOp_270_in1;
	wire [0:0] andOp_270_out;
	andOp #(.WIDTH(1)) andOp_270(.in0(andOp_270_in0), .in1(andOp_270_in1), .out(andOp_270_out));

	reg [0:0] notOp_271_in0;
	wire [0:0] notOp_271_out;
	notOp #(.WIDTH(1)) notOp_271(.in(notOp_271_in0), .out(notOp_271_out));

	reg [0:0] andOp_272_in0;
	reg [0:0] andOp_272_in1;
	wire [0:0] andOp_272_out;
	andOp #(.WIDTH(1)) andOp_272(.in0(andOp_272_in0), .in1(andOp_272_in1), .out(andOp_272_out));

	reg [0:0] andOp_273_in0;
	reg [0:0] andOp_273_in1;
	wire [0:0] andOp_273_out;
	andOp #(.WIDTH(1)) andOp_273(.in0(andOp_273_in0), .in1(andOp_273_in1), .out(andOp_273_out));

	reg [31:0] eq_274_in0;
	reg [31:0] eq_274_in1;
	wire [0:0] eq_274_out;
	eq #(.WIDTH(32)) eq_274(.in0(eq_274_in0), .in1(eq_274_in1), .out(eq_274_out));

	reg [0:0] andOp_275_in0;
	reg [0:0] andOp_275_in1;
	wire [0:0] andOp_275_out;
	andOp #(.WIDTH(1)) andOp_275(.in0(andOp_275_in0), .in1(andOp_275_in1), .out(andOp_275_out));

	reg [0:0] notOp_276_in0;
	wire [0:0] notOp_276_out;
	notOp #(.WIDTH(1)) notOp_276(.in(notOp_276_in0), .out(notOp_276_out));

	reg [0:0] andOp_277_in0;
	reg [0:0] andOp_277_in1;
	wire [0:0] andOp_277_out;
	andOp #(.WIDTH(1)) andOp_277(.in0(andOp_277_in0), .in1(andOp_277_in1), .out(andOp_277_out));

	reg [0:0] andOp_278_in0;
	reg [0:0] andOp_278_in1;
	wire [0:0] andOp_278_out;
	andOp #(.WIDTH(1)) andOp_278(.in0(andOp_278_in0), .in1(andOp_278_in1), .out(andOp_278_out));

	reg [31:0] eq_279_in0;
	reg [31:0] eq_279_in1;
	wire [0:0] eq_279_out;
	eq #(.WIDTH(32)) eq_279(.in0(eq_279_in0), .in1(eq_279_in1), .out(eq_279_out));

	reg [0:0] andOp_280_in0;
	reg [0:0] andOp_280_in1;
	wire [0:0] andOp_280_out;
	andOp #(.WIDTH(1)) andOp_280(.in0(andOp_280_in0), .in1(andOp_280_in1), .out(andOp_280_out));

	reg [0:0] notOp_281_in0;
	wire [0:0] notOp_281_out;
	notOp #(.WIDTH(1)) notOp_281(.in(notOp_281_in0), .out(notOp_281_out));

	reg [0:0] andOp_282_in0;
	reg [0:0] andOp_282_in1;
	wire [0:0] andOp_282_out;
	andOp #(.WIDTH(1)) andOp_282(.in0(andOp_282_in0), .in1(andOp_282_in1), .out(andOp_282_out));

	reg [0:0] andOp_283_in0;
	reg [0:0] andOp_283_in1;
	wire [0:0] andOp_283_out;
	andOp #(.WIDTH(1)) andOp_283(.in0(andOp_283_in0), .in1(andOp_283_in1), .out(andOp_283_out));

	reg [31:0] eq_284_in0;
	reg [31:0] eq_284_in1;
	wire [0:0] eq_284_out;
	eq #(.WIDTH(32)) eq_284(.in0(eq_284_in0), .in1(eq_284_in1), .out(eq_284_out));

	reg [0:0] andOp_285_in0;
	reg [0:0] andOp_285_in1;
	wire [0:0] andOp_285_out;
	andOp #(.WIDTH(1)) andOp_285(.in0(andOp_285_in0), .in1(andOp_285_in1), .out(andOp_285_out));

	reg [0:0] notOp_286_in0;
	wire [0:0] notOp_286_out;
	notOp #(.WIDTH(1)) notOp_286(.in(notOp_286_in0), .out(notOp_286_out));

	reg [0:0] andOp_287_in0;
	reg [0:0] andOp_287_in1;
	wire [0:0] andOp_287_out;
	andOp #(.WIDTH(1)) andOp_287(.in0(andOp_287_in0), .in1(andOp_287_in1), .out(andOp_287_out));

	reg [0:0] andOp_288_in0;
	reg [0:0] andOp_288_in1;
	wire [0:0] andOp_288_out;
	andOp #(.WIDTH(1)) andOp_288(.in0(andOp_288_in0), .in1(andOp_288_in1), .out(andOp_288_out));

	reg [31:0] eq_289_in0;
	reg [31:0] eq_289_in1;
	wire [0:0] eq_289_out;
	eq #(.WIDTH(32)) eq_289(.in0(eq_289_in0), .in1(eq_289_in1), .out(eq_289_out));

	reg [0:0] andOp_290_in0;
	reg [0:0] andOp_290_in1;
	wire [0:0] andOp_290_out;
	andOp #(.WIDTH(1)) andOp_290(.in0(andOp_290_in0), .in1(andOp_290_in1), .out(andOp_290_out));

	reg [0:0] notOp_291_in0;
	wire [0:0] notOp_291_out;
	notOp #(.WIDTH(1)) notOp_291(.in(notOp_291_in0), .out(notOp_291_out));

	reg [0:0] andOp_292_in0;
	reg [0:0] andOp_292_in1;
	wire [0:0] andOp_292_out;
	andOp #(.WIDTH(1)) andOp_292(.in0(andOp_292_in0), .in1(andOp_292_in1), .out(andOp_292_out));

	reg [0:0] andOp_293_in0;
	reg [0:0] andOp_293_in1;
	wire [0:0] andOp_293_out;
	andOp #(.WIDTH(1)) andOp_293(.in0(andOp_293_in0), .in1(andOp_293_in1), .out(andOp_293_out));

	reg [31:0] eq_294_in0;
	reg [31:0] eq_294_in1;
	wire [0:0] eq_294_out;
	eq #(.WIDTH(32)) eq_294(.in0(eq_294_in0), .in1(eq_294_in1), .out(eq_294_out));

	reg [0:0] andOp_295_in0;
	reg [0:0] andOp_295_in1;
	wire [0:0] andOp_295_out;
	andOp #(.WIDTH(1)) andOp_295(.in0(andOp_295_in0), .in1(andOp_295_in1), .out(andOp_295_out));

	reg [0:0] notOp_296_in0;
	wire [0:0] notOp_296_out;
	notOp #(.WIDTH(1)) notOp_296(.in(notOp_296_in0), .out(notOp_296_out));

	reg [0:0] andOp_297_in0;
	reg [0:0] andOp_297_in1;
	wire [0:0] andOp_297_out;
	andOp #(.WIDTH(1)) andOp_297(.in0(andOp_297_in0), .in1(andOp_297_in1), .out(andOp_297_out));

	reg [31:0] eq_298_in0;
	reg [31:0] eq_298_in1;
	wire [0:0] eq_298_out;
	eq #(.WIDTH(32)) eq_298(.in0(eq_298_in0), .in1(eq_298_in1), .out(eq_298_out));

	reg [0:0] andOp_299_in0;
	reg [0:0] andOp_299_in1;
	wire [0:0] andOp_299_out;
	andOp #(.WIDTH(1)) andOp_299(.in0(andOp_299_in0), .in1(andOp_299_in1), .out(andOp_299_out));

	reg [31:0] eq_300_in0;
	reg [31:0] eq_300_in1;
	wire [0:0] eq_300_out;
	eq #(.WIDTH(32)) eq_300(.in0(eq_300_in0), .in1(eq_300_in1), .out(eq_300_out));

	reg [0:0] andOp_301_in0;
	reg [0:0] andOp_301_in1;
	wire [0:0] andOp_301_out;
	andOp #(.WIDTH(1)) andOp_301(.in0(andOp_301_in0), .in1(andOp_301_in1), .out(andOp_301_out));

	reg [31:0] eq_302_in0;
	reg [31:0] eq_302_in1;
	wire [0:0] eq_302_out;
	eq #(.WIDTH(32)) eq_302(.in0(eq_302_in0), .in1(eq_302_in1), .out(eq_302_out));

	reg [0:0] andOp_303_in0;
	reg [0:0] andOp_303_in1;
	wire [0:0] andOp_303_out;
	andOp #(.WIDTH(1)) andOp_303(.in0(andOp_303_in0), .in1(andOp_303_in1), .out(andOp_303_out));

	reg [31:0] eq_304_in0;
	reg [31:0] eq_304_in1;
	wire [0:0] eq_304_out;
	eq #(.WIDTH(32)) eq_304(.in0(eq_304_in0), .in1(eq_304_in1), .out(eq_304_out));

	reg [0:0] andOp_305_in0;
	reg [0:0] andOp_305_in1;
	wire [0:0] andOp_305_out;
	andOp #(.WIDTH(1)) andOp_305(.in0(andOp_305_in0), .in1(andOp_305_in1), .out(andOp_305_out));

	reg [31:0] eq_306_in0;
	reg [31:0] eq_306_in1;
	wire [0:0] eq_306_out;
	eq #(.WIDTH(32)) eq_306(.in0(eq_306_in0), .in1(eq_306_in1), .out(eq_306_out));

	reg [0:0] andOp_307_in0;
	reg [0:0] andOp_307_in1;
	wire [0:0] andOp_307_out;
	andOp #(.WIDTH(1)) andOp_307(.in0(andOp_307_in0), .in1(andOp_307_in1), .out(andOp_307_out));

	reg [0:0] andOp_308_in0;
	reg [0:0] andOp_308_in1;
	wire [0:0] andOp_308_out;
	andOp #(.WIDTH(1)) andOp_308(.in0(andOp_308_in0), .in1(andOp_308_in1), .out(andOp_308_out));

	reg [31:0] eq_309_in0;
	reg [31:0] eq_309_in1;
	wire [0:0] eq_309_out;
	eq #(.WIDTH(32)) eq_309(.in0(eq_309_in0), .in1(eq_309_in1), .out(eq_309_out));

	reg [0:0] andOp_310_in0;
	reg [0:0] andOp_310_in1;
	wire [0:0] andOp_310_out;
	andOp #(.WIDTH(1)) andOp_310(.in0(andOp_310_in0), .in1(andOp_310_in1), .out(andOp_310_out));

	reg [0:0] notOp_311_in0;
	wire [0:0] notOp_311_out;
	notOp #(.WIDTH(1)) notOp_311(.in(notOp_311_in0), .out(notOp_311_out));

	reg [0:0] andOp_312_in0;
	reg [0:0] andOp_312_in1;
	wire [0:0] andOp_312_out;
	andOp #(.WIDTH(1)) andOp_312(.in0(andOp_312_in0), .in1(andOp_312_in1), .out(andOp_312_out));

	reg [0:0] andOp_313_in0;
	reg [0:0] andOp_313_in1;
	wire [0:0] andOp_313_out;
	andOp #(.WIDTH(1)) andOp_313(.in0(andOp_313_in0), .in1(andOp_313_in1), .out(andOp_313_out));

	reg [31:0] eq_314_in0;
	reg [31:0] eq_314_in1;
	wire [0:0] eq_314_out;
	eq #(.WIDTH(32)) eq_314(.in0(eq_314_in0), .in1(eq_314_in1), .out(eq_314_out));

	reg [0:0] andOp_315_in0;
	reg [0:0] andOp_315_in1;
	wire [0:0] andOp_315_out;
	andOp #(.WIDTH(1)) andOp_315(.in0(andOp_315_in0), .in1(andOp_315_in1), .out(andOp_315_out));

	reg [0:0] notOp_316_in0;
	wire [0:0] notOp_316_out;
	notOp #(.WIDTH(1)) notOp_316(.in(notOp_316_in0), .out(notOp_316_out));

	reg [0:0] andOp_317_in0;
	reg [0:0] andOp_317_in1;
	wire [0:0] andOp_317_out;
	andOp #(.WIDTH(1)) andOp_317(.in0(andOp_317_in0), .in1(andOp_317_in1), .out(andOp_317_out));

	reg [0:0] andOp_318_in0;
	reg [0:0] andOp_318_in1;
	wire [0:0] andOp_318_out;
	andOp #(.WIDTH(1)) andOp_318(.in0(andOp_318_in0), .in1(andOp_318_in1), .out(andOp_318_out));

	reg [31:0] eq_319_in0;
	reg [31:0] eq_319_in1;
	wire [0:0] eq_319_out;
	eq #(.WIDTH(32)) eq_319(.in0(eq_319_in0), .in1(eq_319_in1), .out(eq_319_out));

	reg [0:0] andOp_320_in0;
	reg [0:0] andOp_320_in1;
	wire [0:0] andOp_320_out;
	andOp #(.WIDTH(1)) andOp_320(.in0(andOp_320_in0), .in1(andOp_320_in1), .out(andOp_320_out));

	reg [0:0] notOp_321_in0;
	wire [0:0] notOp_321_out;
	notOp #(.WIDTH(1)) notOp_321(.in(notOp_321_in0), .out(notOp_321_out));

	reg [0:0] andOp_322_in0;
	reg [0:0] andOp_322_in1;
	wire [0:0] andOp_322_out;
	andOp #(.WIDTH(1)) andOp_322(.in0(andOp_322_in0), .in1(andOp_322_in1), .out(andOp_322_out));

	reg [0:0] andOp_323_in0;
	reg [0:0] andOp_323_in1;
	wire [0:0] andOp_323_out;
	andOp #(.WIDTH(1)) andOp_323(.in0(andOp_323_in0), .in1(andOp_323_in1), .out(andOp_323_out));

	reg [31:0] eq_324_in0;
	reg [31:0] eq_324_in1;
	wire [0:0] eq_324_out;
	eq #(.WIDTH(32)) eq_324(.in0(eq_324_in0), .in1(eq_324_in1), .out(eq_324_out));

	reg [0:0] andOp_325_in0;
	reg [0:0] andOp_325_in1;
	wire [0:0] andOp_325_out;
	andOp #(.WIDTH(1)) andOp_325(.in0(andOp_325_in0), .in1(andOp_325_in1), .out(andOp_325_out));

	reg [0:0] notOp_326_in0;
	wire [0:0] notOp_326_out;
	notOp #(.WIDTH(1)) notOp_326(.in(notOp_326_in0), .out(notOp_326_out));

	reg [0:0] andOp_327_in0;
	reg [0:0] andOp_327_in1;
	wire [0:0] andOp_327_out;
	andOp #(.WIDTH(1)) andOp_327(.in0(andOp_327_in0), .in1(andOp_327_in1), .out(andOp_327_out));

	reg [0:0] andOp_328_in0;
	reg [0:0] andOp_328_in1;
	wire [0:0] andOp_328_out;
	andOp #(.WIDTH(1)) andOp_328(.in0(andOp_328_in0), .in1(andOp_328_in1), .out(andOp_328_out));

	reg [31:0] eq_329_in0;
	reg [31:0] eq_329_in1;
	wire [0:0] eq_329_out;
	eq #(.WIDTH(32)) eq_329(.in0(eq_329_in0), .in1(eq_329_in1), .out(eq_329_out));

	reg [0:0] andOp_330_in0;
	reg [0:0] andOp_330_in1;
	wire [0:0] andOp_330_out;
	andOp #(.WIDTH(1)) andOp_330(.in0(andOp_330_in0), .in1(andOp_330_in1), .out(andOp_330_out));

	reg [0:0] notOp_331_in0;
	wire [0:0] notOp_331_out;
	notOp #(.WIDTH(1)) notOp_331(.in(notOp_331_in0), .out(notOp_331_out));

	reg [0:0] andOp_332_in0;
	reg [0:0] andOp_332_in1;
	wire [0:0] andOp_332_out;
	andOp #(.WIDTH(1)) andOp_332(.in0(andOp_332_in0), .in1(andOp_332_in1), .out(andOp_332_out));

	reg [0:0] andOp_333_in0;
	reg [0:0] andOp_333_in1;
	wire [0:0] andOp_333_out;
	andOp #(.WIDTH(1)) andOp_333(.in0(andOp_333_in0), .in1(andOp_333_in1), .out(andOp_333_out));

	reg [31:0] eq_334_in0;
	reg [31:0] eq_334_in1;
	wire [0:0] eq_334_out;
	eq #(.WIDTH(32)) eq_334(.in0(eq_334_in0), .in1(eq_334_in1), .out(eq_334_out));

	reg [0:0] andOp_335_in0;
	reg [0:0] andOp_335_in1;
	wire [0:0] andOp_335_out;
	andOp #(.WIDTH(1)) andOp_335(.in0(andOp_335_in0), .in1(andOp_335_in1), .out(andOp_335_out));

	reg [0:0] notOp_336_in0;
	wire [0:0] notOp_336_out;
	notOp #(.WIDTH(1)) notOp_336(.in(notOp_336_in0), .out(notOp_336_out));

	reg [0:0] andOp_337_in0;
	reg [0:0] andOp_337_in1;
	wire [0:0] andOp_337_out;
	andOp #(.WIDTH(1)) andOp_337(.in0(andOp_337_in0), .in1(andOp_337_in1), .out(andOp_337_out));

	reg [0:0] andOp_338_in0;
	reg [0:0] andOp_338_in1;
	wire [0:0] andOp_338_out;
	andOp #(.WIDTH(1)) andOp_338(.in0(andOp_338_in0), .in1(andOp_338_in1), .out(andOp_338_out));

	reg [31:0] eq_339_in0;
	reg [31:0] eq_339_in1;
	wire [0:0] eq_339_out;
	eq #(.WIDTH(32)) eq_339(.in0(eq_339_in0), .in1(eq_339_in1), .out(eq_339_out));

	reg [0:0] andOp_340_in0;
	reg [0:0] andOp_340_in1;
	wire [0:0] andOp_340_out;
	andOp #(.WIDTH(1)) andOp_340(.in0(andOp_340_in0), .in1(andOp_340_in1), .out(andOp_340_out));

	reg [0:0] notOp_341_in0;
	wire [0:0] notOp_341_out;
	notOp #(.WIDTH(1)) notOp_341(.in(notOp_341_in0), .out(notOp_341_out));

	reg [0:0] andOp_342_in0;
	reg [0:0] andOp_342_in1;
	wire [0:0] andOp_342_out;
	andOp #(.WIDTH(1)) andOp_342(.in0(andOp_342_in0), .in1(andOp_342_in1), .out(andOp_342_out));

	reg [0:0] andOp_343_in0;
	reg [0:0] andOp_343_in1;
	wire [0:0] andOp_343_out;
	andOp #(.WIDTH(1)) andOp_343(.in0(andOp_343_in0), .in1(andOp_343_in1), .out(andOp_343_out));

	reg [31:0] eq_344_in0;
	reg [31:0] eq_344_in1;
	wire [0:0] eq_344_out;
	eq #(.WIDTH(32)) eq_344(.in0(eq_344_in0), .in1(eq_344_in1), .out(eq_344_out));

	reg [0:0] andOp_345_in0;
	reg [0:0] andOp_345_in1;
	wire [0:0] andOp_345_out;
	andOp #(.WIDTH(1)) andOp_345(.in0(andOp_345_in0), .in1(andOp_345_in1), .out(andOp_345_out));

	reg [0:0] notOp_346_in0;
	wire [0:0] notOp_346_out;
	notOp #(.WIDTH(1)) notOp_346(.in(notOp_346_in0), .out(notOp_346_out));

	reg [0:0] andOp_347_in0;
	reg [0:0] andOp_347_in1;
	wire [0:0] andOp_347_out;
	andOp #(.WIDTH(1)) andOp_347(.in0(andOp_347_in0), .in1(andOp_347_in1), .out(andOp_347_out));

	reg [0:0] andOp_348_in0;
	reg [0:0] andOp_348_in1;
	wire [0:0] andOp_348_out;
	andOp #(.WIDTH(1)) andOp_348(.in0(andOp_348_in0), .in1(andOp_348_in1), .out(andOp_348_out));

	reg [31:0] eq_349_in0;
	reg [31:0] eq_349_in1;
	wire [0:0] eq_349_out;
	eq #(.WIDTH(32)) eq_349(.in0(eq_349_in0), .in1(eq_349_in1), .out(eq_349_out));

	reg [0:0] andOp_350_in0;
	reg [0:0] andOp_350_in1;
	wire [0:0] andOp_350_out;
	andOp #(.WIDTH(1)) andOp_350(.in0(andOp_350_in0), .in1(andOp_350_in1), .out(andOp_350_out));

	reg [0:0] notOp_351_in0;
	wire [0:0] notOp_351_out;
	notOp #(.WIDTH(1)) notOp_351(.in(notOp_351_in0), .out(notOp_351_out));

	reg [0:0] andOp_352_in0;
	reg [0:0] andOp_352_in1;
	wire [0:0] andOp_352_out;
	andOp #(.WIDTH(1)) andOp_352(.in0(andOp_352_in0), .in1(andOp_352_in1), .out(andOp_352_out));

	reg [31:0] eq_353_in0;
	reg [31:0] eq_353_in1;
	wire [0:0] eq_353_out;
	eq #(.WIDTH(32)) eq_353(.in0(eq_353_in0), .in1(eq_353_in1), .out(eq_353_out));

	reg [0:0] andOp_354_in0;
	reg [0:0] andOp_354_in1;
	wire [0:0] andOp_354_out;
	andOp #(.WIDTH(1)) andOp_354(.in0(andOp_354_in0), .in1(andOp_354_in1), .out(andOp_354_out));

	reg [31:0] eq_355_in0;
	reg [31:0] eq_355_in1;
	wire [0:0] eq_355_out;
	eq #(.WIDTH(32)) eq_355(.in0(eq_355_in0), .in1(eq_355_in1), .out(eq_355_out));

	reg [0:0] andOp_356_in0;
	reg [0:0] andOp_356_in1;
	wire [0:0] andOp_356_out;
	andOp #(.WIDTH(1)) andOp_356(.in0(andOp_356_in0), .in1(andOp_356_in1), .out(andOp_356_out));

	reg [31:0] eq_357_in0;
	reg [31:0] eq_357_in1;
	wire [0:0] eq_357_out;
	eq #(.WIDTH(32)) eq_357(.in0(eq_357_in0), .in1(eq_357_in1), .out(eq_357_out));

	reg [0:0] andOp_358_in0;
	reg [0:0] andOp_358_in1;
	wire [0:0] andOp_358_out;
	andOp #(.WIDTH(1)) andOp_358(.in0(andOp_358_in0), .in1(andOp_358_in1), .out(andOp_358_out));

	reg [31:0] eq_359_in0;
	reg [31:0] eq_359_in1;
	wire [0:0] eq_359_out;
	eq #(.WIDTH(32)) eq_359(.in0(eq_359_in0), .in1(eq_359_in1), .out(eq_359_out));

	reg [0:0] andOp_360_in0;
	reg [0:0] andOp_360_in1;
	wire [0:0] andOp_360_out;
	andOp #(.WIDTH(1)) andOp_360(.in0(andOp_360_in0), .in1(andOp_360_in1), .out(andOp_360_out));

	reg [31:0] eq_361_in0;
	reg [31:0] eq_361_in1;
	wire [0:0] eq_361_out;
	eq #(.WIDTH(32)) eq_361(.in0(eq_361_in0), .in1(eq_361_in1), .out(eq_361_out));

	reg [0:0] andOp_362_in0;
	reg [0:0] andOp_362_in1;
	wire [0:0] andOp_362_out;
	andOp #(.WIDTH(1)) andOp_362(.in0(andOp_362_in0), .in1(andOp_362_in1), .out(andOp_362_out));

	reg [0:0] andOp_363_in0;
	reg [0:0] andOp_363_in1;
	wire [0:0] andOp_363_out;
	andOp #(.WIDTH(1)) andOp_363(.in0(andOp_363_in0), .in1(andOp_363_in1), .out(andOp_363_out));

	reg [31:0] eq_364_in0;
	reg [31:0] eq_364_in1;
	wire [0:0] eq_364_out;
	eq #(.WIDTH(32)) eq_364(.in0(eq_364_in0), .in1(eq_364_in1), .out(eq_364_out));

	reg [0:0] andOp_365_in0;
	reg [0:0] andOp_365_in1;
	wire [0:0] andOp_365_out;
	andOp #(.WIDTH(1)) andOp_365(.in0(andOp_365_in0), .in1(andOp_365_in1), .out(andOp_365_out));

	reg [0:0] notOp_366_in0;
	wire [0:0] notOp_366_out;
	notOp #(.WIDTH(1)) notOp_366(.in(notOp_366_in0), .out(notOp_366_out));

	reg [0:0] andOp_367_in0;
	reg [0:0] andOp_367_in1;
	wire [0:0] andOp_367_out;
	andOp #(.WIDTH(1)) andOp_367(.in0(andOp_367_in0), .in1(andOp_367_in1), .out(andOp_367_out));

	reg [0:0] andOp_368_in0;
	reg [0:0] andOp_368_in1;
	wire [0:0] andOp_368_out;
	andOp #(.WIDTH(1)) andOp_368(.in0(andOp_368_in0), .in1(andOp_368_in1), .out(andOp_368_out));

	reg [31:0] eq_369_in0;
	reg [31:0] eq_369_in1;
	wire [0:0] eq_369_out;
	eq #(.WIDTH(32)) eq_369(.in0(eq_369_in0), .in1(eq_369_in1), .out(eq_369_out));

	reg [0:0] andOp_370_in0;
	reg [0:0] andOp_370_in1;
	wire [0:0] andOp_370_out;
	andOp #(.WIDTH(1)) andOp_370(.in0(andOp_370_in0), .in1(andOp_370_in1), .out(andOp_370_out));

	reg [0:0] notOp_371_in0;
	wire [0:0] notOp_371_out;
	notOp #(.WIDTH(1)) notOp_371(.in(notOp_371_in0), .out(notOp_371_out));

	reg [0:0] andOp_372_in0;
	reg [0:0] andOp_372_in1;
	wire [0:0] andOp_372_out;
	andOp #(.WIDTH(1)) andOp_372(.in0(andOp_372_in0), .in1(andOp_372_in1), .out(andOp_372_out));

	reg [0:0] andOp_373_in0;
	reg [0:0] andOp_373_in1;
	wire [0:0] andOp_373_out;
	andOp #(.WIDTH(1)) andOp_373(.in0(andOp_373_in0), .in1(andOp_373_in1), .out(andOp_373_out));

	reg [31:0] eq_374_in0;
	reg [31:0] eq_374_in1;
	wire [0:0] eq_374_out;
	eq #(.WIDTH(32)) eq_374(.in0(eq_374_in0), .in1(eq_374_in1), .out(eq_374_out));

	reg [0:0] andOp_375_in0;
	reg [0:0] andOp_375_in1;
	wire [0:0] andOp_375_out;
	andOp #(.WIDTH(1)) andOp_375(.in0(andOp_375_in0), .in1(andOp_375_in1), .out(andOp_375_out));

	reg [0:0] notOp_376_in0;
	wire [0:0] notOp_376_out;
	notOp #(.WIDTH(1)) notOp_376(.in(notOp_376_in0), .out(notOp_376_out));

	reg [0:0] andOp_377_in0;
	reg [0:0] andOp_377_in1;
	wire [0:0] andOp_377_out;
	andOp #(.WIDTH(1)) andOp_377(.in0(andOp_377_in0), .in1(andOp_377_in1), .out(andOp_377_out));

	reg [0:0] andOp_378_in0;
	reg [0:0] andOp_378_in1;
	wire [0:0] andOp_378_out;
	andOp #(.WIDTH(1)) andOp_378(.in0(andOp_378_in0), .in1(andOp_378_in1), .out(andOp_378_out));

	reg [31:0] eq_379_in0;
	reg [31:0] eq_379_in1;
	wire [0:0] eq_379_out;
	eq #(.WIDTH(32)) eq_379(.in0(eq_379_in0), .in1(eq_379_in1), .out(eq_379_out));

	reg [0:0] andOp_380_in0;
	reg [0:0] andOp_380_in1;
	wire [0:0] andOp_380_out;
	andOp #(.WIDTH(1)) andOp_380(.in0(andOp_380_in0), .in1(andOp_380_in1), .out(andOp_380_out));

	reg [0:0] notOp_381_in0;
	wire [0:0] notOp_381_out;
	notOp #(.WIDTH(1)) notOp_381(.in(notOp_381_in0), .out(notOp_381_out));

	reg [0:0] andOp_382_in0;
	reg [0:0] andOp_382_in1;
	wire [0:0] andOp_382_out;
	andOp #(.WIDTH(1)) andOp_382(.in0(andOp_382_in0), .in1(andOp_382_in1), .out(andOp_382_out));

	reg [0:0] andOp_383_in0;
	reg [0:0] andOp_383_in1;
	wire [0:0] andOp_383_out;
	andOp #(.WIDTH(1)) andOp_383(.in0(andOp_383_in0), .in1(andOp_383_in1), .out(andOp_383_out));

	reg [31:0] eq_384_in0;
	reg [31:0] eq_384_in1;
	wire [0:0] eq_384_out;
	eq #(.WIDTH(32)) eq_384(.in0(eq_384_in0), .in1(eq_384_in1), .out(eq_384_out));

	reg [0:0] andOp_385_in0;
	reg [0:0] andOp_385_in1;
	wire [0:0] andOp_385_out;
	andOp #(.WIDTH(1)) andOp_385(.in0(andOp_385_in0), .in1(andOp_385_in1), .out(andOp_385_out));

	reg [0:0] notOp_386_in0;
	wire [0:0] notOp_386_out;
	notOp #(.WIDTH(1)) notOp_386(.in(notOp_386_in0), .out(notOp_386_out));

	reg [0:0] andOp_387_in0;
	reg [0:0] andOp_387_in1;
	wire [0:0] andOp_387_out;
	andOp #(.WIDTH(1)) andOp_387(.in0(andOp_387_in0), .in1(andOp_387_in1), .out(andOp_387_out));

	reg [0:0] andOp_388_in0;
	reg [0:0] andOp_388_in1;
	wire [0:0] andOp_388_out;
	andOp #(.WIDTH(1)) andOp_388(.in0(andOp_388_in0), .in1(andOp_388_in1), .out(andOp_388_out));

	reg [31:0] eq_389_in0;
	reg [31:0] eq_389_in1;
	wire [0:0] eq_389_out;
	eq #(.WIDTH(32)) eq_389(.in0(eq_389_in0), .in1(eq_389_in1), .out(eq_389_out));

	reg [0:0] andOp_390_in0;
	reg [0:0] andOp_390_in1;
	wire [0:0] andOp_390_out;
	andOp #(.WIDTH(1)) andOp_390(.in0(andOp_390_in0), .in1(andOp_390_in1), .out(andOp_390_out));

	reg [0:0] notOp_391_in0;
	wire [0:0] notOp_391_out;
	notOp #(.WIDTH(1)) notOp_391(.in(notOp_391_in0), .out(notOp_391_out));

	reg [0:0] andOp_392_in0;
	reg [0:0] andOp_392_in1;
	wire [0:0] andOp_392_out;
	andOp #(.WIDTH(1)) andOp_392(.in0(andOp_392_in0), .in1(andOp_392_in1), .out(andOp_392_out));

	reg [0:0] andOp_393_in0;
	reg [0:0] andOp_393_in1;
	wire [0:0] andOp_393_out;
	andOp #(.WIDTH(1)) andOp_393(.in0(andOp_393_in0), .in1(andOp_393_in1), .out(andOp_393_out));

	reg [31:0] eq_394_in0;
	reg [31:0] eq_394_in1;
	wire [0:0] eq_394_out;
	eq #(.WIDTH(32)) eq_394(.in0(eq_394_in0), .in1(eq_394_in1), .out(eq_394_out));

	reg [0:0] andOp_395_in0;
	reg [0:0] andOp_395_in1;
	wire [0:0] andOp_395_out;
	andOp #(.WIDTH(1)) andOp_395(.in0(andOp_395_in0), .in1(andOp_395_in1), .out(andOp_395_out));

	reg [0:0] notOp_396_in0;
	wire [0:0] notOp_396_out;
	notOp #(.WIDTH(1)) notOp_396(.in(notOp_396_in0), .out(notOp_396_out));

	reg [0:0] andOp_397_in0;
	reg [0:0] andOp_397_in1;
	wire [0:0] andOp_397_out;
	andOp #(.WIDTH(1)) andOp_397(.in0(andOp_397_in0), .in1(andOp_397_in1), .out(andOp_397_out));

	reg [0:0] andOp_398_in0;
	reg [0:0] andOp_398_in1;
	wire [0:0] andOp_398_out;
	andOp #(.WIDTH(1)) andOp_398(.in0(andOp_398_in0), .in1(andOp_398_in1), .out(andOp_398_out));

	reg [31:0] eq_399_in0;
	reg [31:0] eq_399_in1;
	wire [0:0] eq_399_out;
	eq #(.WIDTH(32)) eq_399(.in0(eq_399_in0), .in1(eq_399_in1), .out(eq_399_out));

	reg [0:0] andOp_400_in0;
	reg [0:0] andOp_400_in1;
	wire [0:0] andOp_400_out;
	andOp #(.WIDTH(1)) andOp_400(.in0(andOp_400_in0), .in1(andOp_400_in1), .out(andOp_400_out));

	reg [0:0] notOp_401_in0;
	wire [0:0] notOp_401_out;
	notOp #(.WIDTH(1)) notOp_401(.in(notOp_401_in0), .out(notOp_401_out));

	reg [0:0] andOp_402_in0;
	reg [0:0] andOp_402_in1;
	wire [0:0] andOp_402_out;
	andOp #(.WIDTH(1)) andOp_402(.in0(andOp_402_in0), .in1(andOp_402_in1), .out(andOp_402_out));

	reg [0:0] andOp_403_in0;
	reg [0:0] andOp_403_in1;
	wire [0:0] andOp_403_out;
	andOp #(.WIDTH(1)) andOp_403(.in0(andOp_403_in0), .in1(andOp_403_in1), .out(andOp_403_out));

	reg [31:0] eq_404_in0;
	reg [31:0] eq_404_in1;
	wire [0:0] eq_404_out;
	eq #(.WIDTH(32)) eq_404(.in0(eq_404_in0), .in1(eq_404_in1), .out(eq_404_out));

	reg [0:0] andOp_405_in0;
	reg [0:0] andOp_405_in1;
	wire [0:0] andOp_405_out;
	andOp #(.WIDTH(1)) andOp_405(.in0(andOp_405_in0), .in1(andOp_405_in1), .out(andOp_405_out));

	reg [0:0] notOp_406_in0;
	wire [0:0] notOp_406_out;
	notOp #(.WIDTH(1)) notOp_406(.in(notOp_406_in0), .out(notOp_406_out));

	reg [0:0] andOp_407_in0;
	reg [0:0] andOp_407_in1;
	wire [0:0] andOp_407_out;
	andOp #(.WIDTH(1)) andOp_407(.in0(andOp_407_in0), .in1(andOp_407_in1), .out(andOp_407_out));

	reg [31:0] eq_408_in0;
	reg [31:0] eq_408_in1;
	wire [0:0] eq_408_out;
	eq #(.WIDTH(32)) eq_408(.in0(eq_408_in0), .in1(eq_408_in1), .out(eq_408_out));

	reg [0:0] andOp_409_in0;
	reg [0:0] andOp_409_in1;
	wire [0:0] andOp_409_out;
	andOp #(.WIDTH(1)) andOp_409(.in0(andOp_409_in0), .in1(andOp_409_in1), .out(andOp_409_out));

	reg [31:0] eq_410_in0;
	reg [31:0] eq_410_in1;
	wire [0:0] eq_410_out;
	eq #(.WIDTH(32)) eq_410(.in0(eq_410_in0), .in1(eq_410_in1), .out(eq_410_out));

	reg [0:0] andOp_411_in0;
	reg [0:0] andOp_411_in1;
	wire [0:0] andOp_411_out;
	andOp #(.WIDTH(1)) andOp_411(.in0(andOp_411_in0), .in1(andOp_411_in1), .out(andOp_411_out));

	reg [31:0] eq_412_in0;
	reg [31:0] eq_412_in1;
	wire [0:0] eq_412_out;
	eq #(.WIDTH(32)) eq_412(.in0(eq_412_in0), .in1(eq_412_in1), .out(eq_412_out));

	reg [0:0] andOp_413_in0;
	reg [0:0] andOp_413_in1;
	wire [0:0] andOp_413_out;
	andOp #(.WIDTH(1)) andOp_413(.in0(andOp_413_in0), .in1(andOp_413_in1), .out(andOp_413_out));

	reg [31:0] eq_414_in0;
	reg [31:0] eq_414_in1;
	wire [0:0] eq_414_out;
	eq #(.WIDTH(32)) eq_414(.in0(eq_414_in0), .in1(eq_414_in1), .out(eq_414_out));

	reg [0:0] andOp_415_in0;
	reg [0:0] andOp_415_in1;
	wire [0:0] andOp_415_out;
	andOp #(.WIDTH(1)) andOp_415(.in0(andOp_415_in0), .in1(andOp_415_in1), .out(andOp_415_out));

	reg [31:0] eq_416_in0;
	reg [31:0] eq_416_in1;
	wire [0:0] eq_416_out;
	eq #(.WIDTH(32)) eq_416(.in0(eq_416_in0), .in1(eq_416_in1), .out(eq_416_out));

	reg [0:0] andOp_417_in0;
	reg [0:0] andOp_417_in1;
	wire [0:0] andOp_417_out;
	andOp #(.WIDTH(1)) andOp_417(.in0(andOp_417_in0), .in1(andOp_417_in1), .out(andOp_417_out));

	reg [0:0] andOp_418_in0;
	reg [0:0] andOp_418_in1;
	wire [0:0] andOp_418_out;
	andOp #(.WIDTH(1)) andOp_418(.in0(andOp_418_in0), .in1(andOp_418_in1), .out(andOp_418_out));

	reg [31:0] eq_419_in0;
	reg [31:0] eq_419_in1;
	wire [0:0] eq_419_out;
	eq #(.WIDTH(32)) eq_419(.in0(eq_419_in0), .in1(eq_419_in1), .out(eq_419_out));

	reg [0:0] andOp_420_in0;
	reg [0:0] andOp_420_in1;
	wire [0:0] andOp_420_out;
	andOp #(.WIDTH(1)) andOp_420(.in0(andOp_420_in0), .in1(andOp_420_in1), .out(andOp_420_out));

	reg [0:0] notOp_421_in0;
	wire [0:0] notOp_421_out;
	notOp #(.WIDTH(1)) notOp_421(.in(notOp_421_in0), .out(notOp_421_out));

	reg [0:0] andOp_422_in0;
	reg [0:0] andOp_422_in1;
	wire [0:0] andOp_422_out;
	andOp #(.WIDTH(1)) andOp_422(.in0(andOp_422_in0), .in1(andOp_422_in1), .out(andOp_422_out));

	reg [0:0] andOp_423_in0;
	reg [0:0] andOp_423_in1;
	wire [0:0] andOp_423_out;
	andOp #(.WIDTH(1)) andOp_423(.in0(andOp_423_in0), .in1(andOp_423_in1), .out(andOp_423_out));

	reg [31:0] eq_424_in0;
	reg [31:0] eq_424_in1;
	wire [0:0] eq_424_out;
	eq #(.WIDTH(32)) eq_424(.in0(eq_424_in0), .in1(eq_424_in1), .out(eq_424_out));

	reg [0:0] andOp_425_in0;
	reg [0:0] andOp_425_in1;
	wire [0:0] andOp_425_out;
	andOp #(.WIDTH(1)) andOp_425(.in0(andOp_425_in0), .in1(andOp_425_in1), .out(andOp_425_out));

	reg [0:0] notOp_426_in0;
	wire [0:0] notOp_426_out;
	notOp #(.WIDTH(1)) notOp_426(.in(notOp_426_in0), .out(notOp_426_out));

	reg [0:0] andOp_427_in0;
	reg [0:0] andOp_427_in1;
	wire [0:0] andOp_427_out;
	andOp #(.WIDTH(1)) andOp_427(.in0(andOp_427_in0), .in1(andOp_427_in1), .out(andOp_427_out));

	reg [0:0] andOp_428_in0;
	reg [0:0] andOp_428_in1;
	wire [0:0] andOp_428_out;
	andOp #(.WIDTH(1)) andOp_428(.in0(andOp_428_in0), .in1(andOp_428_in1), .out(andOp_428_out));

	reg [31:0] eq_429_in0;
	reg [31:0] eq_429_in1;
	wire [0:0] eq_429_out;
	eq #(.WIDTH(32)) eq_429(.in0(eq_429_in0), .in1(eq_429_in1), .out(eq_429_out));

	reg [0:0] andOp_430_in0;
	reg [0:0] andOp_430_in1;
	wire [0:0] andOp_430_out;
	andOp #(.WIDTH(1)) andOp_430(.in0(andOp_430_in0), .in1(andOp_430_in1), .out(andOp_430_out));

	reg [0:0] notOp_431_in0;
	wire [0:0] notOp_431_out;
	notOp #(.WIDTH(1)) notOp_431(.in(notOp_431_in0), .out(notOp_431_out));

	reg [0:0] andOp_432_in0;
	reg [0:0] andOp_432_in1;
	wire [0:0] andOp_432_out;
	andOp #(.WIDTH(1)) andOp_432(.in0(andOp_432_in0), .in1(andOp_432_in1), .out(andOp_432_out));

	reg [0:0] andOp_433_in0;
	reg [0:0] andOp_433_in1;
	wire [0:0] andOp_433_out;
	andOp #(.WIDTH(1)) andOp_433(.in0(andOp_433_in0), .in1(andOp_433_in1), .out(andOp_433_out));

	reg [31:0] eq_434_in0;
	reg [31:0] eq_434_in1;
	wire [0:0] eq_434_out;
	eq #(.WIDTH(32)) eq_434(.in0(eq_434_in0), .in1(eq_434_in1), .out(eq_434_out));

	reg [0:0] andOp_435_in0;
	reg [0:0] andOp_435_in1;
	wire [0:0] andOp_435_out;
	andOp #(.WIDTH(1)) andOp_435(.in0(andOp_435_in0), .in1(andOp_435_in1), .out(andOp_435_out));

	reg [0:0] notOp_436_in0;
	wire [0:0] notOp_436_out;
	notOp #(.WIDTH(1)) notOp_436(.in(notOp_436_in0), .out(notOp_436_out));

	reg [0:0] andOp_437_in0;
	reg [0:0] andOp_437_in1;
	wire [0:0] andOp_437_out;
	andOp #(.WIDTH(1)) andOp_437(.in0(andOp_437_in0), .in1(andOp_437_in1), .out(andOp_437_out));

	reg [0:0] andOp_438_in0;
	reg [0:0] andOp_438_in1;
	wire [0:0] andOp_438_out;
	andOp #(.WIDTH(1)) andOp_438(.in0(andOp_438_in0), .in1(andOp_438_in1), .out(andOp_438_out));

	reg [31:0] eq_439_in0;
	reg [31:0] eq_439_in1;
	wire [0:0] eq_439_out;
	eq #(.WIDTH(32)) eq_439(.in0(eq_439_in0), .in1(eq_439_in1), .out(eq_439_out));

	reg [0:0] andOp_440_in0;
	reg [0:0] andOp_440_in1;
	wire [0:0] andOp_440_out;
	andOp #(.WIDTH(1)) andOp_440(.in0(andOp_440_in0), .in1(andOp_440_in1), .out(andOp_440_out));

	reg [0:0] notOp_441_in0;
	wire [0:0] notOp_441_out;
	notOp #(.WIDTH(1)) notOp_441(.in(notOp_441_in0), .out(notOp_441_out));

	reg [0:0] andOp_442_in0;
	reg [0:0] andOp_442_in1;
	wire [0:0] andOp_442_out;
	andOp #(.WIDTH(1)) andOp_442(.in0(andOp_442_in0), .in1(andOp_442_in1), .out(andOp_442_out));

	reg [0:0] andOp_443_in0;
	reg [0:0] andOp_443_in1;
	wire [0:0] andOp_443_out;
	andOp #(.WIDTH(1)) andOp_443(.in0(andOp_443_in0), .in1(andOp_443_in1), .out(andOp_443_out));

	reg [31:0] eq_444_in0;
	reg [31:0] eq_444_in1;
	wire [0:0] eq_444_out;
	eq #(.WIDTH(32)) eq_444(.in0(eq_444_in0), .in1(eq_444_in1), .out(eq_444_out));

	reg [0:0] andOp_445_in0;
	reg [0:0] andOp_445_in1;
	wire [0:0] andOp_445_out;
	andOp #(.WIDTH(1)) andOp_445(.in0(andOp_445_in0), .in1(andOp_445_in1), .out(andOp_445_out));

	reg [0:0] notOp_446_in0;
	wire [0:0] notOp_446_out;
	notOp #(.WIDTH(1)) notOp_446(.in(notOp_446_in0), .out(notOp_446_out));

	reg [0:0] andOp_447_in0;
	reg [0:0] andOp_447_in1;
	wire [0:0] andOp_447_out;
	andOp #(.WIDTH(1)) andOp_447(.in0(andOp_447_in0), .in1(andOp_447_in1), .out(andOp_447_out));

	reg [0:0] andOp_448_in0;
	reg [0:0] andOp_448_in1;
	wire [0:0] andOp_448_out;
	andOp #(.WIDTH(1)) andOp_448(.in0(andOp_448_in0), .in1(andOp_448_in1), .out(andOp_448_out));

	reg [31:0] eq_449_in0;
	reg [31:0] eq_449_in1;
	wire [0:0] eq_449_out;
	eq #(.WIDTH(32)) eq_449(.in0(eq_449_in0), .in1(eq_449_in1), .out(eq_449_out));

	reg [0:0] andOp_450_in0;
	reg [0:0] andOp_450_in1;
	wire [0:0] andOp_450_out;
	andOp #(.WIDTH(1)) andOp_450(.in0(andOp_450_in0), .in1(andOp_450_in1), .out(andOp_450_out));

	reg [0:0] notOp_451_in0;
	wire [0:0] notOp_451_out;
	notOp #(.WIDTH(1)) notOp_451(.in(notOp_451_in0), .out(notOp_451_out));

	reg [0:0] andOp_452_in0;
	reg [0:0] andOp_452_in1;
	wire [0:0] andOp_452_out;
	andOp #(.WIDTH(1)) andOp_452(.in0(andOp_452_in0), .in1(andOp_452_in1), .out(andOp_452_out));

	reg [0:0] andOp_453_in0;
	reg [0:0] andOp_453_in1;
	wire [0:0] andOp_453_out;
	andOp #(.WIDTH(1)) andOp_453(.in0(andOp_453_in0), .in1(andOp_453_in1), .out(andOp_453_out));

	reg [31:0] eq_454_in0;
	reg [31:0] eq_454_in1;
	wire [0:0] eq_454_out;
	eq #(.WIDTH(32)) eq_454(.in0(eq_454_in0), .in1(eq_454_in1), .out(eq_454_out));

	reg [0:0] andOp_455_in0;
	reg [0:0] andOp_455_in1;
	wire [0:0] andOp_455_out;
	andOp #(.WIDTH(1)) andOp_455(.in0(andOp_455_in0), .in1(andOp_455_in1), .out(andOp_455_out));

	reg [0:0] notOp_456_in0;
	wire [0:0] notOp_456_out;
	notOp #(.WIDTH(1)) notOp_456(.in(notOp_456_in0), .out(notOp_456_out));

	reg [0:0] andOp_457_in0;
	reg [0:0] andOp_457_in1;
	wire [0:0] andOp_457_out;
	andOp #(.WIDTH(1)) andOp_457(.in0(andOp_457_in0), .in1(andOp_457_in1), .out(andOp_457_out));

	reg [0:0] andOp_458_in0;
	reg [0:0] andOp_458_in1;
	wire [0:0] andOp_458_out;
	andOp #(.WIDTH(1)) andOp_458(.in0(andOp_458_in0), .in1(andOp_458_in1), .out(andOp_458_out));

	reg [31:0] eq_459_in0;
	reg [31:0] eq_459_in1;
	wire [0:0] eq_459_out;
	eq #(.WIDTH(32)) eq_459(.in0(eq_459_in0), .in1(eq_459_in1), .out(eq_459_out));

	reg [0:0] andOp_460_in0;
	reg [0:0] andOp_460_in1;
	wire [0:0] andOp_460_out;
	andOp #(.WIDTH(1)) andOp_460(.in0(andOp_460_in0), .in1(andOp_460_in1), .out(andOp_460_out));

	reg [0:0] notOp_461_in0;
	wire [0:0] notOp_461_out;
	notOp #(.WIDTH(1)) notOp_461(.in(notOp_461_in0), .out(notOp_461_out));

	reg [0:0] andOp_462_in0;
	reg [0:0] andOp_462_in1;
	wire [0:0] andOp_462_out;
	andOp #(.WIDTH(1)) andOp_462(.in0(andOp_462_in0), .in1(andOp_462_in1), .out(andOp_462_out));

	reg [31:0] eq_463_in0;
	reg [31:0] eq_463_in1;
	wire [0:0] eq_463_out;
	eq #(.WIDTH(32)) eq_463(.in0(eq_463_in0), .in1(eq_463_in1), .out(eq_463_out));

	reg [0:0] andOp_464_in0;
	reg [0:0] andOp_464_in1;
	wire [0:0] andOp_464_out;
	andOp #(.WIDTH(1)) andOp_464(.in0(andOp_464_in0), .in1(andOp_464_in1), .out(andOp_464_out));

	reg [31:0] eq_465_in0;
	reg [31:0] eq_465_in1;
	wire [0:0] eq_465_out;
	eq #(.WIDTH(32)) eq_465(.in0(eq_465_in0), .in1(eq_465_in1), .out(eq_465_out));

	reg [0:0] andOp_466_in0;
	reg [0:0] andOp_466_in1;
	wire [0:0] andOp_466_out;
	andOp #(.WIDTH(1)) andOp_466(.in0(andOp_466_in0), .in1(andOp_466_in1), .out(andOp_466_out));

	reg [31:0] eq_467_in0;
	reg [31:0] eq_467_in1;
	wire [0:0] eq_467_out;
	eq #(.WIDTH(32)) eq_467(.in0(eq_467_in0), .in1(eq_467_in1), .out(eq_467_out));

	reg [0:0] andOp_468_in0;
	reg [0:0] andOp_468_in1;
	wire [0:0] andOp_468_out;
	andOp #(.WIDTH(1)) andOp_468(.in0(andOp_468_in0), .in1(andOp_468_in1), .out(andOp_468_out));

	reg [31:0] eq_469_in0;
	reg [31:0] eq_469_in1;
	wire [0:0] eq_469_out;
	eq #(.WIDTH(32)) eq_469(.in0(eq_469_in0), .in1(eq_469_in1), .out(eq_469_out));

	reg [0:0] andOp_470_in0;
	reg [0:0] andOp_470_in1;
	wire [0:0] andOp_470_out;
	andOp #(.WIDTH(1)) andOp_470(.in0(andOp_470_in0), .in1(andOp_470_in1), .out(andOp_470_out));

	reg [31:0] eq_471_in0;
	reg [31:0] eq_471_in1;
	wire [0:0] eq_471_out;
	eq #(.WIDTH(32)) eq_471(.in0(eq_471_in0), .in1(eq_471_in1), .out(eq_471_out));

	reg [0:0] andOp_472_in0;
	reg [0:0] andOp_472_in1;
	wire [0:0] andOp_472_out;
	andOp #(.WIDTH(1)) andOp_472(.in0(andOp_472_in0), .in1(andOp_472_in1), .out(andOp_472_out));

	reg [0:0] andOp_473_in0;
	reg [0:0] andOp_473_in1;
	wire [0:0] andOp_473_out;
	andOp #(.WIDTH(1)) andOp_473(.in0(andOp_473_in0), .in1(andOp_473_in1), .out(andOp_473_out));

	reg [31:0] eq_474_in0;
	reg [31:0] eq_474_in1;
	wire [0:0] eq_474_out;
	eq #(.WIDTH(32)) eq_474(.in0(eq_474_in0), .in1(eq_474_in1), .out(eq_474_out));

	reg [0:0] andOp_475_in0;
	reg [0:0] andOp_475_in1;
	wire [0:0] andOp_475_out;
	andOp #(.WIDTH(1)) andOp_475(.in0(andOp_475_in0), .in1(andOp_475_in1), .out(andOp_475_out));

	reg [0:0] notOp_476_in0;
	wire [0:0] notOp_476_out;
	notOp #(.WIDTH(1)) notOp_476(.in(notOp_476_in0), .out(notOp_476_out));

	reg [0:0] andOp_477_in0;
	reg [0:0] andOp_477_in1;
	wire [0:0] andOp_477_out;
	andOp #(.WIDTH(1)) andOp_477(.in0(andOp_477_in0), .in1(andOp_477_in1), .out(andOp_477_out));

	reg [0:0] andOp_478_in0;
	reg [0:0] andOp_478_in1;
	wire [0:0] andOp_478_out;
	andOp #(.WIDTH(1)) andOp_478(.in0(andOp_478_in0), .in1(andOp_478_in1), .out(andOp_478_out));

	reg [31:0] eq_479_in0;
	reg [31:0] eq_479_in1;
	wire [0:0] eq_479_out;
	eq #(.WIDTH(32)) eq_479(.in0(eq_479_in0), .in1(eq_479_in1), .out(eq_479_out));

	reg [0:0] andOp_480_in0;
	reg [0:0] andOp_480_in1;
	wire [0:0] andOp_480_out;
	andOp #(.WIDTH(1)) andOp_480(.in0(andOp_480_in0), .in1(andOp_480_in1), .out(andOp_480_out));

	reg [0:0] notOp_481_in0;
	wire [0:0] notOp_481_out;
	notOp #(.WIDTH(1)) notOp_481(.in(notOp_481_in0), .out(notOp_481_out));

	reg [0:0] andOp_482_in0;
	reg [0:0] andOp_482_in1;
	wire [0:0] andOp_482_out;
	andOp #(.WIDTH(1)) andOp_482(.in0(andOp_482_in0), .in1(andOp_482_in1), .out(andOp_482_out));

	reg [0:0] andOp_483_in0;
	reg [0:0] andOp_483_in1;
	wire [0:0] andOp_483_out;
	andOp #(.WIDTH(1)) andOp_483(.in0(andOp_483_in0), .in1(andOp_483_in1), .out(andOp_483_out));

	reg [31:0] eq_484_in0;
	reg [31:0] eq_484_in1;
	wire [0:0] eq_484_out;
	eq #(.WIDTH(32)) eq_484(.in0(eq_484_in0), .in1(eq_484_in1), .out(eq_484_out));

	reg [0:0] andOp_485_in0;
	reg [0:0] andOp_485_in1;
	wire [0:0] andOp_485_out;
	andOp #(.WIDTH(1)) andOp_485(.in0(andOp_485_in0), .in1(andOp_485_in1), .out(andOp_485_out));

	reg [0:0] notOp_486_in0;
	wire [0:0] notOp_486_out;
	notOp #(.WIDTH(1)) notOp_486(.in(notOp_486_in0), .out(notOp_486_out));

	reg [0:0] andOp_487_in0;
	reg [0:0] andOp_487_in1;
	wire [0:0] andOp_487_out;
	andOp #(.WIDTH(1)) andOp_487(.in0(andOp_487_in0), .in1(andOp_487_in1), .out(andOp_487_out));

	reg [0:0] andOp_488_in0;
	reg [0:0] andOp_488_in1;
	wire [0:0] andOp_488_out;
	andOp #(.WIDTH(1)) andOp_488(.in0(andOp_488_in0), .in1(andOp_488_in1), .out(andOp_488_out));

	reg [31:0] eq_489_in0;
	reg [31:0] eq_489_in1;
	wire [0:0] eq_489_out;
	eq #(.WIDTH(32)) eq_489(.in0(eq_489_in0), .in1(eq_489_in1), .out(eq_489_out));

	reg [0:0] andOp_490_in0;
	reg [0:0] andOp_490_in1;
	wire [0:0] andOp_490_out;
	andOp #(.WIDTH(1)) andOp_490(.in0(andOp_490_in0), .in1(andOp_490_in1), .out(andOp_490_out));

	reg [0:0] notOp_491_in0;
	wire [0:0] notOp_491_out;
	notOp #(.WIDTH(1)) notOp_491(.in(notOp_491_in0), .out(notOp_491_out));

	reg [0:0] andOp_492_in0;
	reg [0:0] andOp_492_in1;
	wire [0:0] andOp_492_out;
	andOp #(.WIDTH(1)) andOp_492(.in0(andOp_492_in0), .in1(andOp_492_in1), .out(andOp_492_out));

	reg [0:0] andOp_493_in0;
	reg [0:0] andOp_493_in1;
	wire [0:0] andOp_493_out;
	andOp #(.WIDTH(1)) andOp_493(.in0(andOp_493_in0), .in1(andOp_493_in1), .out(andOp_493_out));

	reg [31:0] eq_494_in0;
	reg [31:0] eq_494_in1;
	wire [0:0] eq_494_out;
	eq #(.WIDTH(32)) eq_494(.in0(eq_494_in0), .in1(eq_494_in1), .out(eq_494_out));

	reg [0:0] andOp_495_in0;
	reg [0:0] andOp_495_in1;
	wire [0:0] andOp_495_out;
	andOp #(.WIDTH(1)) andOp_495(.in0(andOp_495_in0), .in1(andOp_495_in1), .out(andOp_495_out));

	reg [0:0] notOp_496_in0;
	wire [0:0] notOp_496_out;
	notOp #(.WIDTH(1)) notOp_496(.in(notOp_496_in0), .out(notOp_496_out));

	reg [0:0] andOp_497_in0;
	reg [0:0] andOp_497_in1;
	wire [0:0] andOp_497_out;
	andOp #(.WIDTH(1)) andOp_497(.in0(andOp_497_in0), .in1(andOp_497_in1), .out(andOp_497_out));

	reg [0:0] andOp_498_in0;
	reg [0:0] andOp_498_in1;
	wire [0:0] andOp_498_out;
	andOp #(.WIDTH(1)) andOp_498(.in0(andOp_498_in0), .in1(andOp_498_in1), .out(andOp_498_out));

	reg [31:0] eq_499_in0;
	reg [31:0] eq_499_in1;
	wire [0:0] eq_499_out;
	eq #(.WIDTH(32)) eq_499(.in0(eq_499_in0), .in1(eq_499_in1), .out(eq_499_out));

	reg [0:0] andOp_500_in0;
	reg [0:0] andOp_500_in1;
	wire [0:0] andOp_500_out;
	andOp #(.WIDTH(1)) andOp_500(.in0(andOp_500_in0), .in1(andOp_500_in1), .out(andOp_500_out));

	reg [0:0] notOp_501_in0;
	wire [0:0] notOp_501_out;
	notOp #(.WIDTH(1)) notOp_501(.in(notOp_501_in0), .out(notOp_501_out));

	reg [0:0] andOp_502_in0;
	reg [0:0] andOp_502_in1;
	wire [0:0] andOp_502_out;
	andOp #(.WIDTH(1)) andOp_502(.in0(andOp_502_in0), .in1(andOp_502_in1), .out(andOp_502_out));

	reg [0:0] andOp_503_in0;
	reg [0:0] andOp_503_in1;
	wire [0:0] andOp_503_out;
	andOp #(.WIDTH(1)) andOp_503(.in0(andOp_503_in0), .in1(andOp_503_in1), .out(andOp_503_out));

	reg [31:0] eq_504_in0;
	reg [31:0] eq_504_in1;
	wire [0:0] eq_504_out;
	eq #(.WIDTH(32)) eq_504(.in0(eq_504_in0), .in1(eq_504_in1), .out(eq_504_out));

	reg [0:0] andOp_505_in0;
	reg [0:0] andOp_505_in1;
	wire [0:0] andOp_505_out;
	andOp #(.WIDTH(1)) andOp_505(.in0(andOp_505_in0), .in1(andOp_505_in1), .out(andOp_505_out));

	reg [0:0] notOp_506_in0;
	wire [0:0] notOp_506_out;
	notOp #(.WIDTH(1)) notOp_506(.in(notOp_506_in0), .out(notOp_506_out));

	reg [0:0] andOp_507_in0;
	reg [0:0] andOp_507_in1;
	wire [0:0] andOp_507_out;
	andOp #(.WIDTH(1)) andOp_507(.in0(andOp_507_in0), .in1(andOp_507_in1), .out(andOp_507_out));

	reg [0:0] andOp_508_in0;
	reg [0:0] andOp_508_in1;
	wire [0:0] andOp_508_out;
	andOp #(.WIDTH(1)) andOp_508(.in0(andOp_508_in0), .in1(andOp_508_in1), .out(andOp_508_out));

	reg [31:0] eq_509_in0;
	reg [31:0] eq_509_in1;
	wire [0:0] eq_509_out;
	eq #(.WIDTH(32)) eq_509(.in0(eq_509_in0), .in1(eq_509_in1), .out(eq_509_out));

	reg [0:0] andOp_510_in0;
	reg [0:0] andOp_510_in1;
	wire [0:0] andOp_510_out;
	andOp #(.WIDTH(1)) andOp_510(.in0(andOp_510_in0), .in1(andOp_510_in1), .out(andOp_510_out));

	reg [0:0] notOp_511_in0;
	wire [0:0] notOp_511_out;
	notOp #(.WIDTH(1)) notOp_511(.in(notOp_511_in0), .out(notOp_511_out));

	reg [0:0] andOp_512_in0;
	reg [0:0] andOp_512_in1;
	wire [0:0] andOp_512_out;
	andOp #(.WIDTH(1)) andOp_512(.in0(andOp_512_in0), .in1(andOp_512_in1), .out(andOp_512_out));

	reg [0:0] andOp_513_in0;
	reg [0:0] andOp_513_in1;
	wire [0:0] andOp_513_out;
	andOp #(.WIDTH(1)) andOp_513(.in0(andOp_513_in0), .in1(andOp_513_in1), .out(andOp_513_out));

	reg [31:0] eq_514_in0;
	reg [31:0] eq_514_in1;
	wire [0:0] eq_514_out;
	eq #(.WIDTH(32)) eq_514(.in0(eq_514_in0), .in1(eq_514_in1), .out(eq_514_out));

	reg [0:0] andOp_515_in0;
	reg [0:0] andOp_515_in1;
	wire [0:0] andOp_515_out;
	andOp #(.WIDTH(1)) andOp_515(.in0(andOp_515_in0), .in1(andOp_515_in1), .out(andOp_515_out));

	reg [0:0] notOp_516_in0;
	wire [0:0] notOp_516_out;
	notOp #(.WIDTH(1)) notOp_516(.in(notOp_516_in0), .out(notOp_516_out));

	reg [0:0] andOp_517_in0;
	reg [0:0] andOp_517_in1;
	wire [0:0] andOp_517_out;
	andOp #(.WIDTH(1)) andOp_517(.in0(andOp_517_in0), .in1(andOp_517_in1), .out(andOp_517_out));

	// End Functional Units

	reg [31:0] add_tmp_4;
	reg [31:0] call_tmp_6;
	reg [31:0] data_store_0_0;
	reg [0:0] data_store_0_10;
	reg [31:0] data_store_0_12;
	reg [0:0] data_store_0_14;
	reg [31:0] data_store_0_16;
	reg [31:0] data_store_0_2;
	reg [31:0] data_store_0_4;
	reg [31:0] data_store_0_6;
	reg [0:0] data_store_0_8;
	reg [31:0] data_store_1_18;
	reg [31:0] data_store_1_20;
	reg [31:0] data_store_1_22;
	reg [31:0] data_store_1_24;
	reg [0:0] data_store_1_26;
	reg [0:0] data_store_1_28;
	reg [31:0] data_store_1_30;
	reg [0:0] data_store_1_32;
	reg [31:0] data_store_1_34;
	reg [31:0] data_store_2_36;
	reg [31:0] data_store_2_38;
	reg [31:0] data_store_2_40;
	reg [31:0] data_store_2_42;
	reg [0:0] data_store_2_44;
	reg [0:0] data_store_2_46;
	reg [31:0] data_store_2_48;
	reg [0:0] data_store_2_50;
	reg [31:0] data_store_2_52;
	reg [31:0] data_store_3_54;
	reg [31:0] data_store_3_56;
	reg [31:0] data_store_3_58;
	reg [31:0] data_store_3_60;
	reg [0:0] data_store_3_62;
	reg [0:0] data_store_3_64;
	reg [31:0] data_store_3_66;
	reg [0:0] data_store_3_68;
	reg [31:0] data_store_3_70;
	reg [31:0] data_store_4_72;
	reg [31:0] data_store_4_74;
	reg [31:0] data_store_4_76;
	reg [31:0] data_store_4_78;
	reg [0:0] data_store_4_80;
	reg [0:0] data_store_4_82;
	reg [31:0] data_store_4_84;
	reg [0:0] data_store_4_86;
	reg [31:0] data_store_4_88;
	reg [31:0] global_state;
	reg [0:0] icmp_tmp_5;
	reg [31:0] phi_tmp_0;
	reg [31:0] state_0_entry_BB_reg;
	reg [0:0] state_0_is_active;
	reg [31:0] state_0_last_BB_reg;
	reg [31:0] state_0_last_state;
	reg [31:0] state_1_entry_BB_reg;
	reg [0:0] state_1_is_active;
	reg [31:0] state_1_last_BB_reg;
	reg [31:0] state_1_last_state;
	reg [31:0] state_2_entry_BB_reg;
	reg [0:0] state_2_is_active;
	reg [31:0] state_2_last_BB_reg;
	reg [31:0] state_2_last_state;
	reg [31:0] state_3_entry_BB_reg;
	reg [0:0] state_3_is_active;
	reg [31:0] state_3_last_BB_reg;
	reg [31:0] state_3_last_state;
	reg [31:0] state_4_entry_BB_reg;
	reg [0:0] state_4_is_active;
	reg [31:0] state_4_last_BB_reg;
	reg [31:0] state_4_last_state;

	// controller for add_add_12.add_in0_add_12
	// controller for add_add_12.add_in1_add_12
	// Insensitive connections
	always @(*) begin
		add_in0_add_12 = valid ? rdata_ram_0 : rdata_ram_0;
		add_in1_add_12 = valid ? tmp_output_210_out_data : tmp_output_210_out_data;
	end
	// controller for add_add_14.add_in0_add_14
	// controller for add_add_14.add_in1_add_14
	// Insensitive connections
	always @(*) begin
		add_in0_add_14 = valid ? data_in_3_55_out_data : data_in_3_55_out_data;
		add_in1_add_14 = valid ? 32'd1 : 32'd1;
	end
	// controller for andOp_100.andOp_100_in0
	// controller for andOp_100.andOp_100_in1
	// Insensitive connections
	always @(*) begin
		andOp_100_in0 = valid ? andOp_99_out : andOp_99_out;
		andOp_100_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_102.andOp_102_in0
	// controller for andOp_102.andOp_102_in1
	// Insensitive connections
	always @(*) begin
		andOp_102_in0 = valid ? andOp_100_out : andOp_100_out;
		andOp_102_in1 = valid ? in_read_ready : in_read_ready;
	end
	// controller for andOp_104.andOp_104_in0
	// controller for andOp_104.andOp_104_in1
	// Insensitive connections
	always @(*) begin
		andOp_104_in0 = valid ? andOp_100_out : andOp_100_out;
		andOp_104_in1 = valid ? notOp_103_out : notOp_103_out;
	end
	// controller for andOp_105.andOp_105_in0
	// controller for andOp_105.andOp_105_in1
	// Insensitive connections
	always @(*) begin
		andOp_105_in0 = valid ? bb_0_active_in_state_1_out_data : bb_0_active_in_state_1_out_data;
		andOp_105_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_106.andOp_106_in0
	// controller for andOp_106.andOp_106_in1
	// Insensitive connections
	always @(*) begin
		andOp_106_in0 = valid ? andOp_105_out : andOp_105_out;
		andOp_106_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_108.andOp_108_in0
	// controller for andOp_108.andOp_108_in1
	// Insensitive connections
	always @(*) begin
		andOp_108_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_108_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_109.andOp_109_in0
	// controller for andOp_109.andOp_109_in1
	// Insensitive connections
	always @(*) begin
		andOp_109_in0 = valid ? andOp_108_out : andOp_108_out;
		andOp_109_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_111.andOp_111_in0
	// controller for andOp_111.andOp_111_in1
	// Insensitive connections
	always @(*) begin
		andOp_111_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_111_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_112.andOp_112_in0
	// controller for andOp_112.andOp_112_in1
	// Insensitive connections
	always @(*) begin
		andOp_112_in0 = valid ? andOp_111_out : andOp_111_out;
		andOp_112_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_114.andOp_114_in0
	// controller for andOp_114.andOp_114_in1
	// Insensitive connections
	always @(*) begin
		andOp_114_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_114_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_115.andOp_115_in0
	// controller for andOp_115.andOp_115_in1
	// Insensitive connections
	always @(*) begin
		andOp_115_in0 = valid ? andOp_114_out : andOp_114_out;
		andOp_115_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_117.andOp_117_in0
	// controller for andOp_117.andOp_117_in1
	// Insensitive connections
	always @(*) begin
		andOp_117_in0 = valid ? andOp_115_out : andOp_115_out;
		andOp_117_in1 = valid ? data_in_4_81_out_data : data_in_4_81_out_data;
	end
	// controller for andOp_119.andOp_119_in0
	// controller for andOp_119.andOp_119_in1
	// Insensitive connections
	always @(*) begin
		andOp_119_in0 = valid ? andOp_115_out : andOp_115_out;
		andOp_119_in1 = valid ? notOp_118_out : notOp_118_out;
	end
	// controller for andOp_120.andOp_120_in0
	// controller for andOp_120.andOp_120_in1
	// Insensitive connections
	always @(*) begin
		andOp_120_in0 = valid ? bb_1_active_in_state_4_out_data : bb_1_active_in_state_4_out_data;
		andOp_120_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_121.andOp_121_in0
	// controller for andOp_121.andOp_121_in1
	// Insensitive connections
	always @(*) begin
		andOp_121_in0 = valid ? andOp_120_out : andOp_120_out;
		andOp_121_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_123.andOp_123_in0
	// controller for andOp_123.andOp_123_in1
	// Insensitive connections
	always @(*) begin
		andOp_123_in0 = valid ? bb_5_active_in_state_4_out_data : bb_5_active_in_state_4_out_data;
		andOp_123_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_124.andOp_124_in0
	// controller for andOp_124.andOp_124_in1
	// Insensitive connections
	always @(*) begin
		andOp_124_in0 = valid ? andOp_123_out : andOp_123_out;
		andOp_124_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_126.andOp_126_in0
	// controller for andOp_126.andOp_126_in1
	// Insensitive connections
	always @(*) begin
		andOp_126_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
		andOp_126_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_127.andOp_127_in0
	// controller for andOp_127.andOp_127_in1
	// Insensitive connections
	always @(*) begin
		andOp_127_in0 = valid ? andOp_126_out : andOp_126_out;
		andOp_127_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_129.andOp_129_in0
	// controller for andOp_129.andOp_129_in1
	// Insensitive connections
	always @(*) begin
		andOp_129_in0 = valid ? andOp_127_out : andOp_127_out;
		andOp_129_in1 = valid ? out_write_ready : out_write_ready;
	end
	// controller for andOp_131.andOp_131_in0
	// controller for andOp_131.andOp_131_in1
	// Insensitive connections
	always @(*) begin
		andOp_131_in0 = valid ? andOp_127_out : andOp_127_out;
		andOp_131_in1 = valid ? notOp_130_out : notOp_130_out;
	end
	// controller for andOp_132.andOp_132_in0
	// controller for andOp_132.andOp_132_in1
	// Insensitive connections
	always @(*) begin
		andOp_132_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_132_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_133.andOp_133_in0
	// controller for andOp_133.andOp_133_in1
	// Insensitive connections
	always @(*) begin
		andOp_133_in0 = valid ? andOp_132_out : andOp_132_out;
		andOp_133_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_135.andOp_135_in0
	// controller for andOp_135.andOp_135_in1
	// Insensitive connections
	always @(*) begin
		andOp_135_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_135_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_136.andOp_136_in0
	// controller for andOp_136.andOp_136_in1
	// Insensitive connections
	always @(*) begin
		andOp_136_in0 = valid ? andOp_135_out : andOp_135_out;
		andOp_136_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_138.andOp_138_in0
	// controller for andOp_138.andOp_138_in1
	// Insensitive connections
	always @(*) begin
		andOp_138_in0 = valid ? andOp_136_out : andOp_136_out;
		andOp_138_in1 = valid ? data_in_4_81_out_data : data_in_4_81_out_data;
	end
	// controller for andOp_140.andOp_140_in0
	// controller for andOp_140.andOp_140_in1
	// Insensitive connections
	always @(*) begin
		andOp_140_in0 = valid ? andOp_136_out : andOp_136_out;
		andOp_140_in1 = valid ? notOp_139_out : notOp_139_out;
	end
	// controller for andOp_167.andOp_167_in0
	// controller for andOp_167.andOp_167_in1
	// Insensitive connections
	always @(*) begin
		andOp_167_in0 = valid ? notOp_166_out : notOp_166_out;
		andOp_167_in1 = valid ? andOp_91_out : andOp_91_out;
	end
	// controller for andOp_170.andOp_170_in0
	// controller for andOp_170.andOp_170_in1
	// Insensitive connections
	always @(*) begin
		andOp_170_in0 = valid ? notOp_169_out : notOp_169_out;
		andOp_170_in1 = valid ? andOp_94_out : andOp_94_out;
	end
	// controller for andOp_173.andOp_173_in0
	// controller for andOp_173.andOp_173_in1
	// Insensitive connections
	always @(*) begin
		andOp_173_in0 = valid ? notOp_172_out : notOp_172_out;
		andOp_173_in1 = valid ? andOp_97_out : andOp_97_out;
	end
	// controller for andOp_179.andOp_179_in0
	// controller for andOp_179.andOp_179_in1
	// Insensitive connections
	always @(*) begin
		andOp_179_in0 = valid ? notOp_178_out : notOp_178_out;
		andOp_179_in1 = valid ? andOp_109_out : andOp_109_out;
	end
	// controller for andOp_182.andOp_182_in0
	// controller for andOp_182.andOp_182_in1
	// Insensitive connections
	always @(*) begin
		andOp_182_in0 = valid ? notOp_181_out : notOp_181_out;
		andOp_182_in1 = valid ? andOp_117_out : andOp_117_out;
	end
	// controller for andOp_185.andOp_185_in0
	// controller for andOp_185.andOp_185_in1
	// Insensitive connections
	always @(*) begin
		andOp_185_in0 = valid ? notOp_184_out : notOp_184_out;
		andOp_185_in1 = valid ? andOp_121_out : andOp_121_out;
	end
	// controller for andOp_188.andOp_188_in0
	// controller for andOp_188.andOp_188_in1
	// Insensitive connections
	always @(*) begin
		andOp_188_in0 = valid ? notOp_187_out : notOp_187_out;
		andOp_188_in1 = valid ? andOp_124_out : andOp_124_out;
	end
	// controller for andOp_191.andOp_191_in0
	// controller for andOp_191.andOp_191_in1
	// Insensitive connections
	always @(*) begin
		andOp_191_in0 = valid ? notOp_190_out : notOp_190_out;
		andOp_191_in1 = valid ? andOp_129_out : andOp_129_out;
	end
	// controller for andOp_195.andOp_195_in0
	// controller for andOp_195.andOp_195_in1
	// Insensitive connections
	always @(*) begin
		andOp_195_in0 = valid ? notOp_194_out : notOp_194_out;
		andOp_195_in1 = valid ? andOp_133_out : andOp_133_out;
	end
	// controller for andOp_196.andOp_196_in0
	// controller for andOp_196.andOp_196_in1
	// Insensitive connections
	always @(*) begin
		andOp_196_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_196_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_197.andOp_197_in0
	// controller for andOp_197.andOp_197_in1
	// Insensitive connections
	always @(*) begin
		andOp_197_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_197_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_198.andOp_198_in0
	// controller for andOp_198.andOp_198_in1
	// Insensitive connections
	always @(*) begin
		andOp_198_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_198_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_199.andOp_199_in0
	// controller for andOp_199.andOp_199_in1
	// Insensitive connections
	always @(*) begin
		andOp_199_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_199_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_200.andOp_200_in0
	// controller for andOp_200.andOp_200_in1
	// Insensitive connections
	always @(*) begin
		andOp_200_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_200_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_201.andOp_201_in0
	// controller for andOp_201.andOp_201_in1
	// Insensitive connections
	always @(*) begin
		andOp_201_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_201_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_202.andOp_202_in0
	// controller for andOp_202.andOp_202_in1
	// Insensitive connections
	always @(*) begin
		andOp_202_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_202_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_203.andOp_203_in0
	// controller for andOp_203.andOp_203_in1
	// Insensitive connections
	always @(*) begin
		andOp_203_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_203_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_206.andOp_206_in0
	// controller for andOp_206.andOp_206_in1
	// Insensitive connections
	always @(*) begin
		andOp_206_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
		andOp_206_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_207.andOp_207_in0
	// controller for andOp_207.andOp_207_in1
	// Insensitive connections
	always @(*) begin
		andOp_207_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_207_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_208.andOp_208_in0
	// controller for andOp_208.andOp_208_in1
	// Insensitive connections
	always @(*) begin
		andOp_208_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_208_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_209.andOp_209_in0
	// controller for andOp_209.andOp_209_in1
	// Insensitive connections
	always @(*) begin
		andOp_209_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_209_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_212.andOp_212_in0
	// controller for andOp_212.andOp_212_in1
	// Insensitive connections
	always @(*) begin
		andOp_212_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_212_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_213.andOp_213_in0
	// controller for andOp_213.andOp_213_in1
	// Insensitive connections
	always @(*) begin
		andOp_213_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_213_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_214.andOp_214_in0
	// controller for andOp_214.andOp_214_in1
	// Insensitive connections
	always @(*) begin
		andOp_214_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_214_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_215.andOp_215_in0
	// controller for andOp_215.andOp_215_in1
	// Insensitive connections
	always @(*) begin
		andOp_215_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_215_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_216.andOp_216_in0
	// controller for andOp_216.andOp_216_in1
	// Insensitive connections
	always @(*) begin
		andOp_216_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_216_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_217.andOp_217_in0
	// controller for andOp_217.andOp_217_in1
	// Insensitive connections
	always @(*) begin
		andOp_217_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
		andOp_217_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_218.andOp_218_in0
	// controller for andOp_218.andOp_218_in1
	// Insensitive connections
	always @(*) begin
		andOp_218_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_218_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_219.andOp_219_in0
	// controller for andOp_219.andOp_219_in1
	// Insensitive connections
	always @(*) begin
		andOp_219_in0 = valid ? bb_0_active_in_state_0_out_data : bb_0_active_in_state_0_out_data;
		andOp_219_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_220.andOp_220_in0
	// controller for andOp_220.andOp_220_in1
	// Insensitive connections
	always @(*) begin
		andOp_220_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_220_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_221.andOp_221_in0
	// controller for andOp_221.andOp_221_in1
	// Insensitive connections
	always @(*) begin
		andOp_221_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_221_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_222.andOp_222_in0
	// controller for andOp_222.andOp_222_in1
	// Insensitive connections
	always @(*) begin
		andOp_222_in0 = valid ? bb_2_active_in_state_4_out_data : bb_2_active_in_state_4_out_data;
		andOp_222_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_224.andOp_224_in0
	// controller for andOp_224.andOp_224_in1
	// Insensitive connections
	always @(*) begin
		andOp_224_in0 = valid ? notOp_223_out : notOp_223_out;
		andOp_224_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_226.andOp_226_in0
	// controller for andOp_226.andOp_226_in1
	// Insensitive connections
	always @(*) begin
		andOp_226_in0 = valid ? notOp_225_out : notOp_225_out;
		andOp_226_in1 = valid ? andOp_224_out : andOp_224_out;
	end
	// controller for andOp_228.andOp_228_in0
	// controller for andOp_228.andOp_228_in1
	// Insensitive connections
	always @(*) begin
		andOp_228_in0 = valid ? notOp_227_out : notOp_227_out;
		andOp_228_in1 = valid ? andOp_226_out : andOp_226_out;
	end
	// controller for andOp_230.andOp_230_in0
	// controller for andOp_230.andOp_230_in1
	// Insensitive connections
	always @(*) begin
		andOp_230_in0 = valid ? notOp_229_out : notOp_229_out;
		andOp_230_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_232.andOp_232_in0
	// controller for andOp_232.andOp_232_in1
	// Insensitive connections
	always @(*) begin
		andOp_232_in0 = valid ? notOp_231_out : notOp_231_out;
		andOp_232_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_234.andOp_234_in0
	// controller for andOp_234.andOp_234_in1
	// Insensitive connections
	always @(*) begin
		andOp_234_in0 = valid ? notOp_233_out : notOp_233_out;
		andOp_234_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_236.andOp_236_in0
	// controller for andOp_236.andOp_236_in1
	// Insensitive connections
	always @(*) begin
		andOp_236_in0 = valid ? notOp_235_out : notOp_235_out;
		andOp_236_in1 = valid ? andOp_234_out : andOp_234_out;
	end
	// controller for andOp_238.andOp_238_in0
	// controller for andOp_238.andOp_238_in1
	// Insensitive connections
	always @(*) begin
		andOp_238_in0 = valid ? notOp_237_out : notOp_237_out;
		andOp_238_in1 = valid ? andOp_236_out : andOp_236_out;
	end
	// controller for andOp_239.andOp_239_in0
	// controller for andOp_239.andOp_239_in1
	// Insensitive connections
	always @(*) begin
		andOp_239_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_239_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_240.andOp_240_in0
	// controller for andOp_240.andOp_240_in1
	// Insensitive connections
	always @(*) begin
		andOp_240_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_240_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_241.andOp_241_in0
	// controller for andOp_241.andOp_241_in1
	// Insensitive connections
	always @(*) begin
		andOp_241_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_241_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_242.andOp_242_in0
	// controller for andOp_242.andOp_242_in1
	// Insensitive connections
	always @(*) begin
		andOp_242_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_242_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_244.andOp_244_in0
	// controller for andOp_244.andOp_244_in1
	// Insensitive connections
	always @(*) begin
		andOp_244_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_244_in1 = valid ? eq_243_out : eq_243_out;
	end
	// controller for andOp_246.andOp_246_in0
	// controller for andOp_246.andOp_246_in1
	// Insensitive connections
	always @(*) begin
		andOp_246_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_246_in1 = valid ? eq_245_out : eq_245_out;
	end
	// controller for andOp_248.andOp_248_in0
	// controller for andOp_248.andOp_248_in1
	// Insensitive connections
	always @(*) begin
		andOp_248_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_248_in1 = valid ? eq_247_out : eq_247_out;
	end
	// controller for andOp_250.andOp_250_in0
	// controller for andOp_250.andOp_250_in1
	// Insensitive connections
	always @(*) begin
		andOp_250_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_250_in1 = valid ? eq_249_out : eq_249_out;
	end
	// controller for andOp_252.andOp_252_in0
	// controller for andOp_252.andOp_252_in1
	// Insensitive connections
	always @(*) begin
		andOp_252_in0 = valid ? state_0_is_active : state_0_is_active;
		andOp_252_in1 = valid ? eq_251_out : eq_251_out;
	end
	// controller for andOp_253.andOp_253_in0
	// controller for andOp_253.andOp_253_in1
	// Insensitive connections
	always @(*) begin
		andOp_253_in0 = valid ? 1'd0 : 1'd0;
		andOp_253_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_255.andOp_255_in0
	// controller for andOp_255.andOp_255_in1
	// Insensitive connections
	always @(*) begin
		andOp_255_in0 = valid ? andOp_253_out : andOp_253_out;
		andOp_255_in1 = valid ? eq_254_out : eq_254_out;
	end
	// controller for andOp_257.andOp_257_in0
	// controller for andOp_257.andOp_257_in1
	// Insensitive connections
	always @(*) begin
		andOp_257_in0 = valid ? andOp_253_out : andOp_253_out;
		andOp_257_in1 = valid ? notOp_256_out : notOp_256_out;
	end
	// controller for andOp_258.andOp_258_in0
	// controller for andOp_258.andOp_258_in1
	// Insensitive connections
	always @(*) begin
		andOp_258_in0 = valid ? 1'd0 : 1'd0;
		andOp_258_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_260.andOp_260_in0
	// controller for andOp_260.andOp_260_in1
	// Insensitive connections
	always @(*) begin
		andOp_260_in0 = valid ? andOp_258_out : andOp_258_out;
		andOp_260_in1 = valid ? eq_259_out : eq_259_out;
	end
	// controller for andOp_262.andOp_262_in0
	// controller for andOp_262.andOp_262_in1
	// Insensitive connections
	always @(*) begin
		andOp_262_in0 = valid ? andOp_258_out : andOp_258_out;
		andOp_262_in1 = valid ? notOp_261_out : notOp_261_out;
	end
	// controller for andOp_263.andOp_263_in0
	// controller for andOp_263.andOp_263_in1
	// Insensitive connections
	always @(*) begin
		andOp_263_in0 = valid ? 1'd0 : 1'd0;
		andOp_263_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_265.andOp_265_in0
	// controller for andOp_265.andOp_265_in1
	// Insensitive connections
	always @(*) begin
		andOp_265_in0 = valid ? andOp_263_out : andOp_263_out;
		andOp_265_in1 = valid ? eq_264_out : eq_264_out;
	end
	// controller for andOp_267.andOp_267_in0
	// controller for andOp_267.andOp_267_in1
	// Insensitive connections
	always @(*) begin
		andOp_267_in0 = valid ? andOp_263_out : andOp_263_out;
		andOp_267_in1 = valid ? notOp_266_out : notOp_266_out;
	end
	// controller for andOp_268.andOp_268_in0
	// controller for andOp_268.andOp_268_in1
	// Insensitive connections
	always @(*) begin
		andOp_268_in0 = valid ? 1'd0 : 1'd0;
		andOp_268_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_270.andOp_270_in0
	// controller for andOp_270.andOp_270_in1
	// Insensitive connections
	always @(*) begin
		andOp_270_in0 = valid ? andOp_268_out : andOp_268_out;
		andOp_270_in1 = valid ? eq_269_out : eq_269_out;
	end
	// controller for andOp_272.andOp_272_in0
	// controller for andOp_272.andOp_272_in1
	// Insensitive connections
	always @(*) begin
		andOp_272_in0 = valid ? andOp_268_out : andOp_268_out;
		andOp_272_in1 = valid ? notOp_271_out : notOp_271_out;
	end
	// controller for andOp_273.andOp_273_in0
	// controller for andOp_273.andOp_273_in1
	// Insensitive connections
	always @(*) begin
		andOp_273_in0 = valid ? 1'd0 : 1'd0;
		andOp_273_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_275.andOp_275_in0
	// controller for andOp_275.andOp_275_in1
	// Insensitive connections
	always @(*) begin
		andOp_275_in0 = valid ? andOp_273_out : andOp_273_out;
		andOp_275_in1 = valid ? eq_274_out : eq_274_out;
	end
	// controller for andOp_277.andOp_277_in0
	// controller for andOp_277.andOp_277_in1
	// Insensitive connections
	always @(*) begin
		andOp_277_in0 = valid ? andOp_273_out : andOp_273_out;
		andOp_277_in1 = valid ? notOp_276_out : notOp_276_out;
	end
	// controller for andOp_278.andOp_278_in0
	// controller for andOp_278.andOp_278_in1
	// Insensitive connections
	always @(*) begin
		andOp_278_in0 = valid ? 1'd0 : 1'd0;
		andOp_278_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_280.andOp_280_in0
	// controller for andOp_280.andOp_280_in1
	// Insensitive connections
	always @(*) begin
		andOp_280_in0 = valid ? andOp_278_out : andOp_278_out;
		andOp_280_in1 = valid ? eq_279_out : eq_279_out;
	end
	// controller for andOp_282.andOp_282_in0
	// controller for andOp_282.andOp_282_in1
	// Insensitive connections
	always @(*) begin
		andOp_282_in0 = valid ? andOp_278_out : andOp_278_out;
		andOp_282_in1 = valid ? notOp_281_out : notOp_281_out;
	end
	// controller for andOp_283.andOp_283_in0
	// controller for andOp_283.andOp_283_in1
	// Insensitive connections
	always @(*) begin
		andOp_283_in0 = valid ? 1'd0 : 1'd0;
		andOp_283_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_285.andOp_285_in0
	// controller for andOp_285.andOp_285_in1
	// Insensitive connections
	always @(*) begin
		andOp_285_in0 = valid ? andOp_283_out : andOp_283_out;
		andOp_285_in1 = valid ? eq_284_out : eq_284_out;
	end
	// controller for andOp_287.andOp_287_in0
	// controller for andOp_287.andOp_287_in1
	// Insensitive connections
	always @(*) begin
		andOp_287_in0 = valid ? andOp_283_out : andOp_283_out;
		andOp_287_in1 = valid ? notOp_286_out : notOp_286_out;
	end
	// controller for andOp_288.andOp_288_in0
	// controller for andOp_288.andOp_288_in1
	// Insensitive connections
	always @(*) begin
		andOp_288_in0 = valid ? 1'd0 : 1'd0;
		andOp_288_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_290.andOp_290_in0
	// controller for andOp_290.andOp_290_in1
	// Insensitive connections
	always @(*) begin
		andOp_290_in0 = valid ? andOp_288_out : andOp_288_out;
		andOp_290_in1 = valid ? eq_289_out : eq_289_out;
	end
	// controller for andOp_292.andOp_292_in0
	// controller for andOp_292.andOp_292_in1
	// Insensitive connections
	always @(*) begin
		andOp_292_in0 = valid ? andOp_288_out : andOp_288_out;
		andOp_292_in1 = valid ? notOp_291_out : notOp_291_out;
	end
	// controller for andOp_293.andOp_293_in0
	// controller for andOp_293.andOp_293_in1
	// Insensitive connections
	always @(*) begin
		andOp_293_in0 = valid ? 1'd0 : 1'd0;
		andOp_293_in1 = valid ? state_0_is_active : state_0_is_active;
	end
	// controller for andOp_295.andOp_295_in0
	// controller for andOp_295.andOp_295_in1
	// Insensitive connections
	always @(*) begin
		andOp_295_in0 = valid ? andOp_293_out : andOp_293_out;
		andOp_295_in1 = valid ? eq_294_out : eq_294_out;
	end
	// controller for andOp_297.andOp_297_in0
	// controller for andOp_297.andOp_297_in1
	// Insensitive connections
	always @(*) begin
		andOp_297_in0 = valid ? andOp_293_out : andOp_293_out;
		andOp_297_in1 = valid ? notOp_296_out : notOp_296_out;
	end
	// controller for andOp_299.andOp_299_in0
	// controller for andOp_299.andOp_299_in1
	// Insensitive connections
	always @(*) begin
		andOp_299_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_299_in1 = valid ? eq_298_out : eq_298_out;
	end
	// controller for andOp_301.andOp_301_in0
	// controller for andOp_301.andOp_301_in1
	// Insensitive connections
	always @(*) begin
		andOp_301_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_301_in1 = valid ? eq_300_out : eq_300_out;
	end
	// controller for andOp_303.andOp_303_in0
	// controller for andOp_303.andOp_303_in1
	// Insensitive connections
	always @(*) begin
		andOp_303_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_303_in1 = valid ? eq_302_out : eq_302_out;
	end
	// controller for andOp_305.andOp_305_in0
	// controller for andOp_305.andOp_305_in1
	// Insensitive connections
	always @(*) begin
		andOp_305_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_305_in1 = valid ? eq_304_out : eq_304_out;
	end
	// controller for andOp_307.andOp_307_in0
	// controller for andOp_307.andOp_307_in1
	// Insensitive connections
	always @(*) begin
		andOp_307_in0 = valid ? state_1_is_active : state_1_is_active;
		andOp_307_in1 = valid ? eq_306_out : eq_306_out;
	end
	// controller for andOp_308.andOp_308_in0
	// controller for andOp_308.andOp_308_in1
	// Insensitive connections
	always @(*) begin
		andOp_308_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_308_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_310.andOp_310_in0
	// controller for andOp_310.andOp_310_in1
	// Insensitive connections
	always @(*) begin
		andOp_310_in0 = valid ? andOp_308_out : andOp_308_out;
		andOp_310_in1 = valid ? eq_309_out : eq_309_out;
	end
	// controller for andOp_312.andOp_312_in0
	// controller for andOp_312.andOp_312_in1
	// Insensitive connections
	always @(*) begin
		andOp_312_in0 = valid ? andOp_308_out : andOp_308_out;
		andOp_312_in1 = valid ? notOp_311_out : notOp_311_out;
	end
	// controller for andOp_313.andOp_313_in0
	// controller for andOp_313.andOp_313_in1
	// Insensitive connections
	always @(*) begin
		andOp_313_in0 = valid ? 1'd0 : 1'd0;
		andOp_313_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_315.andOp_315_in0
	// controller for andOp_315.andOp_315_in1
	// Insensitive connections
	always @(*) begin
		andOp_315_in0 = valid ? andOp_313_out : andOp_313_out;
		andOp_315_in1 = valid ? eq_314_out : eq_314_out;
	end
	// controller for andOp_317.andOp_317_in0
	// controller for andOp_317.andOp_317_in1
	// Insensitive connections
	always @(*) begin
		andOp_317_in0 = valid ? andOp_313_out : andOp_313_out;
		andOp_317_in1 = valid ? notOp_316_out : notOp_316_out;
	end
	// controller for andOp_318.andOp_318_in0
	// controller for andOp_318.andOp_318_in1
	// Insensitive connections
	always @(*) begin
		andOp_318_in0 = valid ? 1'd0 : 1'd0;
		andOp_318_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_320.andOp_320_in0
	// controller for andOp_320.andOp_320_in1
	// Insensitive connections
	always @(*) begin
		andOp_320_in0 = valid ? andOp_318_out : andOp_318_out;
		andOp_320_in1 = valid ? eq_319_out : eq_319_out;
	end
	// controller for andOp_322.andOp_322_in0
	// controller for andOp_322.andOp_322_in1
	// Insensitive connections
	always @(*) begin
		andOp_322_in0 = valid ? andOp_318_out : andOp_318_out;
		andOp_322_in1 = valid ? notOp_321_out : notOp_321_out;
	end
	// controller for andOp_323.andOp_323_in0
	// controller for andOp_323.andOp_323_in1
	// Insensitive connections
	always @(*) begin
		andOp_323_in0 = valid ? 1'd0 : 1'd0;
		andOp_323_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_325.andOp_325_in0
	// controller for andOp_325.andOp_325_in1
	// Insensitive connections
	always @(*) begin
		andOp_325_in0 = valid ? andOp_323_out : andOp_323_out;
		andOp_325_in1 = valid ? eq_324_out : eq_324_out;
	end
	// controller for andOp_327.andOp_327_in0
	// controller for andOp_327.andOp_327_in1
	// Insensitive connections
	always @(*) begin
		andOp_327_in0 = valid ? andOp_323_out : andOp_323_out;
		andOp_327_in1 = valid ? notOp_326_out : notOp_326_out;
	end
	// controller for andOp_328.andOp_328_in0
	// controller for andOp_328.andOp_328_in1
	// Insensitive connections
	always @(*) begin
		andOp_328_in0 = valid ? 1'd0 : 1'd0;
		andOp_328_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_330.andOp_330_in0
	// controller for andOp_330.andOp_330_in1
	// Insensitive connections
	always @(*) begin
		andOp_330_in0 = valid ? andOp_328_out : andOp_328_out;
		andOp_330_in1 = valid ? eq_329_out : eq_329_out;
	end
	// controller for andOp_332.andOp_332_in0
	// controller for andOp_332.andOp_332_in1
	// Insensitive connections
	always @(*) begin
		andOp_332_in0 = valid ? andOp_328_out : andOp_328_out;
		andOp_332_in1 = valid ? notOp_331_out : notOp_331_out;
	end
	// controller for andOp_333.andOp_333_in0
	// controller for andOp_333.andOp_333_in1
	// Insensitive connections
	always @(*) begin
		andOp_333_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
		andOp_333_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_335.andOp_335_in0
	// controller for andOp_335.andOp_335_in1
	// Insensitive connections
	always @(*) begin
		andOp_335_in0 = valid ? andOp_333_out : andOp_333_out;
		andOp_335_in1 = valid ? eq_334_out : eq_334_out;
	end
	// controller for andOp_337.andOp_337_in0
	// controller for andOp_337.andOp_337_in1
	// Insensitive connections
	always @(*) begin
		andOp_337_in0 = valid ? andOp_333_out : andOp_333_out;
		andOp_337_in1 = valid ? notOp_336_out : notOp_336_out;
	end
	// controller for andOp_338.andOp_338_in0
	// controller for andOp_338.andOp_338_in1
	// Insensitive connections
	always @(*) begin
		andOp_338_in0 = valid ? 1'd0 : 1'd0;
		andOp_338_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_340.andOp_340_in0
	// controller for andOp_340.andOp_340_in1
	// Insensitive connections
	always @(*) begin
		andOp_340_in0 = valid ? andOp_338_out : andOp_338_out;
		andOp_340_in1 = valid ? eq_339_out : eq_339_out;
	end
	// controller for andOp_342.andOp_342_in0
	// controller for andOp_342.andOp_342_in1
	// Insensitive connections
	always @(*) begin
		andOp_342_in0 = valid ? andOp_338_out : andOp_338_out;
		andOp_342_in1 = valid ? notOp_341_out : notOp_341_out;
	end
	// controller for andOp_343.andOp_343_in0
	// controller for andOp_343.andOp_343_in1
	// Insensitive connections
	always @(*) begin
		andOp_343_in0 = valid ? 1'd0 : 1'd0;
		andOp_343_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_345.andOp_345_in0
	// controller for andOp_345.andOp_345_in1
	// Insensitive connections
	always @(*) begin
		andOp_345_in0 = valid ? andOp_343_out : andOp_343_out;
		andOp_345_in1 = valid ? eq_344_out : eq_344_out;
	end
	// controller for andOp_347.andOp_347_in0
	// controller for andOp_347.andOp_347_in1
	// Insensitive connections
	always @(*) begin
		andOp_347_in0 = valid ? andOp_343_out : andOp_343_out;
		andOp_347_in1 = valid ? notOp_346_out : notOp_346_out;
	end
	// controller for andOp_348.andOp_348_in0
	// controller for andOp_348.andOp_348_in1
	// Insensitive connections
	always @(*) begin
		andOp_348_in0 = valid ? 1'd0 : 1'd0;
		andOp_348_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_350.andOp_350_in0
	// controller for andOp_350.andOp_350_in1
	// Insensitive connections
	always @(*) begin
		andOp_350_in0 = valid ? andOp_348_out : andOp_348_out;
		andOp_350_in1 = valid ? eq_349_out : eq_349_out;
	end
	// controller for andOp_352.andOp_352_in0
	// controller for andOp_352.andOp_352_in1
	// Insensitive connections
	always @(*) begin
		andOp_352_in0 = valid ? andOp_348_out : andOp_348_out;
		andOp_352_in1 = valid ? notOp_351_out : notOp_351_out;
	end
	// controller for andOp_354.andOp_354_in0
	// controller for andOp_354.andOp_354_in1
	// Insensitive connections
	always @(*) begin
		andOp_354_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_354_in1 = valid ? eq_353_out : eq_353_out;
	end
	// controller for andOp_356.andOp_356_in0
	// controller for andOp_356.andOp_356_in1
	// Insensitive connections
	always @(*) begin
		andOp_356_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_356_in1 = valid ? eq_355_out : eq_355_out;
	end
	// controller for andOp_358.andOp_358_in0
	// controller for andOp_358.andOp_358_in1
	// Insensitive connections
	always @(*) begin
		andOp_358_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_358_in1 = valid ? eq_357_out : eq_357_out;
	end
	// controller for andOp_360.andOp_360_in0
	// controller for andOp_360.andOp_360_in1
	// Insensitive connections
	always @(*) begin
		andOp_360_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_360_in1 = valid ? eq_359_out : eq_359_out;
	end
	// controller for andOp_362.andOp_362_in0
	// controller for andOp_362.andOp_362_in1
	// Insensitive connections
	always @(*) begin
		andOp_362_in0 = valid ? state_2_is_active : state_2_is_active;
		andOp_362_in1 = valid ? eq_361_out : eq_361_out;
	end
	// controller for andOp_363.andOp_363_in0
	// controller for andOp_363.andOp_363_in1
	// Insensitive connections
	always @(*) begin
		andOp_363_in0 = valid ? 1'd0 : 1'd0;
		andOp_363_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_365.andOp_365_in0
	// controller for andOp_365.andOp_365_in1
	// Insensitive connections
	always @(*) begin
		andOp_365_in0 = valid ? andOp_363_out : andOp_363_out;
		andOp_365_in1 = valid ? eq_364_out : eq_364_out;
	end
	// controller for andOp_367.andOp_367_in0
	// controller for andOp_367.andOp_367_in1
	// Insensitive connections
	always @(*) begin
		andOp_367_in0 = valid ? andOp_363_out : andOp_363_out;
		andOp_367_in1 = valid ? notOp_366_out : notOp_366_out;
	end
	// controller for andOp_368.andOp_368_in0
	// controller for andOp_368.andOp_368_in1
	// Insensitive connections
	always @(*) begin
		andOp_368_in0 = valid ? 1'd0 : 1'd0;
		andOp_368_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_370.andOp_370_in0
	// controller for andOp_370.andOp_370_in1
	// Insensitive connections
	always @(*) begin
		andOp_370_in0 = valid ? andOp_368_out : andOp_368_out;
		andOp_370_in1 = valid ? eq_369_out : eq_369_out;
	end
	// controller for andOp_372.andOp_372_in0
	// controller for andOp_372.andOp_372_in1
	// Insensitive connections
	always @(*) begin
		andOp_372_in0 = valid ? andOp_368_out : andOp_368_out;
		andOp_372_in1 = valid ? notOp_371_out : notOp_371_out;
	end
	// controller for andOp_373.andOp_373_in0
	// controller for andOp_373.andOp_373_in1
	// Insensitive connections
	always @(*) begin
		andOp_373_in0 = valid ? 1'd0 : 1'd0;
		andOp_373_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_375.andOp_375_in0
	// controller for andOp_375.andOp_375_in1
	// Insensitive connections
	always @(*) begin
		andOp_375_in0 = valid ? andOp_373_out : andOp_373_out;
		andOp_375_in1 = valid ? eq_374_out : eq_374_out;
	end
	// controller for andOp_377.andOp_377_in0
	// controller for andOp_377.andOp_377_in1
	// Insensitive connections
	always @(*) begin
		andOp_377_in0 = valid ? andOp_373_out : andOp_373_out;
		andOp_377_in1 = valid ? notOp_376_out : notOp_376_out;
	end
	// controller for andOp_378.andOp_378_in0
	// controller for andOp_378.andOp_378_in1
	// Insensitive connections
	always @(*) begin
		andOp_378_in0 = valid ? 1'd0 : 1'd0;
		andOp_378_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_380.andOp_380_in0
	// controller for andOp_380.andOp_380_in1
	// Insensitive connections
	always @(*) begin
		andOp_380_in0 = valid ? andOp_378_out : andOp_378_out;
		andOp_380_in1 = valid ? eq_379_out : eq_379_out;
	end
	// controller for andOp_382.andOp_382_in0
	// controller for andOp_382.andOp_382_in1
	// Insensitive connections
	always @(*) begin
		andOp_382_in0 = valid ? andOp_378_out : andOp_378_out;
		andOp_382_in1 = valid ? notOp_381_out : notOp_381_out;
	end
	// controller for andOp_383.andOp_383_in0
	// controller for andOp_383.andOp_383_in1
	// Insensitive connections
	always @(*) begin
		andOp_383_in0 = valid ? 1'd0 : 1'd0;
		andOp_383_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_385.andOp_385_in0
	// controller for andOp_385.andOp_385_in1
	// Insensitive connections
	always @(*) begin
		andOp_385_in0 = valid ? andOp_383_out : andOp_383_out;
		andOp_385_in1 = valid ? eq_384_out : eq_384_out;
	end
	// controller for andOp_387.andOp_387_in0
	// controller for andOp_387.andOp_387_in1
	// Insensitive connections
	always @(*) begin
		andOp_387_in0 = valid ? andOp_383_out : andOp_383_out;
		andOp_387_in1 = valid ? notOp_386_out : notOp_386_out;
	end
	// controller for andOp_388.andOp_388_in0
	// controller for andOp_388.andOp_388_in1
	// Insensitive connections
	always @(*) begin
		andOp_388_in0 = valid ? 1'd0 : 1'd0;
		andOp_388_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_390.andOp_390_in0
	// controller for andOp_390.andOp_390_in1
	// Insensitive connections
	always @(*) begin
		andOp_390_in0 = valid ? andOp_388_out : andOp_388_out;
		andOp_390_in1 = valid ? eq_389_out : eq_389_out;
	end
	// controller for andOp_392.andOp_392_in0
	// controller for andOp_392.andOp_392_in1
	// Insensitive connections
	always @(*) begin
		andOp_392_in0 = valid ? andOp_388_out : andOp_388_out;
		andOp_392_in1 = valid ? notOp_391_out : notOp_391_out;
	end
	// controller for andOp_393.andOp_393_in0
	// controller for andOp_393.andOp_393_in1
	// Insensitive connections
	always @(*) begin
		andOp_393_in0 = valid ? bb_10_active_in_state_2_out_data : bb_10_active_in_state_2_out_data;
		andOp_393_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_395.andOp_395_in0
	// controller for andOp_395.andOp_395_in1
	// Insensitive connections
	always @(*) begin
		andOp_395_in0 = valid ? andOp_393_out : andOp_393_out;
		andOp_395_in1 = valid ? eq_394_out : eq_394_out;
	end
	// controller for andOp_397.andOp_397_in0
	// controller for andOp_397.andOp_397_in1
	// Insensitive connections
	always @(*) begin
		andOp_397_in0 = valid ? andOp_393_out : andOp_393_out;
		andOp_397_in1 = valid ? notOp_396_out : notOp_396_out;
	end
	// controller for andOp_398.andOp_398_in0
	// controller for andOp_398.andOp_398_in1
	// Insensitive connections
	always @(*) begin
		andOp_398_in0 = valid ? 1'd0 : 1'd0;
		andOp_398_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_400.andOp_400_in0
	// controller for andOp_400.andOp_400_in1
	// Insensitive connections
	always @(*) begin
		andOp_400_in0 = valid ? andOp_398_out : andOp_398_out;
		andOp_400_in1 = valid ? eq_399_out : eq_399_out;
	end
	// controller for andOp_402.andOp_402_in0
	// controller for andOp_402.andOp_402_in1
	// Insensitive connections
	always @(*) begin
		andOp_402_in0 = valid ? andOp_398_out : andOp_398_out;
		andOp_402_in1 = valid ? notOp_401_out : notOp_401_out;
	end
	// controller for andOp_403.andOp_403_in0
	// controller for andOp_403.andOp_403_in1
	// Insensitive connections
	always @(*) begin
		andOp_403_in0 = valid ? 1'd0 : 1'd0;
		andOp_403_in1 = valid ? state_2_is_active : state_2_is_active;
	end
	// controller for andOp_405.andOp_405_in0
	// controller for andOp_405.andOp_405_in1
	// Insensitive connections
	always @(*) begin
		andOp_405_in0 = valid ? andOp_403_out : andOp_403_out;
		andOp_405_in1 = valid ? eq_404_out : eq_404_out;
	end
	// controller for andOp_407.andOp_407_in0
	// controller for andOp_407.andOp_407_in1
	// Insensitive connections
	always @(*) begin
		andOp_407_in0 = valid ? andOp_403_out : andOp_403_out;
		andOp_407_in1 = valid ? notOp_406_out : notOp_406_out;
	end
	// controller for andOp_409.andOp_409_in0
	// controller for andOp_409.andOp_409_in1
	// Insensitive connections
	always @(*) begin
		andOp_409_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_409_in1 = valid ? eq_408_out : eq_408_out;
	end
	// controller for andOp_411.andOp_411_in0
	// controller for andOp_411.andOp_411_in1
	// Insensitive connections
	always @(*) begin
		andOp_411_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_411_in1 = valid ? eq_410_out : eq_410_out;
	end
	// controller for andOp_413.andOp_413_in0
	// controller for andOp_413.andOp_413_in1
	// Insensitive connections
	always @(*) begin
		andOp_413_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_413_in1 = valid ? eq_412_out : eq_412_out;
	end
	// controller for andOp_415.andOp_415_in0
	// controller for andOp_415.andOp_415_in1
	// Insensitive connections
	always @(*) begin
		andOp_415_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_415_in1 = valid ? eq_414_out : eq_414_out;
	end
	// controller for andOp_417.andOp_417_in0
	// controller for andOp_417.andOp_417_in1
	// Insensitive connections
	always @(*) begin
		andOp_417_in0 = valid ? state_3_is_active : state_3_is_active;
		andOp_417_in1 = valid ? eq_416_out : eq_416_out;
	end
	// controller for andOp_418.andOp_418_in0
	// controller for andOp_418.andOp_418_in1
	// Insensitive connections
	always @(*) begin
		andOp_418_in0 = valid ? 1'd0 : 1'd0;
		andOp_418_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_420.andOp_420_in0
	// controller for andOp_420.andOp_420_in1
	// Insensitive connections
	always @(*) begin
		andOp_420_in0 = valid ? andOp_418_out : andOp_418_out;
		andOp_420_in1 = valid ? eq_419_out : eq_419_out;
	end
	// controller for andOp_422.andOp_422_in0
	// controller for andOp_422.andOp_422_in1
	// Insensitive connections
	always @(*) begin
		andOp_422_in0 = valid ? andOp_418_out : andOp_418_out;
		andOp_422_in1 = valid ? notOp_421_out : notOp_421_out;
	end
	// controller for andOp_423.andOp_423_in0
	// controller for andOp_423.andOp_423_in1
	// Insensitive connections
	always @(*) begin
		andOp_423_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_423_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_425.andOp_425_in0
	// controller for andOp_425.andOp_425_in1
	// Insensitive connections
	always @(*) begin
		andOp_425_in0 = valid ? andOp_423_out : andOp_423_out;
		andOp_425_in1 = valid ? eq_424_out : eq_424_out;
	end
	// controller for andOp_427.andOp_427_in0
	// controller for andOp_427.andOp_427_in1
	// Insensitive connections
	always @(*) begin
		andOp_427_in0 = valid ? andOp_423_out : andOp_423_out;
		andOp_427_in1 = valid ? notOp_426_out : notOp_426_out;
	end
	// controller for andOp_428.andOp_428_in0
	// controller for andOp_428.andOp_428_in1
	// Insensitive connections
	always @(*) begin
		andOp_428_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_428_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_430.andOp_430_in0
	// controller for andOp_430.andOp_430_in1
	// Insensitive connections
	always @(*) begin
		andOp_430_in0 = valid ? andOp_428_out : andOp_428_out;
		andOp_430_in1 = valid ? eq_429_out : eq_429_out;
	end
	// controller for andOp_432.andOp_432_in0
	// controller for andOp_432.andOp_432_in1
	// Insensitive connections
	always @(*) begin
		andOp_432_in0 = valid ? andOp_428_out : andOp_428_out;
		andOp_432_in1 = valid ? notOp_431_out : notOp_431_out;
	end
	// controller for andOp_433.andOp_433_in0
	// controller for andOp_433.andOp_433_in1
	// Insensitive connections
	always @(*) begin
		andOp_433_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_433_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_435.andOp_435_in0
	// controller for andOp_435.andOp_435_in1
	// Insensitive connections
	always @(*) begin
		andOp_435_in0 = valid ? andOp_433_out : andOp_433_out;
		andOp_435_in1 = valid ? eq_434_out : eq_434_out;
	end
	// controller for andOp_437.andOp_437_in0
	// controller for andOp_437.andOp_437_in1
	// Insensitive connections
	always @(*) begin
		andOp_437_in0 = valid ? andOp_433_out : andOp_433_out;
		andOp_437_in1 = valid ? notOp_436_out : notOp_436_out;
	end
	// controller for andOp_438.andOp_438_in0
	// controller for andOp_438.andOp_438_in1
	// Insensitive connections
	always @(*) begin
		andOp_438_in0 = valid ? bb_4_active_in_state_3_out_data : bb_4_active_in_state_3_out_data;
		andOp_438_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_440.andOp_440_in0
	// controller for andOp_440.andOp_440_in1
	// Insensitive connections
	always @(*) begin
		andOp_440_in0 = valid ? andOp_438_out : andOp_438_out;
		andOp_440_in1 = valid ? eq_439_out : eq_439_out;
	end
	// controller for andOp_442.andOp_442_in0
	// controller for andOp_442.andOp_442_in1
	// Insensitive connections
	always @(*) begin
		andOp_442_in0 = valid ? andOp_438_out : andOp_438_out;
		andOp_442_in1 = valid ? notOp_441_out : notOp_441_out;
	end
	// controller for andOp_443.andOp_443_in0
	// controller for andOp_443.andOp_443_in1
	// Insensitive connections
	always @(*) begin
		andOp_443_in0 = valid ? 1'd0 : 1'd0;
		andOp_443_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_445.andOp_445_in0
	// controller for andOp_445.andOp_445_in1
	// Insensitive connections
	always @(*) begin
		andOp_445_in0 = valid ? andOp_443_out : andOp_443_out;
		andOp_445_in1 = valid ? eq_444_out : eq_444_out;
	end
	// controller for andOp_447.andOp_447_in0
	// controller for andOp_447.andOp_447_in1
	// Insensitive connections
	always @(*) begin
		andOp_447_in0 = valid ? andOp_443_out : andOp_443_out;
		andOp_447_in1 = valid ? notOp_446_out : notOp_446_out;
	end
	// controller for andOp_448.andOp_448_in0
	// controller for andOp_448.andOp_448_in1
	// Insensitive connections
	always @(*) begin
		andOp_448_in0 = valid ? bb_10_active_in_state_3_out_data : bb_10_active_in_state_3_out_data;
		andOp_448_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_450.andOp_450_in0
	// controller for andOp_450.andOp_450_in1
	// Insensitive connections
	always @(*) begin
		andOp_450_in0 = valid ? andOp_448_out : andOp_448_out;
		andOp_450_in1 = valid ? eq_449_out : eq_449_out;
	end
	// controller for andOp_452.andOp_452_in0
	// controller for andOp_452.andOp_452_in1
	// Insensitive connections
	always @(*) begin
		andOp_452_in0 = valid ? andOp_448_out : andOp_448_out;
		andOp_452_in1 = valid ? notOp_451_out : notOp_451_out;
	end
	// controller for andOp_453.andOp_453_in0
	// controller for andOp_453.andOp_453_in1
	// Insensitive connections
	always @(*) begin
		andOp_453_in0 = valid ? 1'd0 : 1'd0;
		andOp_453_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_455.andOp_455_in0
	// controller for andOp_455.andOp_455_in1
	// Insensitive connections
	always @(*) begin
		andOp_455_in0 = valid ? andOp_453_out : andOp_453_out;
		andOp_455_in1 = valid ? eq_454_out : eq_454_out;
	end
	// controller for andOp_457.andOp_457_in0
	// controller for andOp_457.andOp_457_in1
	// Insensitive connections
	always @(*) begin
		andOp_457_in0 = valid ? andOp_453_out : andOp_453_out;
		andOp_457_in1 = valid ? notOp_456_out : notOp_456_out;
	end
	// controller for andOp_458.andOp_458_in0
	// controller for andOp_458.andOp_458_in1
	// Insensitive connections
	always @(*) begin
		andOp_458_in0 = valid ? 1'd0 : 1'd0;
		andOp_458_in1 = valid ? state_3_is_active : state_3_is_active;
	end
	// controller for andOp_460.andOp_460_in0
	// controller for andOp_460.andOp_460_in1
	// Insensitive connections
	always @(*) begin
		andOp_460_in0 = valid ? andOp_458_out : andOp_458_out;
		andOp_460_in1 = valid ? eq_459_out : eq_459_out;
	end
	// controller for andOp_462.andOp_462_in0
	// controller for andOp_462.andOp_462_in1
	// Insensitive connections
	always @(*) begin
		andOp_462_in0 = valid ? andOp_458_out : andOp_458_out;
		andOp_462_in1 = valid ? notOp_461_out : notOp_461_out;
	end
	// controller for andOp_464.andOp_464_in0
	// controller for andOp_464.andOp_464_in1
	// Insensitive connections
	always @(*) begin
		andOp_464_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_464_in1 = valid ? eq_463_out : eq_463_out;
	end
	// controller for andOp_466.andOp_466_in0
	// controller for andOp_466.andOp_466_in1
	// Insensitive connections
	always @(*) begin
		andOp_466_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_466_in1 = valid ? eq_465_out : eq_465_out;
	end
	// controller for andOp_468.andOp_468_in0
	// controller for andOp_468.andOp_468_in1
	// Insensitive connections
	always @(*) begin
		andOp_468_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_468_in1 = valid ? eq_467_out : eq_467_out;
	end
	// controller for andOp_470.andOp_470_in0
	// controller for andOp_470.andOp_470_in1
	// Insensitive connections
	always @(*) begin
		andOp_470_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_470_in1 = valid ? eq_469_out : eq_469_out;
	end
	// controller for andOp_472.andOp_472_in0
	// controller for andOp_472.andOp_472_in1
	// Insensitive connections
	always @(*) begin
		andOp_472_in0 = valid ? state_4_is_active : state_4_is_active;
		andOp_472_in1 = valid ? eq_471_out : eq_471_out;
	end
	// controller for andOp_473.andOp_473_in0
	// controller for andOp_473.andOp_473_in1
	// Insensitive connections
	always @(*) begin
		andOp_473_in0 = valid ? 1'd0 : 1'd0;
		andOp_473_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_475.andOp_475_in0
	// controller for andOp_475.andOp_475_in1
	// Insensitive connections
	always @(*) begin
		andOp_475_in0 = valid ? andOp_473_out : andOp_473_out;
		andOp_475_in1 = valid ? eq_474_out : eq_474_out;
	end
	// controller for andOp_477.andOp_477_in0
	// controller for andOp_477.andOp_477_in1
	// Insensitive connections
	always @(*) begin
		andOp_477_in0 = valid ? andOp_473_out : andOp_473_out;
		andOp_477_in1 = valid ? notOp_476_out : notOp_476_out;
	end
	// controller for andOp_478.andOp_478_in0
	// controller for andOp_478.andOp_478_in1
	// Insensitive connections
	always @(*) begin
		andOp_478_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_478_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_480.andOp_480_in0
	// controller for andOp_480.andOp_480_in1
	// Insensitive connections
	always @(*) begin
		andOp_480_in0 = valid ? andOp_478_out : andOp_478_out;
		andOp_480_in1 = valid ? eq_479_out : eq_479_out;
	end
	// controller for andOp_482.andOp_482_in0
	// controller for andOp_482.andOp_482_in1
	// Insensitive connections
	always @(*) begin
		andOp_482_in0 = valid ? andOp_478_out : andOp_478_out;
		andOp_482_in1 = valid ? notOp_481_out : notOp_481_out;
	end
	// controller for andOp_483.andOp_483_in0
	// controller for andOp_483.andOp_483_in1
	// Insensitive connections
	always @(*) begin
		andOp_483_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_483_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_485.andOp_485_in0
	// controller for andOp_485.andOp_485_in1
	// Insensitive connections
	always @(*) begin
		andOp_485_in0 = valid ? andOp_483_out : andOp_483_out;
		andOp_485_in1 = valid ? eq_484_out : eq_484_out;
	end
	// controller for andOp_487.andOp_487_in0
	// controller for andOp_487.andOp_487_in1
	// Insensitive connections
	always @(*) begin
		andOp_487_in0 = valid ? andOp_483_out : andOp_483_out;
		andOp_487_in1 = valid ? notOp_486_out : notOp_486_out;
	end
	// controller for andOp_488.andOp_488_in0
	// controller for andOp_488.andOp_488_in1
	// Insensitive connections
	always @(*) begin
		andOp_488_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_488_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_490.andOp_490_in0
	// controller for andOp_490.andOp_490_in1
	// Insensitive connections
	always @(*) begin
		andOp_490_in0 = valid ? andOp_488_out : andOp_488_out;
		andOp_490_in1 = valid ? eq_489_out : eq_489_out;
	end
	// controller for andOp_492.andOp_492_in0
	// controller for andOp_492.andOp_492_in1
	// Insensitive connections
	always @(*) begin
		andOp_492_in0 = valid ? andOp_488_out : andOp_488_out;
		andOp_492_in1 = valid ? notOp_491_out : notOp_491_out;
	end
	// controller for andOp_493.andOp_493_in0
	// controller for andOp_493.andOp_493_in1
	// Insensitive connections
	always @(*) begin
		andOp_493_in0 = valid ? bb_4_active_in_state_4_out_data : bb_4_active_in_state_4_out_data;
		andOp_493_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_495.andOp_495_in0
	// controller for andOp_495.andOp_495_in1
	// Insensitive connections
	always @(*) begin
		andOp_495_in0 = valid ? andOp_493_out : andOp_493_out;
		andOp_495_in1 = valid ? eq_494_out : eq_494_out;
	end
	// controller for andOp_497.andOp_497_in0
	// controller for andOp_497.andOp_497_in1
	// Insensitive connections
	always @(*) begin
		andOp_497_in0 = valid ? andOp_493_out : andOp_493_out;
		andOp_497_in1 = valid ? notOp_496_out : notOp_496_out;
	end
	// controller for andOp_498.andOp_498_in0
	// controller for andOp_498.andOp_498_in1
	// Insensitive connections
	always @(*) begin
		andOp_498_in0 = valid ? 1'd0 : 1'd0;
		andOp_498_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_500.andOp_500_in0
	// controller for andOp_500.andOp_500_in1
	// Insensitive connections
	always @(*) begin
		andOp_500_in0 = valid ? andOp_498_out : andOp_498_out;
		andOp_500_in1 = valid ? eq_499_out : eq_499_out;
	end
	// controller for andOp_502.andOp_502_in0
	// controller for andOp_502.andOp_502_in1
	// Insensitive connections
	always @(*) begin
		andOp_502_in0 = valid ? andOp_498_out : andOp_498_out;
		andOp_502_in1 = valid ? notOp_501_out : notOp_501_out;
	end
	// controller for andOp_503.andOp_503_in0
	// controller for andOp_503.andOp_503_in1
	// Insensitive connections
	always @(*) begin
		andOp_503_in0 = valid ? 1'd0 : 1'd0;
		andOp_503_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_505.andOp_505_in0
	// controller for andOp_505.andOp_505_in1
	// Insensitive connections
	always @(*) begin
		andOp_505_in0 = valid ? andOp_503_out : andOp_503_out;
		andOp_505_in1 = valid ? eq_504_out : eq_504_out;
	end
	// controller for andOp_507.andOp_507_in0
	// controller for andOp_507.andOp_507_in1
	// Insensitive connections
	always @(*) begin
		andOp_507_in0 = valid ? andOp_503_out : andOp_503_out;
		andOp_507_in1 = valid ? notOp_506_out : notOp_506_out;
	end
	// controller for andOp_508.andOp_508_in0
	// controller for andOp_508.andOp_508_in1
	// Insensitive connections
	always @(*) begin
		andOp_508_in0 = valid ? bb_6_active_in_state_4_out_data : bb_6_active_in_state_4_out_data;
		andOp_508_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_510.andOp_510_in0
	// controller for andOp_510.andOp_510_in1
	// Insensitive connections
	always @(*) begin
		andOp_510_in0 = valid ? andOp_508_out : andOp_508_out;
		andOp_510_in1 = valid ? eq_509_out : eq_509_out;
	end
	// controller for andOp_512.andOp_512_in0
	// controller for andOp_512.andOp_512_in1
	// Insensitive connections
	always @(*) begin
		andOp_512_in0 = valid ? andOp_508_out : andOp_508_out;
		andOp_512_in1 = valid ? notOp_511_out : notOp_511_out;
	end
	// controller for andOp_513.andOp_513_in0
	// controller for andOp_513.andOp_513_in1
	// Insensitive connections
	always @(*) begin
		andOp_513_in0 = valid ? bb_7_active_in_state_4_out_data : bb_7_active_in_state_4_out_data;
		andOp_513_in1 = valid ? state_4_is_active : state_4_is_active;
	end
	// controller for andOp_515.andOp_515_in0
	// controller for andOp_515.andOp_515_in1
	// Insensitive connections
	always @(*) begin
		andOp_515_in0 = valid ? andOp_513_out : andOp_513_out;
		andOp_515_in1 = valid ? eq_514_out : eq_514_out;
	end
	// controller for andOp_517.andOp_517_in0
	// controller for andOp_517.andOp_517_in1
	// Insensitive connections
	always @(*) begin
		andOp_517_in0 = valid ? andOp_513_out : andOp_513_out;
		andOp_517_in1 = valid ? notOp_516_out : notOp_516_out;
	end
	// controller for andOp_90.andOp_90_in0
	// controller for andOp_90.andOp_90_in1
	// Insensitive connections
	always @(*) begin
		andOp_90_in0 = valid ? bb_0_active_in_state_1_out_data : bb_0_active_in_state_1_out_data;
		andOp_90_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_91.andOp_91_in0
	// controller for andOp_91.andOp_91_in1
	// Insensitive connections
	always @(*) begin
		andOp_91_in0 = valid ? andOp_90_out : andOp_90_out;
		andOp_91_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_93.andOp_93_in0
	// controller for andOp_93.andOp_93_in1
	// Insensitive connections
	always @(*) begin
		andOp_93_in0 = valid ? bb_3_active_in_state_1_out_data : bb_3_active_in_state_1_out_data;
		andOp_93_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_94.andOp_94_in0
	// controller for andOp_94.andOp_94_in1
	// Insensitive connections
	always @(*) begin
		andOp_94_in0 = valid ? andOp_93_out : andOp_93_out;
		andOp_94_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_96.andOp_96_in0
	// controller for andOp_96.andOp_96_in1
	// Insensitive connections
	always @(*) begin
		andOp_96_in0 = valid ? bb_8_active_in_state_1_out_data : bb_8_active_in_state_1_out_data;
		andOp_96_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for andOp_97.andOp_97_in0
	// controller for andOp_97.andOp_97_in1
	// Insensitive connections
	always @(*) begin
		andOp_97_in0 = valid ? andOp_96_out : andOp_96_out;
		andOp_97_in1 = valid ? 1'd1 : 1'd1;
	end
	// controller for andOp_99.andOp_99_in0
	// controller for andOp_99.andOp_99_in1
	// Insensitive connections
	always @(*) begin
		andOp_99_in0 = valid ? bb_9_active_in_state_1_out_data : bb_9_active_in_state_1_out_data;
		andOp_99_in1 = valid ? state_1_is_active : state_1_is_active;
	end
	// controller for bb_0_active_in_state_0.bb_0_active_in_state_0_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_0_in_data = eq_141_out;
		end else begin
			bb_0_active_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_active_in_state_1.bb_0_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_0_active_in_state_1_in_data = eq_148_out;
		end else begin
			bb_0_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_0.bb_0_predecessor_in_state_0_in_data
	always @(*) begin
		if (eq_164_out) begin 
			bb_0_predecessor_in_state_0_in_data = state_0_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_0_in_data = 0;
		end
	end
	// controller for bb_0_predecessor_in_state_1.bb_0_predecessor_in_state_1_in_data
	always @(*) begin
		if (eq_174_out) begin 
			bb_0_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_0_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_2.bb_10_active_in_state_2_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_2_in_data = eq_149_out;
		end else begin
			bb_10_active_in_state_2_in_data = 0;
		end
	end
	// controller for bb_10_active_in_state_3.bb_10_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_10_active_in_state_3_in_data = eq_150_out;
		end else begin
			bb_10_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_2.bb_10_predecessor_in_state_2_in_data
	always @(*) begin
		if (eq_175_out) begin 
			bb_10_predecessor_in_state_2_in_data = state_2_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_2_in_data = 0;
		end
	end
	// controller for bb_10_predecessor_in_state_3.bb_10_predecessor_in_state_3_in_data
	always @(*) begin
		if (eq_176_out) begin 
			bb_10_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_10_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_1_active_in_state_4.bb_1_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_1_active_in_state_4_in_data = orOp_154_out;
		end else begin
			bb_1_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_1_predecessor_in_state_4.bb_1_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_182_out) begin 
			bb_1_predecessor_in_state_4_in_data = 32'd4;
		end else if (eq_180_out) begin 
			bb_1_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_1_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_active_in_state_4.bb_2_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_2_active_in_state_4_in_data = orOp_163_out;
		end else begin
			bb_2_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_2_predecessor_in_state_4.bb_2_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_195_out) begin 
			bb_2_predecessor_in_state_4_in_data = 32'd7;
		end else if (eq_193_out) begin 
			bb_2_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_2_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_3_active_in_state_1.bb_3_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_3_active_in_state_1_in_data = orOp_143_out;
		end else begin
			bb_3_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_3_predecessor_in_state_1.bb_3_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_167_out) begin 
			bb_3_predecessor_in_state_1_in_data = 32'd0;
		end else if (eq_165_out) begin 
			bb_3_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_3_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_3.bb_4_active_in_state_3_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_3_in_data = orOp_152_out;
		end else begin
			bb_4_active_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_active_in_state_4.bb_4_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_4_active_in_state_4_in_data = eq_161_out;
		end else begin
			bb_4_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_3.bb_4_predecessor_in_state_3_in_data
	always @(*) begin
		if (andOp_179_out) begin 
			bb_4_predecessor_in_state_3_in_data = 32'd10;
		end else if (eq_177_out) begin 
			bb_4_predecessor_in_state_3_in_data = state_3_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_3_in_data = 0;
		end
	end
	// controller for bb_4_predecessor_in_state_4.bb_4_predecessor_in_state_4_in_data
	always @(*) begin
		if (eq_192_out) begin 
			bb_4_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_4_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_5_active_in_state_4.bb_5_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_5_active_in_state_4_in_data = orOp_156_out;
		end else begin
			bb_5_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_5_predecessor_in_state_4.bb_5_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_185_out) begin 
			bb_5_predecessor_in_state_4_in_data = 32'd1;
		end else if (eq_183_out) begin 
			bb_5_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_5_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_6_active_in_state_4.bb_6_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_6_active_in_state_4_in_data = orOp_158_out;
		end else begin
			bb_6_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_6_predecessor_in_state_4.bb_6_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_188_out) begin 
			bb_6_predecessor_in_state_4_in_data = 32'd5;
		end else if (eq_186_out) begin 
			bb_6_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_6_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_7_active_in_state_4.bb_7_active_in_state_4_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_7_active_in_state_4_in_data = orOp_160_out;
		end else begin
			bb_7_active_in_state_4_in_data = 0;
		end
	end
	// controller for bb_7_predecessor_in_state_4.bb_7_predecessor_in_state_4_in_data
	always @(*) begin
		if (andOp_191_out) begin 
			bb_7_predecessor_in_state_4_in_data = 32'd6;
		end else if (eq_189_out) begin 
			bb_7_predecessor_in_state_4_in_data = state_4_last_BB_reg;
		end else begin
			bb_7_predecessor_in_state_4_in_data = 0;
		end
	end
	// controller for bb_8_active_in_state_1.bb_8_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_8_active_in_state_1_in_data = orOp_145_out;
		end else begin
			bb_8_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_8_predecessor_in_state_1.bb_8_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_170_out) begin 
			bb_8_predecessor_in_state_1_in_data = 32'd3;
		end else if (eq_168_out) begin 
			bb_8_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_8_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for bb_9_active_in_state_1.bb_9_active_in_state_1_in_data
	always @(*) begin
		if (1'd1) begin 
			bb_9_active_in_state_1_in_data = orOp_147_out;
		end else begin
			bb_9_active_in_state_1_in_data = 0;
		end
	end
	// controller for bb_9_predecessor_in_state_1.bb_9_predecessor_in_state_1_in_data
	always @(*) begin
		if (andOp_173_out) begin 
			bb_9_predecessor_in_state_1_in_data = 32'd8;
		end else if (eq_171_out) begin 
			bb_9_predecessor_in_state_1_in_data = state_1_last_BB_reg;
		end else begin
			bb_9_predecessor_in_state_1_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_0.br_0_happened_in_state_0_in_data
	always @(*) begin
		if (andOp_91_out) begin 
			br_0_happened_in_state_0_in_data = 1'd1;
		end else if (notOp_92_out) begin 
			br_0_happened_in_state_0_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_0_in_data = 0;
		end
	end
	// controller for br_0_happened_in_state_1.br_0_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_106_out) begin 
			br_0_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_107_out) begin 
			br_0_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_0_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_2.br_10_happened_in_state_2_in_data
	always @(*) begin
		if (andOp_109_out) begin 
			br_10_happened_in_state_2_in_data = 1'd1;
		end else if (notOp_110_out) begin 
			br_10_happened_in_state_2_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_2_in_data = 0;
		end
	end
	// controller for br_10_happened_in_state_3.br_10_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_112_out) begin 
			br_10_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_113_out) begin 
			br_10_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_10_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_1_happened_in_state_4.br_1_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_121_out) begin 
			br_1_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_122_out) begin 
			br_1_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_1_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_3_happened_in_state_1.br_3_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_94_out) begin 
			br_3_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_95_out) begin 
			br_3_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_3_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_3.br_4_happened_in_state_3_in_data
	always @(*) begin
		if (andOp_115_out) begin 
			br_4_happened_in_state_3_in_data = 1'd1;
		end else if (notOp_116_out) begin 
			br_4_happened_in_state_3_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_3_in_data = 0;
		end
	end
	// controller for br_4_happened_in_state_4.br_4_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_136_out) begin 
			br_4_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_137_out) begin 
			br_4_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_4_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_5_happened_in_state_4.br_5_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_124_out) begin 
			br_5_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_125_out) begin 
			br_5_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_5_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_6_happened_in_state_4.br_6_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_127_out) begin 
			br_6_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_128_out) begin 
			br_6_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_6_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_7_happened_in_state_4.br_7_happened_in_state_4_in_data
	always @(*) begin
		if (andOp_133_out) begin 
			br_7_happened_in_state_4_in_data = 1'd1;
		end else if (notOp_134_out) begin 
			br_7_happened_in_state_4_in_data = 1'd0;
		end else begin
			br_7_happened_in_state_4_in_data = 0;
		end
	end
	// controller for br_8_happened_in_state_1.br_8_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_97_out) begin 
			br_8_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_98_out) begin 
			br_8_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_8_happened_in_state_1_in_data = 0;
		end
	end
	// controller for br_9_happened_in_state_1.br_9_happened_in_state_1_in_data
	always @(*) begin
		if (andOp_100_out) begin 
			br_9_happened_in_state_1_in_data = 1'd1;
		end else if (notOp_101_out) begin 
			br_9_happened_in_state_1_in_data = 1'd0;
		end else begin
			br_9_happened_in_state_1_in_data = 0;
		end
	end
	// controller for concat_204.concat_204_in0
	// controller for concat_204.concat_204_in1
	// Insensitive connections
	always @(*) begin
		concat_204_in0 = valid ? data_in_1_25_out_data : data_in_1_25_out_data;
		concat_204_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for concat_205.concat_205_in0
	// controller for concat_205.concat_205_in1
	// Insensitive connections
	always @(*) begin
		concat_205_in0 = valid ? 32'd4 : 32'd4;
		concat_205_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for data_in_0_1.data_in_0_1_in_data
	always @(*) begin
		if (andOp_244_out) begin 
			data_in_0_1_in_data = data_store_0_0;
		end else if (andOp_246_out) begin 
			data_in_0_1_in_data = data_store_1_18;
		end else if (andOp_248_out) begin 
			data_in_0_1_in_data = data_store_2_36;
		end else if (andOp_250_out) begin 
			data_in_0_1_in_data = data_store_3_54;
		end else if (andOp_252_out) begin 
			data_in_0_1_in_data = data_store_4_72;
		end else begin
			data_in_0_1_in_data = 0;
		end
	end
	// controller for data_in_0_11.data_in_0_11_in_data
	always @(*) begin
		if (andOp_244_out) begin 
			data_in_0_11_in_data = data_store_0_10;
		end else if (andOp_246_out) begin 
			data_in_0_11_in_data = data_store_1_28;
		end else if (andOp_248_out) begin 
			data_in_0_11_in_data = data_store_2_46;
		end else if (andOp_250_out) begin 
			data_in_0_11_in_data = data_store_3_64;
		end else if (andOp_252_out) begin 
			data_in_0_11_in_data = data_store_4_82;
		end else begin
			data_in_0_11_in_data = 0;
		end
	end
	// controller for data_in_0_13.data_in_0_13_in_data
	always @(*) begin
		if (andOp_244_out) begin 
			data_in_0_13_in_data = data_store_0_12;
		end else if (andOp_246_out) begin 
			data_in_0_13_in_data = data_store_1_30;
		end else if (andOp_248_out) begin 
			data_in_0_13_in_data = data_store_2_48;
		end else if (andOp_250_out) begin 
			data_in_0_13_in_data = data_store_3_66;
		end else if (andOp_252_out) begin 
			data_in_0_13_in_data = data_store_4_84;
		end else begin
			data_in_0_13_in_data = 0;
		end
	end
	// controller for data_in_0_15.data_in_0_15_in_data
	always @(*) begin
		if (andOp_244_out) begin 
			data_in_0_15_in_data = data_store_0_14;
		end else if (andOp_246_out) begin 
			data_in_0_15_in_data = data_store_1_32;
		end else if (andOp_248_out) begin 
			data_in_0_15_in_data = data_store_2_50;
		end else if (andOp_250_out) begin 
			data_in_0_15_in_data = data_store_3_68;
		end else if (andOp_252_out) begin 
			data_in_0_15_in_data = data_store_4_86;
		end else begin
			data_in_0_15_in_data = 0;
		end
	end
	// controller for data_in_0_17.data_in_0_17_in_data
	always @(*) begin
		if (andOp_244_out) begin 
			data_in_0_17_in_data = data_store_0_16;
		end else if (andOp_246_out) begin 
			data_in_0_17_in_data = data_store_1_34;
		end else if (andOp_248_out) begin 
			data_in_0_17_in_data = data_store_2_52;
		end else if (andOp_250_out) begin 
			data_in_0_17_in_data = data_store_3_70;
		end else if (andOp_252_out) begin 
			data_in_0_17_in_data = data_store_4_88;
		end else begin
			data_in_0_17_in_data = 0;
		end
	end
	// controller for data_in_0_3.data_in_0_3_in_data
	always @(*) begin
		if (andOp_244_out) begin 
			data_in_0_3_in_data = data_store_0_2;
		end else if (andOp_246_out) begin 
			data_in_0_3_in_data = data_store_1_20;
		end else if (andOp_248_out) begin 
			data_in_0_3_in_data = data_store_2_38;
		end else if (andOp_250_out) begin 
			data_in_0_3_in_data = data_store_3_56;
		end else if (andOp_252_out) begin 
			data_in_0_3_in_data = data_store_4_74;
		end else begin
			data_in_0_3_in_data = 0;
		end
	end
	// controller for data_in_0_5.data_in_0_5_in_data
	always @(*) begin
		if (andOp_244_out) begin 
			data_in_0_5_in_data = data_store_0_4;
		end else if (andOp_246_out) begin 
			data_in_0_5_in_data = data_store_1_22;
		end else if (andOp_248_out) begin 
			data_in_0_5_in_data = data_store_2_40;
		end else if (andOp_250_out) begin 
			data_in_0_5_in_data = data_store_3_58;
		end else if (andOp_252_out) begin 
			data_in_0_5_in_data = data_store_4_76;
		end else begin
			data_in_0_5_in_data = 0;
		end
	end
	// controller for data_in_0_7.data_in_0_7_in_data
	always @(*) begin
		if (andOp_244_out) begin 
			data_in_0_7_in_data = data_store_0_6;
		end else if (andOp_246_out) begin 
			data_in_0_7_in_data = data_store_1_24;
		end else if (andOp_248_out) begin 
			data_in_0_7_in_data = data_store_2_42;
		end else if (andOp_250_out) begin 
			data_in_0_7_in_data = data_store_3_60;
		end else if (andOp_252_out) begin 
			data_in_0_7_in_data = data_store_4_78;
		end else begin
			data_in_0_7_in_data = 0;
		end
	end
	// controller for data_in_0_9.data_in_0_9_in_data
	always @(*) begin
		if (andOp_244_out) begin 
			data_in_0_9_in_data = data_store_0_8;
		end else if (andOp_246_out) begin 
			data_in_0_9_in_data = data_store_1_26;
		end else if (andOp_248_out) begin 
			data_in_0_9_in_data = data_store_2_44;
		end else if (andOp_250_out) begin 
			data_in_0_9_in_data = data_store_3_62;
		end else if (andOp_252_out) begin 
			data_in_0_9_in_data = data_store_4_80;
		end else begin
			data_in_0_9_in_data = 0;
		end
	end
	// controller for data_in_1_19.data_in_1_19_in_data
	always @(*) begin
		if (andOp_299_out) begin 
			data_in_1_19_in_data = data_store_0_0;
		end else if (andOp_301_out) begin 
			data_in_1_19_in_data = data_store_1_18;
		end else if (andOp_303_out) begin 
			data_in_1_19_in_data = data_store_2_36;
		end else if (andOp_305_out) begin 
			data_in_1_19_in_data = data_store_3_54;
		end else if (andOp_307_out) begin 
			data_in_1_19_in_data = data_store_4_72;
		end else begin
			data_in_1_19_in_data = 0;
		end
	end
	// controller for data_in_1_21.data_in_1_21_in_data
	always @(*) begin
		if (andOp_299_out) begin 
			data_in_1_21_in_data = data_store_0_2;
		end else if (andOp_301_out) begin 
			data_in_1_21_in_data = data_store_1_20;
		end else if (andOp_303_out) begin 
			data_in_1_21_in_data = data_store_2_38;
		end else if (andOp_305_out) begin 
			data_in_1_21_in_data = data_store_3_56;
		end else if (andOp_307_out) begin 
			data_in_1_21_in_data = data_store_4_74;
		end else begin
			data_in_1_21_in_data = 0;
		end
	end
	// controller for data_in_1_23.data_in_1_23_in_data
	always @(*) begin
		if (andOp_299_out) begin 
			data_in_1_23_in_data = data_store_0_4;
		end else if (andOp_301_out) begin 
			data_in_1_23_in_data = data_store_1_22;
		end else if (andOp_303_out) begin 
			data_in_1_23_in_data = data_store_2_40;
		end else if (andOp_305_out) begin 
			data_in_1_23_in_data = data_store_3_58;
		end else if (andOp_307_out) begin 
			data_in_1_23_in_data = data_store_4_76;
		end else begin
			data_in_1_23_in_data = 0;
		end
	end
	// controller for data_in_1_25.data_in_1_25_in_data
	always @(*) begin
		if (andOp_299_out) begin 
			data_in_1_25_in_data = data_store_0_6;
		end else if (andOp_301_out) begin 
			data_in_1_25_in_data = data_store_1_24;
		end else if (andOp_303_out) begin 
			data_in_1_25_in_data = data_store_2_42;
		end else if (andOp_305_out) begin 
			data_in_1_25_in_data = data_store_3_60;
		end else if (andOp_307_out) begin 
			data_in_1_25_in_data = data_store_4_78;
		end else begin
			data_in_1_25_in_data = 0;
		end
	end
	// controller for data_in_1_27.data_in_1_27_in_data
	always @(*) begin
		if (andOp_299_out) begin 
			data_in_1_27_in_data = data_store_0_8;
		end else if (andOp_301_out) begin 
			data_in_1_27_in_data = data_store_1_26;
		end else if (andOp_303_out) begin 
			data_in_1_27_in_data = data_store_2_44;
		end else if (andOp_305_out) begin 
			data_in_1_27_in_data = data_store_3_62;
		end else if (andOp_307_out) begin 
			data_in_1_27_in_data = data_store_4_80;
		end else begin
			data_in_1_27_in_data = 0;
		end
	end
	// controller for data_in_1_29.data_in_1_29_in_data
	always @(*) begin
		if (andOp_299_out) begin 
			data_in_1_29_in_data = data_store_0_10;
		end else if (andOp_301_out) begin 
			data_in_1_29_in_data = data_store_1_28;
		end else if (andOp_303_out) begin 
			data_in_1_29_in_data = data_store_2_46;
		end else if (andOp_305_out) begin 
			data_in_1_29_in_data = data_store_3_64;
		end else if (andOp_307_out) begin 
			data_in_1_29_in_data = data_store_4_82;
		end else begin
			data_in_1_29_in_data = 0;
		end
	end
	// controller for data_in_1_31.data_in_1_31_in_data
	always @(*) begin
		if (andOp_299_out) begin 
			data_in_1_31_in_data = data_store_0_12;
		end else if (andOp_301_out) begin 
			data_in_1_31_in_data = data_store_1_30;
		end else if (andOp_303_out) begin 
			data_in_1_31_in_data = data_store_2_48;
		end else if (andOp_305_out) begin 
			data_in_1_31_in_data = data_store_3_66;
		end else if (andOp_307_out) begin 
			data_in_1_31_in_data = data_store_4_84;
		end else begin
			data_in_1_31_in_data = 0;
		end
	end
	// controller for data_in_1_33.data_in_1_33_in_data
	always @(*) begin
		if (andOp_299_out) begin 
			data_in_1_33_in_data = data_store_0_14;
		end else if (andOp_301_out) begin 
			data_in_1_33_in_data = data_store_1_32;
		end else if (andOp_303_out) begin 
			data_in_1_33_in_data = data_store_2_50;
		end else if (andOp_305_out) begin 
			data_in_1_33_in_data = data_store_3_68;
		end else if (andOp_307_out) begin 
			data_in_1_33_in_data = data_store_4_86;
		end else begin
			data_in_1_33_in_data = 0;
		end
	end
	// controller for data_in_1_35.data_in_1_35_in_data
	always @(*) begin
		if (andOp_299_out) begin 
			data_in_1_35_in_data = data_store_0_16;
		end else if (andOp_301_out) begin 
			data_in_1_35_in_data = data_store_1_34;
		end else if (andOp_303_out) begin 
			data_in_1_35_in_data = data_store_2_52;
		end else if (andOp_305_out) begin 
			data_in_1_35_in_data = data_store_3_70;
		end else if (andOp_307_out) begin 
			data_in_1_35_in_data = data_store_4_88;
		end else begin
			data_in_1_35_in_data = 0;
		end
	end
	// controller for data_in_2_37.data_in_2_37_in_data
	always @(*) begin
		if (andOp_354_out) begin 
			data_in_2_37_in_data = data_store_0_0;
		end else if (andOp_356_out) begin 
			data_in_2_37_in_data = data_store_1_18;
		end else if (andOp_358_out) begin 
			data_in_2_37_in_data = data_store_2_36;
		end else if (andOp_360_out) begin 
			data_in_2_37_in_data = data_store_3_54;
		end else if (andOp_362_out) begin 
			data_in_2_37_in_data = data_store_4_72;
		end else begin
			data_in_2_37_in_data = 0;
		end
	end
	// controller for data_in_2_39.data_in_2_39_in_data
	always @(*) begin
		if (andOp_354_out) begin 
			data_in_2_39_in_data = data_store_0_2;
		end else if (andOp_356_out) begin 
			data_in_2_39_in_data = data_store_1_20;
		end else if (andOp_358_out) begin 
			data_in_2_39_in_data = data_store_2_38;
		end else if (andOp_360_out) begin 
			data_in_2_39_in_data = data_store_3_56;
		end else if (andOp_362_out) begin 
			data_in_2_39_in_data = data_store_4_74;
		end else begin
			data_in_2_39_in_data = 0;
		end
	end
	// controller for data_in_2_41.data_in_2_41_in_data
	always @(*) begin
		if (andOp_354_out) begin 
			data_in_2_41_in_data = data_store_0_4;
		end else if (andOp_356_out) begin 
			data_in_2_41_in_data = data_store_1_22;
		end else if (andOp_358_out) begin 
			data_in_2_41_in_data = data_store_2_40;
		end else if (andOp_360_out) begin 
			data_in_2_41_in_data = data_store_3_58;
		end else if (andOp_362_out) begin 
			data_in_2_41_in_data = data_store_4_76;
		end else begin
			data_in_2_41_in_data = 0;
		end
	end
	// controller for data_in_2_43.data_in_2_43_in_data
	always @(*) begin
		if (andOp_354_out) begin 
			data_in_2_43_in_data = data_store_0_6;
		end else if (andOp_356_out) begin 
			data_in_2_43_in_data = data_store_1_24;
		end else if (andOp_358_out) begin 
			data_in_2_43_in_data = data_store_2_42;
		end else if (andOp_360_out) begin 
			data_in_2_43_in_data = data_store_3_60;
		end else if (andOp_362_out) begin 
			data_in_2_43_in_data = data_store_4_78;
		end else begin
			data_in_2_43_in_data = 0;
		end
	end
	// controller for data_in_2_45.data_in_2_45_in_data
	always @(*) begin
		if (andOp_354_out) begin 
			data_in_2_45_in_data = data_store_0_8;
		end else if (andOp_356_out) begin 
			data_in_2_45_in_data = data_store_1_26;
		end else if (andOp_358_out) begin 
			data_in_2_45_in_data = data_store_2_44;
		end else if (andOp_360_out) begin 
			data_in_2_45_in_data = data_store_3_62;
		end else if (andOp_362_out) begin 
			data_in_2_45_in_data = data_store_4_80;
		end else begin
			data_in_2_45_in_data = 0;
		end
	end
	// controller for data_in_2_47.data_in_2_47_in_data
	always @(*) begin
		if (andOp_354_out) begin 
			data_in_2_47_in_data = data_store_0_10;
		end else if (andOp_356_out) begin 
			data_in_2_47_in_data = data_store_1_28;
		end else if (andOp_358_out) begin 
			data_in_2_47_in_data = data_store_2_46;
		end else if (andOp_360_out) begin 
			data_in_2_47_in_data = data_store_3_64;
		end else if (andOp_362_out) begin 
			data_in_2_47_in_data = data_store_4_82;
		end else begin
			data_in_2_47_in_data = 0;
		end
	end
	// controller for data_in_2_49.data_in_2_49_in_data
	always @(*) begin
		if (andOp_354_out) begin 
			data_in_2_49_in_data = data_store_0_12;
		end else if (andOp_356_out) begin 
			data_in_2_49_in_data = data_store_1_30;
		end else if (andOp_358_out) begin 
			data_in_2_49_in_data = data_store_2_48;
		end else if (andOp_360_out) begin 
			data_in_2_49_in_data = data_store_3_66;
		end else if (andOp_362_out) begin 
			data_in_2_49_in_data = data_store_4_84;
		end else begin
			data_in_2_49_in_data = 0;
		end
	end
	// controller for data_in_2_51.data_in_2_51_in_data
	always @(*) begin
		if (andOp_354_out) begin 
			data_in_2_51_in_data = data_store_0_14;
		end else if (andOp_356_out) begin 
			data_in_2_51_in_data = data_store_1_32;
		end else if (andOp_358_out) begin 
			data_in_2_51_in_data = data_store_2_50;
		end else if (andOp_360_out) begin 
			data_in_2_51_in_data = data_store_3_68;
		end else if (andOp_362_out) begin 
			data_in_2_51_in_data = data_store_4_86;
		end else begin
			data_in_2_51_in_data = 0;
		end
	end
	// controller for data_in_2_53.data_in_2_53_in_data
	always @(*) begin
		if (andOp_354_out) begin 
			data_in_2_53_in_data = data_store_0_16;
		end else if (andOp_356_out) begin 
			data_in_2_53_in_data = data_store_1_34;
		end else if (andOp_358_out) begin 
			data_in_2_53_in_data = data_store_2_52;
		end else if (andOp_360_out) begin 
			data_in_2_53_in_data = data_store_3_70;
		end else if (andOp_362_out) begin 
			data_in_2_53_in_data = data_store_4_88;
		end else begin
			data_in_2_53_in_data = 0;
		end
	end
	// controller for data_in_3_55.data_in_3_55_in_data
	always @(*) begin
		if (andOp_409_out) begin 
			data_in_3_55_in_data = data_store_0_0;
		end else if (andOp_411_out) begin 
			data_in_3_55_in_data = data_store_1_18;
		end else if (andOp_413_out) begin 
			data_in_3_55_in_data = data_store_2_36;
		end else if (andOp_415_out) begin 
			data_in_3_55_in_data = data_store_3_54;
		end else if (andOp_417_out) begin 
			data_in_3_55_in_data = data_store_4_72;
		end else begin
			data_in_3_55_in_data = 0;
		end
	end
	// controller for data_in_3_57.data_in_3_57_in_data
	always @(*) begin
		if (andOp_409_out) begin 
			data_in_3_57_in_data = data_store_0_2;
		end else if (andOp_411_out) begin 
			data_in_3_57_in_data = data_store_1_20;
		end else if (andOp_413_out) begin 
			data_in_3_57_in_data = data_store_2_38;
		end else if (andOp_415_out) begin 
			data_in_3_57_in_data = data_store_3_56;
		end else if (andOp_417_out) begin 
			data_in_3_57_in_data = data_store_4_74;
		end else begin
			data_in_3_57_in_data = 0;
		end
	end
	// controller for data_in_3_59.data_in_3_59_in_data
	always @(*) begin
		if (andOp_409_out) begin 
			data_in_3_59_in_data = data_store_0_4;
		end else if (andOp_411_out) begin 
			data_in_3_59_in_data = data_store_1_22;
		end else if (andOp_413_out) begin 
			data_in_3_59_in_data = data_store_2_40;
		end else if (andOp_415_out) begin 
			data_in_3_59_in_data = data_store_3_58;
		end else if (andOp_417_out) begin 
			data_in_3_59_in_data = data_store_4_76;
		end else begin
			data_in_3_59_in_data = 0;
		end
	end
	// controller for data_in_3_61.data_in_3_61_in_data
	always @(*) begin
		if (andOp_409_out) begin 
			data_in_3_61_in_data = data_store_0_6;
		end else if (andOp_411_out) begin 
			data_in_3_61_in_data = data_store_1_24;
		end else if (andOp_413_out) begin 
			data_in_3_61_in_data = data_store_2_42;
		end else if (andOp_415_out) begin 
			data_in_3_61_in_data = data_store_3_60;
		end else if (andOp_417_out) begin 
			data_in_3_61_in_data = data_store_4_78;
		end else begin
			data_in_3_61_in_data = 0;
		end
	end
	// controller for data_in_3_63.data_in_3_63_in_data
	always @(*) begin
		if (andOp_409_out) begin 
			data_in_3_63_in_data = data_store_0_8;
		end else if (andOp_411_out) begin 
			data_in_3_63_in_data = data_store_1_26;
		end else if (andOp_413_out) begin 
			data_in_3_63_in_data = data_store_2_44;
		end else if (andOp_415_out) begin 
			data_in_3_63_in_data = data_store_3_62;
		end else if (andOp_417_out) begin 
			data_in_3_63_in_data = data_store_4_80;
		end else begin
			data_in_3_63_in_data = 0;
		end
	end
	// controller for data_in_3_65.data_in_3_65_in_data
	always @(*) begin
		if (andOp_409_out) begin 
			data_in_3_65_in_data = data_store_0_10;
		end else if (andOp_411_out) begin 
			data_in_3_65_in_data = data_store_1_28;
		end else if (andOp_413_out) begin 
			data_in_3_65_in_data = data_store_2_46;
		end else if (andOp_415_out) begin 
			data_in_3_65_in_data = data_store_3_64;
		end else if (andOp_417_out) begin 
			data_in_3_65_in_data = data_store_4_82;
		end else begin
			data_in_3_65_in_data = 0;
		end
	end
	// controller for data_in_3_67.data_in_3_67_in_data
	always @(*) begin
		if (andOp_409_out) begin 
			data_in_3_67_in_data = data_store_0_12;
		end else if (andOp_411_out) begin 
			data_in_3_67_in_data = data_store_1_30;
		end else if (andOp_413_out) begin 
			data_in_3_67_in_data = data_store_2_48;
		end else if (andOp_415_out) begin 
			data_in_3_67_in_data = data_store_3_66;
		end else if (andOp_417_out) begin 
			data_in_3_67_in_data = data_store_4_84;
		end else begin
			data_in_3_67_in_data = 0;
		end
	end
	// controller for data_in_3_69.data_in_3_69_in_data
	always @(*) begin
		if (andOp_409_out) begin 
			data_in_3_69_in_data = data_store_0_14;
		end else if (andOp_411_out) begin 
			data_in_3_69_in_data = data_store_1_32;
		end else if (andOp_413_out) begin 
			data_in_3_69_in_data = data_store_2_50;
		end else if (andOp_415_out) begin 
			data_in_3_69_in_data = data_store_3_68;
		end else if (andOp_417_out) begin 
			data_in_3_69_in_data = data_store_4_86;
		end else begin
			data_in_3_69_in_data = 0;
		end
	end
	// controller for data_in_3_71.data_in_3_71_in_data
	always @(*) begin
		if (andOp_409_out) begin 
			data_in_3_71_in_data = data_store_0_16;
		end else if (andOp_411_out) begin 
			data_in_3_71_in_data = data_store_1_34;
		end else if (andOp_413_out) begin 
			data_in_3_71_in_data = data_store_2_52;
		end else if (andOp_415_out) begin 
			data_in_3_71_in_data = data_store_3_70;
		end else if (andOp_417_out) begin 
			data_in_3_71_in_data = data_store_4_88;
		end else begin
			data_in_3_71_in_data = 0;
		end
	end
	// controller for data_in_4_73.data_in_4_73_in_data
	always @(*) begin
		if (andOp_464_out) begin 
			data_in_4_73_in_data = data_store_0_0;
		end else if (andOp_466_out) begin 
			data_in_4_73_in_data = data_store_1_18;
		end else if (andOp_468_out) begin 
			data_in_4_73_in_data = data_store_2_36;
		end else if (andOp_470_out) begin 
			data_in_4_73_in_data = data_store_3_54;
		end else if (andOp_472_out) begin 
			data_in_4_73_in_data = data_store_4_72;
		end else begin
			data_in_4_73_in_data = 0;
		end
	end
	// controller for data_in_4_75.data_in_4_75_in_data
	always @(*) begin
		if (andOp_464_out) begin 
			data_in_4_75_in_data = data_store_0_2;
		end else if (andOp_466_out) begin 
			data_in_4_75_in_data = data_store_1_20;
		end else if (andOp_468_out) begin 
			data_in_4_75_in_data = data_store_2_38;
		end else if (andOp_470_out) begin 
			data_in_4_75_in_data = data_store_3_56;
		end else if (andOp_472_out) begin 
			data_in_4_75_in_data = data_store_4_74;
		end else begin
			data_in_4_75_in_data = 0;
		end
	end
	// controller for data_in_4_77.data_in_4_77_in_data
	always @(*) begin
		if (andOp_464_out) begin 
			data_in_4_77_in_data = data_store_0_4;
		end else if (andOp_466_out) begin 
			data_in_4_77_in_data = data_store_1_22;
		end else if (andOp_468_out) begin 
			data_in_4_77_in_data = data_store_2_40;
		end else if (andOp_470_out) begin 
			data_in_4_77_in_data = data_store_3_58;
		end else if (andOp_472_out) begin 
			data_in_4_77_in_data = data_store_4_76;
		end else begin
			data_in_4_77_in_data = 0;
		end
	end
	// controller for data_in_4_79.data_in_4_79_in_data
	always @(*) begin
		if (andOp_464_out) begin 
			data_in_4_79_in_data = data_store_0_6;
		end else if (andOp_466_out) begin 
			data_in_4_79_in_data = data_store_1_24;
		end else if (andOp_468_out) begin 
			data_in_4_79_in_data = data_store_2_42;
		end else if (andOp_470_out) begin 
			data_in_4_79_in_data = data_store_3_60;
		end else if (andOp_472_out) begin 
			data_in_4_79_in_data = data_store_4_78;
		end else begin
			data_in_4_79_in_data = 0;
		end
	end
	// controller for data_in_4_81.data_in_4_81_in_data
	always @(*) begin
		if (andOp_464_out) begin 
			data_in_4_81_in_data = data_store_0_8;
		end else if (andOp_466_out) begin 
			data_in_4_81_in_data = data_store_1_26;
		end else if (andOp_468_out) begin 
			data_in_4_81_in_data = data_store_2_44;
		end else if (andOp_470_out) begin 
			data_in_4_81_in_data = data_store_3_62;
		end else if (andOp_472_out) begin 
			data_in_4_81_in_data = data_store_4_80;
		end else begin
			data_in_4_81_in_data = 0;
		end
	end
	// controller for data_in_4_83.data_in_4_83_in_data
	always @(*) begin
		if (andOp_464_out) begin 
			data_in_4_83_in_data = data_store_0_10;
		end else if (andOp_466_out) begin 
			data_in_4_83_in_data = data_store_1_28;
		end else if (andOp_468_out) begin 
			data_in_4_83_in_data = data_store_2_46;
		end else if (andOp_470_out) begin 
			data_in_4_83_in_data = data_store_3_64;
		end else if (andOp_472_out) begin 
			data_in_4_83_in_data = data_store_4_82;
		end else begin
			data_in_4_83_in_data = 0;
		end
	end
	// controller for data_in_4_85.data_in_4_85_in_data
	always @(*) begin
		if (andOp_464_out) begin 
			data_in_4_85_in_data = data_store_0_12;
		end else if (andOp_466_out) begin 
			data_in_4_85_in_data = data_store_1_30;
		end else if (andOp_468_out) begin 
			data_in_4_85_in_data = data_store_2_48;
		end else if (andOp_470_out) begin 
			data_in_4_85_in_data = data_store_3_66;
		end else if (andOp_472_out) begin 
			data_in_4_85_in_data = data_store_4_84;
		end else begin
			data_in_4_85_in_data = 0;
		end
	end
	// controller for data_in_4_87.data_in_4_87_in_data
	always @(*) begin
		if (andOp_464_out) begin 
			data_in_4_87_in_data = data_store_0_14;
		end else if (andOp_466_out) begin 
			data_in_4_87_in_data = data_store_1_32;
		end else if (andOp_468_out) begin 
			data_in_4_87_in_data = data_store_2_50;
		end else if (andOp_470_out) begin 
			data_in_4_87_in_data = data_store_3_68;
		end else if (andOp_472_out) begin 
			data_in_4_87_in_data = data_store_4_86;
		end else begin
			data_in_4_87_in_data = 0;
		end
	end
	// controller for data_in_4_89.data_in_4_89_in_data
	always @(*) begin
		if (andOp_464_out) begin 
			data_in_4_89_in_data = data_store_0_16;
		end else if (andOp_466_out) begin 
			data_in_4_89_in_data = data_store_1_34;
		end else if (andOp_468_out) begin 
			data_in_4_89_in_data = data_store_2_52;
		end else if (andOp_470_out) begin 
			data_in_4_89_in_data = data_store_3_70;
		end else if (andOp_472_out) begin 
			data_in_4_89_in_data = data_store_4_88;
		end else begin
			data_in_4_89_in_data = 0;
		end
	end
	// controller for eq_141.eq_141_in0
	// controller for eq_141.eq_141_in1
	// Insensitive connections
	always @(*) begin
		eq_141_in0 = valid ? 32'd0 : 32'd0;
		eq_141_in1 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
	end
	// controller for eq_142.eq_142_in0
	// controller for eq_142.eq_142_in1
	// Insensitive connections
	always @(*) begin
		eq_142_in0 = valid ? 32'd3 : 32'd3;
		eq_142_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_144.eq_144_in0
	// controller for eq_144.eq_144_in1
	// Insensitive connections
	always @(*) begin
		eq_144_in0 = valid ? 32'd8 : 32'd8;
		eq_144_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_146.eq_146_in0
	// controller for eq_146.eq_146_in1
	// Insensitive connections
	always @(*) begin
		eq_146_in0 = valid ? 32'd9 : 32'd9;
		eq_146_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_148.eq_148_in0
	// controller for eq_148.eq_148_in1
	// Insensitive connections
	always @(*) begin
		eq_148_in0 = valid ? 32'd0 : 32'd0;
		eq_148_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_149.eq_149_in0
	// controller for eq_149.eq_149_in1
	// Insensitive connections
	always @(*) begin
		eq_149_in0 = valid ? 32'd10 : 32'd10;
		eq_149_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_150.eq_150_in0
	// controller for eq_150.eq_150_in1
	// Insensitive connections
	always @(*) begin
		eq_150_in0 = valid ? 32'd10 : 32'd10;
		eq_150_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_151.eq_151_in0
	// controller for eq_151.eq_151_in1
	// Insensitive connections
	always @(*) begin
		eq_151_in0 = valid ? 32'd4 : 32'd4;
		eq_151_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_153.eq_153_in0
	// controller for eq_153.eq_153_in1
	// Insensitive connections
	always @(*) begin
		eq_153_in0 = valid ? 32'd1 : 32'd1;
		eq_153_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_155.eq_155_in0
	// controller for eq_155.eq_155_in1
	// Insensitive connections
	always @(*) begin
		eq_155_in0 = valid ? 32'd5 : 32'd5;
		eq_155_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_157.eq_157_in0
	// controller for eq_157.eq_157_in1
	// Insensitive connections
	always @(*) begin
		eq_157_in0 = valid ? 32'd6 : 32'd6;
		eq_157_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_159.eq_159_in0
	// controller for eq_159.eq_159_in1
	// Insensitive connections
	always @(*) begin
		eq_159_in0 = valid ? 32'd7 : 32'd7;
		eq_159_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_161.eq_161_in0
	// controller for eq_161.eq_161_in1
	// Insensitive connections
	always @(*) begin
		eq_161_in0 = valid ? 32'd4 : 32'd4;
		eq_161_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_162.eq_162_in0
	// controller for eq_162.eq_162_in1
	// Insensitive connections
	always @(*) begin
		eq_162_in0 = valid ? 32'd2 : 32'd2;
		eq_162_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_164.eq_164_in0
	// controller for eq_164.eq_164_in1
	// Insensitive connections
	always @(*) begin
		eq_164_in0 = valid ? 32'd0 : 32'd0;
		eq_164_in1 = valid ? state_0_entry_BB_reg : state_0_entry_BB_reg;
	end
	// controller for eq_165.eq_165_in0
	// controller for eq_165.eq_165_in1
	// Insensitive connections
	always @(*) begin
		eq_165_in0 = valid ? 32'd3 : 32'd3;
		eq_165_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_168.eq_168_in0
	// controller for eq_168.eq_168_in1
	// Insensitive connections
	always @(*) begin
		eq_168_in0 = valid ? 32'd8 : 32'd8;
		eq_168_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_171.eq_171_in0
	// controller for eq_171.eq_171_in1
	// Insensitive connections
	always @(*) begin
		eq_171_in0 = valid ? 32'd9 : 32'd9;
		eq_171_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_174.eq_174_in0
	// controller for eq_174.eq_174_in1
	// Insensitive connections
	always @(*) begin
		eq_174_in0 = valid ? 32'd0 : 32'd0;
		eq_174_in1 = valid ? state_1_entry_BB_reg : state_1_entry_BB_reg;
	end
	// controller for eq_175.eq_175_in0
	// controller for eq_175.eq_175_in1
	// Insensitive connections
	always @(*) begin
		eq_175_in0 = valid ? 32'd10 : 32'd10;
		eq_175_in1 = valid ? state_2_entry_BB_reg : state_2_entry_BB_reg;
	end
	// controller for eq_176.eq_176_in0
	// controller for eq_176.eq_176_in1
	// Insensitive connections
	always @(*) begin
		eq_176_in0 = valid ? 32'd10 : 32'd10;
		eq_176_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_177.eq_177_in0
	// controller for eq_177.eq_177_in1
	// Insensitive connections
	always @(*) begin
		eq_177_in0 = valid ? 32'd4 : 32'd4;
		eq_177_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_180.eq_180_in0
	// controller for eq_180.eq_180_in1
	// Insensitive connections
	always @(*) begin
		eq_180_in0 = valid ? 32'd1 : 32'd1;
		eq_180_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_183.eq_183_in0
	// controller for eq_183.eq_183_in1
	// Insensitive connections
	always @(*) begin
		eq_183_in0 = valid ? 32'd5 : 32'd5;
		eq_183_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_186.eq_186_in0
	// controller for eq_186.eq_186_in1
	// Insensitive connections
	always @(*) begin
		eq_186_in0 = valid ? 32'd6 : 32'd6;
		eq_186_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_189.eq_189_in0
	// controller for eq_189.eq_189_in1
	// Insensitive connections
	always @(*) begin
		eq_189_in0 = valid ? 32'd7 : 32'd7;
		eq_189_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_192.eq_192_in0
	// controller for eq_192.eq_192_in1
	// Insensitive connections
	always @(*) begin
		eq_192_in0 = valid ? 32'd4 : 32'd4;
		eq_192_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_193.eq_193_in0
	// controller for eq_193.eq_193_in1
	// Insensitive connections
	always @(*) begin
		eq_193_in0 = valid ? 32'd2 : 32'd2;
		eq_193_in1 = valid ? state_4_entry_BB_reg : state_4_entry_BB_reg;
	end
	// controller for eq_211.eq_211_in0
	// controller for eq_211.eq_211_in1
	// Insensitive connections
	always @(*) begin
		eq_211_in0 = valid ? 32'd10 : 32'd10;
		eq_211_in1 = valid ? state_3_entry_BB_reg : state_3_entry_BB_reg;
	end
	// controller for eq_243.eq_243_in0
	// controller for eq_243.eq_243_in1
	// Insensitive connections
	always @(*) begin
		eq_243_in0 = valid ? 32'd0 : 32'd0;
		eq_243_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_245.eq_245_in0
	// controller for eq_245.eq_245_in1
	// Insensitive connections
	always @(*) begin
		eq_245_in0 = valid ? 32'd1 : 32'd1;
		eq_245_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_247.eq_247_in0
	// controller for eq_247.eq_247_in1
	// Insensitive connections
	always @(*) begin
		eq_247_in0 = valid ? 32'd2 : 32'd2;
		eq_247_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_249.eq_249_in0
	// controller for eq_249.eq_249_in1
	// Insensitive connections
	always @(*) begin
		eq_249_in0 = valid ? 32'd3 : 32'd3;
		eq_249_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_251.eq_251_in0
	// controller for eq_251.eq_251_in1
	// Insensitive connections
	always @(*) begin
		eq_251_in0 = valid ? 32'd4 : 32'd4;
		eq_251_in1 = valid ? state_0_last_state : state_0_last_state;
	end
	// controller for eq_254.eq_254_in0
	// controller for eq_254.eq_254_in1
	// Insensitive connections
	always @(*) begin
		eq_254_in0 = valid ? 32'd1 : 32'd1;
		eq_254_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_259.eq_259_in0
	// controller for eq_259.eq_259_in1
	// Insensitive connections
	always @(*) begin
		eq_259_in0 = valid ? 32'd3 : 32'd3;
		eq_259_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_264.eq_264_in0
	// controller for eq_264.eq_264_in1
	// Insensitive connections
	always @(*) begin
		eq_264_in0 = valid ? 32'd3 : 32'd3;
		eq_264_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_269.eq_269_in0
	// controller for eq_269.eq_269_in1
	// Insensitive connections
	always @(*) begin
		eq_269_in0 = valid ? 32'd3 : 32'd3;
		eq_269_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_274.eq_274_in0
	// controller for eq_274.eq_274_in1
	// Insensitive connections
	always @(*) begin
		eq_274_in0 = valid ? 32'd3 : 32'd3;
		eq_274_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_279.eq_279_in0
	// controller for eq_279.eq_279_in1
	// Insensitive connections
	always @(*) begin
		eq_279_in0 = valid ? 32'd1 : 32'd1;
		eq_279_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_284.eq_284_in0
	// controller for eq_284.eq_284_in1
	// Insensitive connections
	always @(*) begin
		eq_284_in0 = valid ? 32'd3 : 32'd3;
		eq_284_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_289.eq_289_in0
	// controller for eq_289.eq_289_in1
	// Insensitive connections
	always @(*) begin
		eq_289_in0 = valid ? 32'd4 : 32'd4;
		eq_289_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_294.eq_294_in0
	// controller for eq_294.eq_294_in1
	// Insensitive connections
	always @(*) begin
		eq_294_in0 = valid ? 32'd4 : 32'd4;
		eq_294_in1 = valid ? 32'd0 : 32'd0;
	end
	// controller for eq_298.eq_298_in0
	// controller for eq_298.eq_298_in1
	// Insensitive connections
	always @(*) begin
		eq_298_in0 = valid ? 32'd0 : 32'd0;
		eq_298_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_300.eq_300_in0
	// controller for eq_300.eq_300_in1
	// Insensitive connections
	always @(*) begin
		eq_300_in0 = valid ? 32'd1 : 32'd1;
		eq_300_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_302.eq_302_in0
	// controller for eq_302.eq_302_in1
	// Insensitive connections
	always @(*) begin
		eq_302_in0 = valid ? 32'd2 : 32'd2;
		eq_302_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_304.eq_304_in0
	// controller for eq_304.eq_304_in1
	// Insensitive connections
	always @(*) begin
		eq_304_in0 = valid ? 32'd3 : 32'd3;
		eq_304_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_306.eq_306_in0
	// controller for eq_306.eq_306_in1
	// Insensitive connections
	always @(*) begin
		eq_306_in0 = valid ? 32'd4 : 32'd4;
		eq_306_in1 = valid ? state_1_last_state : state_1_last_state;
	end
	// controller for eq_309.eq_309_in0
	// controller for eq_309.eq_309_in1
	// Insensitive connections
	always @(*) begin
		eq_309_in0 = valid ? 32'd1 : 32'd1;
		eq_309_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_314.eq_314_in0
	// controller for eq_314.eq_314_in1
	// Insensitive connections
	always @(*) begin
		eq_314_in0 = valid ? 32'd3 : 32'd3;
		eq_314_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_319.eq_319_in0
	// controller for eq_319.eq_319_in1
	// Insensitive connections
	always @(*) begin
		eq_319_in0 = valid ? 32'd3 : 32'd3;
		eq_319_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_324.eq_324_in0
	// controller for eq_324.eq_324_in1
	// Insensitive connections
	always @(*) begin
		eq_324_in0 = valid ? 32'd3 : 32'd3;
		eq_324_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_329.eq_329_in0
	// controller for eq_329.eq_329_in1
	// Insensitive connections
	always @(*) begin
		eq_329_in0 = valid ? 32'd3 : 32'd3;
		eq_329_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_334.eq_334_in0
	// controller for eq_334.eq_334_in1
	// Insensitive connections
	always @(*) begin
		eq_334_in0 = valid ? 32'd1 : 32'd1;
		eq_334_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_339.eq_339_in0
	// controller for eq_339.eq_339_in1
	// Insensitive connections
	always @(*) begin
		eq_339_in0 = valid ? 32'd3 : 32'd3;
		eq_339_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_344.eq_344_in0
	// controller for eq_344.eq_344_in1
	// Insensitive connections
	always @(*) begin
		eq_344_in0 = valid ? 32'd4 : 32'd4;
		eq_344_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_349.eq_349_in0
	// controller for eq_349.eq_349_in1
	// Insensitive connections
	always @(*) begin
		eq_349_in0 = valid ? 32'd4 : 32'd4;
		eq_349_in1 = valid ? 32'd1 : 32'd1;
	end
	// controller for eq_353.eq_353_in0
	// controller for eq_353.eq_353_in1
	// Insensitive connections
	always @(*) begin
		eq_353_in0 = valid ? 32'd0 : 32'd0;
		eq_353_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_355.eq_355_in0
	// controller for eq_355.eq_355_in1
	// Insensitive connections
	always @(*) begin
		eq_355_in0 = valid ? 32'd1 : 32'd1;
		eq_355_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_357.eq_357_in0
	// controller for eq_357.eq_357_in1
	// Insensitive connections
	always @(*) begin
		eq_357_in0 = valid ? 32'd2 : 32'd2;
		eq_357_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_359.eq_359_in0
	// controller for eq_359.eq_359_in1
	// Insensitive connections
	always @(*) begin
		eq_359_in0 = valid ? 32'd3 : 32'd3;
		eq_359_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_361.eq_361_in0
	// controller for eq_361.eq_361_in1
	// Insensitive connections
	always @(*) begin
		eq_361_in0 = valid ? 32'd4 : 32'd4;
		eq_361_in1 = valid ? state_2_last_state : state_2_last_state;
	end
	// controller for eq_364.eq_364_in0
	// controller for eq_364.eq_364_in1
	// Insensitive connections
	always @(*) begin
		eq_364_in0 = valid ? 32'd1 : 32'd1;
		eq_364_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_369.eq_369_in0
	// controller for eq_369.eq_369_in1
	// Insensitive connections
	always @(*) begin
		eq_369_in0 = valid ? 32'd3 : 32'd3;
		eq_369_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_374.eq_374_in0
	// controller for eq_374.eq_374_in1
	// Insensitive connections
	always @(*) begin
		eq_374_in0 = valid ? 32'd3 : 32'd3;
		eq_374_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_379.eq_379_in0
	// controller for eq_379.eq_379_in1
	// Insensitive connections
	always @(*) begin
		eq_379_in0 = valid ? 32'd3 : 32'd3;
		eq_379_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_384.eq_384_in0
	// controller for eq_384.eq_384_in1
	// Insensitive connections
	always @(*) begin
		eq_384_in0 = valid ? 32'd3 : 32'd3;
		eq_384_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_389.eq_389_in0
	// controller for eq_389.eq_389_in1
	// Insensitive connections
	always @(*) begin
		eq_389_in0 = valid ? 32'd1 : 32'd1;
		eq_389_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_394.eq_394_in0
	// controller for eq_394.eq_394_in1
	// Insensitive connections
	always @(*) begin
		eq_394_in0 = valid ? 32'd3 : 32'd3;
		eq_394_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_399.eq_399_in0
	// controller for eq_399.eq_399_in1
	// Insensitive connections
	always @(*) begin
		eq_399_in0 = valid ? 32'd4 : 32'd4;
		eq_399_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_404.eq_404_in0
	// controller for eq_404.eq_404_in1
	// Insensitive connections
	always @(*) begin
		eq_404_in0 = valid ? 32'd4 : 32'd4;
		eq_404_in1 = valid ? 32'd2 : 32'd2;
	end
	// controller for eq_408.eq_408_in0
	// controller for eq_408.eq_408_in1
	// Insensitive connections
	always @(*) begin
		eq_408_in0 = valid ? 32'd0 : 32'd0;
		eq_408_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_410.eq_410_in0
	// controller for eq_410.eq_410_in1
	// Insensitive connections
	always @(*) begin
		eq_410_in0 = valid ? 32'd1 : 32'd1;
		eq_410_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_412.eq_412_in0
	// controller for eq_412.eq_412_in1
	// Insensitive connections
	always @(*) begin
		eq_412_in0 = valid ? 32'd2 : 32'd2;
		eq_412_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_414.eq_414_in0
	// controller for eq_414.eq_414_in1
	// Insensitive connections
	always @(*) begin
		eq_414_in0 = valid ? 32'd3 : 32'd3;
		eq_414_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_416.eq_416_in0
	// controller for eq_416.eq_416_in1
	// Insensitive connections
	always @(*) begin
		eq_416_in0 = valid ? 32'd4 : 32'd4;
		eq_416_in1 = valid ? state_3_last_state : state_3_last_state;
	end
	// controller for eq_419.eq_419_in0
	// controller for eq_419.eq_419_in1
	// Insensitive connections
	always @(*) begin
		eq_419_in0 = valid ? 32'd1 : 32'd1;
		eq_419_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_424.eq_424_in0
	// controller for eq_424.eq_424_in1
	// Insensitive connections
	always @(*) begin
		eq_424_in0 = valid ? 32'd3 : 32'd3;
		eq_424_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_429.eq_429_in0
	// controller for eq_429.eq_429_in1
	// Insensitive connections
	always @(*) begin
		eq_429_in0 = valid ? 32'd3 : 32'd3;
		eq_429_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_434.eq_434_in0
	// controller for eq_434.eq_434_in1
	// Insensitive connections
	always @(*) begin
		eq_434_in0 = valid ? 32'd3 : 32'd3;
		eq_434_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_439.eq_439_in0
	// controller for eq_439.eq_439_in1
	// Insensitive connections
	always @(*) begin
		eq_439_in0 = valid ? 32'd3 : 32'd3;
		eq_439_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_444.eq_444_in0
	// controller for eq_444.eq_444_in1
	// Insensitive connections
	always @(*) begin
		eq_444_in0 = valid ? 32'd1 : 32'd1;
		eq_444_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_449.eq_449_in0
	// controller for eq_449.eq_449_in1
	// Insensitive connections
	always @(*) begin
		eq_449_in0 = valid ? 32'd3 : 32'd3;
		eq_449_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_454.eq_454_in0
	// controller for eq_454.eq_454_in1
	// Insensitive connections
	always @(*) begin
		eq_454_in0 = valid ? 32'd4 : 32'd4;
		eq_454_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_459.eq_459_in0
	// controller for eq_459.eq_459_in1
	// Insensitive connections
	always @(*) begin
		eq_459_in0 = valid ? 32'd4 : 32'd4;
		eq_459_in1 = valid ? 32'd3 : 32'd3;
	end
	// controller for eq_463.eq_463_in0
	// controller for eq_463.eq_463_in1
	// Insensitive connections
	always @(*) begin
		eq_463_in0 = valid ? 32'd0 : 32'd0;
		eq_463_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_465.eq_465_in0
	// controller for eq_465.eq_465_in1
	// Insensitive connections
	always @(*) begin
		eq_465_in0 = valid ? 32'd1 : 32'd1;
		eq_465_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_467.eq_467_in0
	// controller for eq_467.eq_467_in1
	// Insensitive connections
	always @(*) begin
		eq_467_in0 = valid ? 32'd2 : 32'd2;
		eq_467_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_469.eq_469_in0
	// controller for eq_469.eq_469_in1
	// Insensitive connections
	always @(*) begin
		eq_469_in0 = valid ? 32'd3 : 32'd3;
		eq_469_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_471.eq_471_in0
	// controller for eq_471.eq_471_in1
	// Insensitive connections
	always @(*) begin
		eq_471_in0 = valid ? 32'd4 : 32'd4;
		eq_471_in1 = valid ? state_4_last_state : state_4_last_state;
	end
	// controller for eq_474.eq_474_in0
	// controller for eq_474.eq_474_in1
	// Insensitive connections
	always @(*) begin
		eq_474_in0 = valid ? 32'd1 : 32'd1;
		eq_474_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_479.eq_479_in0
	// controller for eq_479.eq_479_in1
	// Insensitive connections
	always @(*) begin
		eq_479_in0 = valid ? 32'd3 : 32'd3;
		eq_479_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_484.eq_484_in0
	// controller for eq_484.eq_484_in1
	// Insensitive connections
	always @(*) begin
		eq_484_in0 = valid ? 32'd3 : 32'd3;
		eq_484_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_489.eq_489_in0
	// controller for eq_489.eq_489_in1
	// Insensitive connections
	always @(*) begin
		eq_489_in0 = valid ? 32'd3 : 32'd3;
		eq_489_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_494.eq_494_in0
	// controller for eq_494.eq_494_in1
	// Insensitive connections
	always @(*) begin
		eq_494_in0 = valid ? 32'd3 : 32'd3;
		eq_494_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_499.eq_499_in0
	// controller for eq_499.eq_499_in1
	// Insensitive connections
	always @(*) begin
		eq_499_in0 = valid ? 32'd1 : 32'd1;
		eq_499_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_504.eq_504_in0
	// controller for eq_504.eq_504_in1
	// Insensitive connections
	always @(*) begin
		eq_504_in0 = valid ? 32'd3 : 32'd3;
		eq_504_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_509.eq_509_in0
	// controller for eq_509.eq_509_in1
	// Insensitive connections
	always @(*) begin
		eq_509_in0 = valid ? 32'd4 : 32'd4;
		eq_509_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for eq_514.eq_514_in0
	// controller for eq_514.eq_514_in1
	// Insensitive connections
	always @(*) begin
		eq_514_in0 = valid ? 32'd4 : 32'd4;
		eq_514_in1 = valid ? 32'd4 : 32'd4;
	end
	// controller for icmp_15.cmp_in0_icmp_15
	// controller for icmp_15.cmp_in1_icmp_15
	// Insensitive connections
	always @(*) begin
		cmp_in0_icmp_15 = valid ? add_out_add_14 : add_out_add_14;
		cmp_in1_icmp_15 = valid ? 32'd4 : 32'd4;
	end
	// controller for in.in_read_valid_reg
	always @(*) begin
		if (andOp_207_out) begin 
			in_read_valid_reg = -(1'd1);
		end else begin
			in_read_valid_reg = 0;
		end
	end
	// controller for notOp_101.notOp_101_in0
	// Insensitive connections
	always @(*) begin
		notOp_101_in0 = valid ? andOp_100_out : andOp_100_out;
	end
	// controller for notOp_103.notOp_103_in0
	// Insensitive connections
	always @(*) begin
		notOp_103_in0 = valid ? in_read_ready : in_read_ready;
	end
	// controller for notOp_107.notOp_107_in0
	// Insensitive connections
	always @(*) begin
		notOp_107_in0 = valid ? andOp_106_out : andOp_106_out;
	end
	// controller for notOp_110.notOp_110_in0
	// Insensitive connections
	always @(*) begin
		notOp_110_in0 = valid ? andOp_109_out : andOp_109_out;
	end
	// controller for notOp_113.notOp_113_in0
	// Insensitive connections
	always @(*) begin
		notOp_113_in0 = valid ? andOp_112_out : andOp_112_out;
	end
	// controller for notOp_116.notOp_116_in0
	// Insensitive connections
	always @(*) begin
		notOp_116_in0 = valid ? andOp_115_out : andOp_115_out;
	end
	// controller for notOp_118.notOp_118_in0
	// Insensitive connections
	always @(*) begin
		notOp_118_in0 = valid ? data_in_4_81_out_data : data_in_4_81_out_data;
	end
	// controller for notOp_122.notOp_122_in0
	// Insensitive connections
	always @(*) begin
		notOp_122_in0 = valid ? andOp_121_out : andOp_121_out;
	end
	// controller for notOp_125.notOp_125_in0
	// Insensitive connections
	always @(*) begin
		notOp_125_in0 = valid ? andOp_124_out : andOp_124_out;
	end
	// controller for notOp_128.notOp_128_in0
	// Insensitive connections
	always @(*) begin
		notOp_128_in0 = valid ? andOp_127_out : andOp_127_out;
	end
	// controller for notOp_130.notOp_130_in0
	// Insensitive connections
	always @(*) begin
		notOp_130_in0 = valid ? out_write_ready : out_write_ready;
	end
	// controller for notOp_134.notOp_134_in0
	// Insensitive connections
	always @(*) begin
		notOp_134_in0 = valid ? andOp_133_out : andOp_133_out;
	end
	// controller for notOp_137.notOp_137_in0
	// Insensitive connections
	always @(*) begin
		notOp_137_in0 = valid ? andOp_136_out : andOp_136_out;
	end
	// controller for notOp_139.notOp_139_in0
	// Insensitive connections
	always @(*) begin
		notOp_139_in0 = valid ? data_in_4_81_out_data : data_in_4_81_out_data;
	end
	// controller for notOp_166.notOp_166_in0
	// Insensitive connections
	always @(*) begin
		notOp_166_in0 = valid ? eq_165_out : eq_165_out;
	end
	// controller for notOp_169.notOp_169_in0
	// Insensitive connections
	always @(*) begin
		notOp_169_in0 = valid ? eq_168_out : eq_168_out;
	end
	// controller for notOp_172.notOp_172_in0
	// Insensitive connections
	always @(*) begin
		notOp_172_in0 = valid ? eq_171_out : eq_171_out;
	end
	// controller for notOp_178.notOp_178_in0
	// Insensitive connections
	always @(*) begin
		notOp_178_in0 = valid ? eq_177_out : eq_177_out;
	end
	// controller for notOp_181.notOp_181_in0
	// Insensitive connections
	always @(*) begin
		notOp_181_in0 = valid ? eq_180_out : eq_180_out;
	end
	// controller for notOp_184.notOp_184_in0
	// Insensitive connections
	always @(*) begin
		notOp_184_in0 = valid ? eq_183_out : eq_183_out;
	end
	// controller for notOp_187.notOp_187_in0
	// Insensitive connections
	always @(*) begin
		notOp_187_in0 = valid ? eq_186_out : eq_186_out;
	end
	// controller for notOp_190.notOp_190_in0
	// Insensitive connections
	always @(*) begin
		notOp_190_in0 = valid ? eq_189_out : eq_189_out;
	end
	// controller for notOp_194.notOp_194_in0
	// Insensitive connections
	always @(*) begin
		notOp_194_in0 = valid ? eq_193_out : eq_193_out;
	end
	// controller for notOp_223.notOp_223_in0
	// Insensitive connections
	always @(*) begin
		notOp_223_in0 = valid ? andOp_104_out : andOp_104_out;
	end
	// controller for notOp_225.notOp_225_in0
	// Insensitive connections
	always @(*) begin
		notOp_225_in0 = valid ? andOp_119_out : andOp_119_out;
	end
	// controller for notOp_227.notOp_227_in0
	// Insensitive connections
	always @(*) begin
		notOp_227_in0 = valid ? andOp_219_out : andOp_219_out;
	end
	// controller for notOp_229.notOp_229_in0
	// Insensitive connections
	always @(*) begin
		notOp_229_in0 = valid ? andOp_102_out : andOp_102_out;
	end
	// controller for notOp_231.notOp_231_in0
	// Insensitive connections
	always @(*) begin
		notOp_231_in0 = valid ? andOp_220_out : andOp_220_out;
	end
	// controller for notOp_233.notOp_233_in0
	// Insensitive connections
	always @(*) begin
		notOp_233_in0 = valid ? andOp_131_out : andOp_131_out;
	end
	// controller for notOp_235.notOp_235_in0
	// Insensitive connections
	always @(*) begin
		notOp_235_in0 = valid ? andOp_221_out : andOp_221_out;
	end
	// controller for notOp_237.notOp_237_in0
	// Insensitive connections
	always @(*) begin
		notOp_237_in0 = valid ? andOp_222_out : andOp_222_out;
	end
	// controller for notOp_256.notOp_256_in0
	// Insensitive connections
	always @(*) begin
		notOp_256_in0 = valid ? eq_254_out : eq_254_out;
	end
	// controller for notOp_261.notOp_261_in0
	// Insensitive connections
	always @(*) begin
		notOp_261_in0 = valid ? eq_259_out : eq_259_out;
	end
	// controller for notOp_266.notOp_266_in0
	// Insensitive connections
	always @(*) begin
		notOp_266_in0 = valid ? eq_264_out : eq_264_out;
	end
	// controller for notOp_271.notOp_271_in0
	// Insensitive connections
	always @(*) begin
		notOp_271_in0 = valid ? eq_269_out : eq_269_out;
	end
	// controller for notOp_276.notOp_276_in0
	// Insensitive connections
	always @(*) begin
		notOp_276_in0 = valid ? eq_274_out : eq_274_out;
	end
	// controller for notOp_281.notOp_281_in0
	// Insensitive connections
	always @(*) begin
		notOp_281_in0 = valid ? eq_279_out : eq_279_out;
	end
	// controller for notOp_286.notOp_286_in0
	// Insensitive connections
	always @(*) begin
		notOp_286_in0 = valid ? eq_284_out : eq_284_out;
	end
	// controller for notOp_291.notOp_291_in0
	// Insensitive connections
	always @(*) begin
		notOp_291_in0 = valid ? eq_289_out : eq_289_out;
	end
	// controller for notOp_296.notOp_296_in0
	// Insensitive connections
	always @(*) begin
		notOp_296_in0 = valid ? eq_294_out : eq_294_out;
	end
	// controller for notOp_311.notOp_311_in0
	// Insensitive connections
	always @(*) begin
		notOp_311_in0 = valid ? eq_309_out : eq_309_out;
	end
	// controller for notOp_316.notOp_316_in0
	// Insensitive connections
	always @(*) begin
		notOp_316_in0 = valid ? eq_314_out : eq_314_out;
	end
	// controller for notOp_321.notOp_321_in0
	// Insensitive connections
	always @(*) begin
		notOp_321_in0 = valid ? eq_319_out : eq_319_out;
	end
	// controller for notOp_326.notOp_326_in0
	// Insensitive connections
	always @(*) begin
		notOp_326_in0 = valid ? eq_324_out : eq_324_out;
	end
	// controller for notOp_331.notOp_331_in0
	// Insensitive connections
	always @(*) begin
		notOp_331_in0 = valid ? eq_329_out : eq_329_out;
	end
	// controller for notOp_336.notOp_336_in0
	// Insensitive connections
	always @(*) begin
		notOp_336_in0 = valid ? eq_334_out : eq_334_out;
	end
	// controller for notOp_341.notOp_341_in0
	// Insensitive connections
	always @(*) begin
		notOp_341_in0 = valid ? eq_339_out : eq_339_out;
	end
	// controller for notOp_346.notOp_346_in0
	// Insensitive connections
	always @(*) begin
		notOp_346_in0 = valid ? eq_344_out : eq_344_out;
	end
	// controller for notOp_351.notOp_351_in0
	// Insensitive connections
	always @(*) begin
		notOp_351_in0 = valid ? eq_349_out : eq_349_out;
	end
	// controller for notOp_366.notOp_366_in0
	// Insensitive connections
	always @(*) begin
		notOp_366_in0 = valid ? eq_364_out : eq_364_out;
	end
	// controller for notOp_371.notOp_371_in0
	// Insensitive connections
	always @(*) begin
		notOp_371_in0 = valid ? eq_369_out : eq_369_out;
	end
	// controller for notOp_376.notOp_376_in0
	// Insensitive connections
	always @(*) begin
		notOp_376_in0 = valid ? eq_374_out : eq_374_out;
	end
	// controller for notOp_381.notOp_381_in0
	// Insensitive connections
	always @(*) begin
		notOp_381_in0 = valid ? eq_379_out : eq_379_out;
	end
	// controller for notOp_386.notOp_386_in0
	// Insensitive connections
	always @(*) begin
		notOp_386_in0 = valid ? eq_384_out : eq_384_out;
	end
	// controller for notOp_391.notOp_391_in0
	// Insensitive connections
	always @(*) begin
		notOp_391_in0 = valid ? eq_389_out : eq_389_out;
	end
	// controller for notOp_396.notOp_396_in0
	// Insensitive connections
	always @(*) begin
		notOp_396_in0 = valid ? eq_394_out : eq_394_out;
	end
	// controller for notOp_401.notOp_401_in0
	// Insensitive connections
	always @(*) begin
		notOp_401_in0 = valid ? eq_399_out : eq_399_out;
	end
	// controller for notOp_406.notOp_406_in0
	// Insensitive connections
	always @(*) begin
		notOp_406_in0 = valid ? eq_404_out : eq_404_out;
	end
	// controller for notOp_421.notOp_421_in0
	// Insensitive connections
	always @(*) begin
		notOp_421_in0 = valid ? eq_419_out : eq_419_out;
	end
	// controller for notOp_426.notOp_426_in0
	// Insensitive connections
	always @(*) begin
		notOp_426_in0 = valid ? eq_424_out : eq_424_out;
	end
	// controller for notOp_431.notOp_431_in0
	// Insensitive connections
	always @(*) begin
		notOp_431_in0 = valid ? eq_429_out : eq_429_out;
	end
	// controller for notOp_436.notOp_436_in0
	// Insensitive connections
	always @(*) begin
		notOp_436_in0 = valid ? eq_434_out : eq_434_out;
	end
	// controller for notOp_441.notOp_441_in0
	// Insensitive connections
	always @(*) begin
		notOp_441_in0 = valid ? eq_439_out : eq_439_out;
	end
	// controller for notOp_446.notOp_446_in0
	// Insensitive connections
	always @(*) begin
		notOp_446_in0 = valid ? eq_444_out : eq_444_out;
	end
	// controller for notOp_451.notOp_451_in0
	// Insensitive connections
	always @(*) begin
		notOp_451_in0 = valid ? eq_449_out : eq_449_out;
	end
	// controller for notOp_456.notOp_456_in0
	// Insensitive connections
	always @(*) begin
		notOp_456_in0 = valid ? eq_454_out : eq_454_out;
	end
	// controller for notOp_461.notOp_461_in0
	// Insensitive connections
	always @(*) begin
		notOp_461_in0 = valid ? eq_459_out : eq_459_out;
	end
	// controller for notOp_476.notOp_476_in0
	// Insensitive connections
	always @(*) begin
		notOp_476_in0 = valid ? eq_474_out : eq_474_out;
	end
	// controller for notOp_481.notOp_481_in0
	// Insensitive connections
	always @(*) begin
		notOp_481_in0 = valid ? eq_479_out : eq_479_out;
	end
	// controller for notOp_486.notOp_486_in0
	// Insensitive connections
	always @(*) begin
		notOp_486_in0 = valid ? eq_484_out : eq_484_out;
	end
	// controller for notOp_491.notOp_491_in0
	// Insensitive connections
	always @(*) begin
		notOp_491_in0 = valid ? eq_489_out : eq_489_out;
	end
	// controller for notOp_496.notOp_496_in0
	// Insensitive connections
	always @(*) begin
		notOp_496_in0 = valid ? eq_494_out : eq_494_out;
	end
	// controller for notOp_501.notOp_501_in0
	// Insensitive connections
	always @(*) begin
		notOp_501_in0 = valid ? eq_499_out : eq_499_out;
	end
	// controller for notOp_506.notOp_506_in0
	// Insensitive connections
	always @(*) begin
		notOp_506_in0 = valid ? eq_504_out : eq_504_out;
	end
	// controller for notOp_511.notOp_511_in0
	// Insensitive connections
	always @(*) begin
		notOp_511_in0 = valid ? eq_509_out : eq_509_out;
	end
	// controller for notOp_516.notOp_516_in0
	// Insensitive connections
	always @(*) begin
		notOp_516_in0 = valid ? eq_514_out : eq_514_out;
	end
	// controller for notOp_92.notOp_92_in0
	// Insensitive connections
	always @(*) begin
		notOp_92_in0 = valid ? andOp_91_out : andOp_91_out;
	end
	// controller for notOp_95.notOp_95_in0
	// Insensitive connections
	always @(*) begin
		notOp_95_in0 = valid ? andOp_94_out : andOp_94_out;
	end
	// controller for notOp_98.notOp_98_in0
	// Insensitive connections
	always @(*) begin
		notOp_98_in0 = valid ? andOp_97_out : andOp_97_out;
	end
	// controller for orOp_143.orOp_143_in0
	// controller for orOp_143.orOp_143_in1
	// Insensitive connections
	always @(*) begin
		orOp_143_in0 = valid ? eq_142_out : eq_142_out;
		orOp_143_in1 = valid ? andOp_91_out : andOp_91_out;
	end
	// controller for orOp_145.orOp_145_in0
	// controller for orOp_145.orOp_145_in1
	// Insensitive connections
	always @(*) begin
		orOp_145_in0 = valid ? eq_144_out : eq_144_out;
		orOp_145_in1 = valid ? andOp_94_out : andOp_94_out;
	end
	// controller for orOp_147.orOp_147_in0
	// controller for orOp_147.orOp_147_in1
	// Insensitive connections
	always @(*) begin
		orOp_147_in0 = valid ? eq_146_out : eq_146_out;
		orOp_147_in1 = valid ? andOp_97_out : andOp_97_out;
	end
	// controller for orOp_152.orOp_152_in0
	// controller for orOp_152.orOp_152_in1
	// Insensitive connections
	always @(*) begin
		orOp_152_in0 = valid ? eq_151_out : eq_151_out;
		orOp_152_in1 = valid ? andOp_109_out : andOp_109_out;
	end
	// controller for orOp_154.orOp_154_in0
	// controller for orOp_154.orOp_154_in1
	// Insensitive connections
	always @(*) begin
		orOp_154_in0 = valid ? eq_153_out : eq_153_out;
		orOp_154_in1 = valid ? andOp_117_out : andOp_117_out;
	end
	// controller for orOp_156.orOp_156_in0
	// controller for orOp_156.orOp_156_in1
	// Insensitive connections
	always @(*) begin
		orOp_156_in0 = valid ? eq_155_out : eq_155_out;
		orOp_156_in1 = valid ? andOp_121_out : andOp_121_out;
	end
	// controller for orOp_158.orOp_158_in0
	// controller for orOp_158.orOp_158_in1
	// Insensitive connections
	always @(*) begin
		orOp_158_in0 = valid ? eq_157_out : eq_157_out;
		orOp_158_in1 = valid ? andOp_124_out : andOp_124_out;
	end
	// controller for orOp_160.orOp_160_in0
	// controller for orOp_160.orOp_160_in1
	// Insensitive connections
	always @(*) begin
		orOp_160_in0 = valid ? eq_159_out : eq_159_out;
		orOp_160_in1 = valid ? andOp_129_out : andOp_129_out;
	end
	// controller for orOp_163.orOp_163_in0
	// controller for orOp_163.orOp_163_in1
	// Insensitive connections
	always @(*) begin
		orOp_163_in0 = valid ? eq_162_out : eq_162_out;
		orOp_163_in1 = valid ? andOp_133_out : andOp_133_out;
	end
	// controller for out.out_in_data_reg
	always @(*) begin
		if (andOp_218_out) begin 
			out_in_data_reg = rdata_ram_0;
		end else begin
			out_in_data_reg = 0;
		end
	end
	// controller for out.out_write_valid_reg
	always @(*) begin
		if (andOp_216_out) begin 
			out_write_valid_reg = -(1'd1);
		end else begin
			out_write_valid_reg = 0;
		end
	end
	// controller for phi_6.phi_in_phi_6
	// controller for phi_6.phi_last_block_phi_6
	// controller for phi_6.phi_s_phi_6
	// Insensitive connections
	always @(*) begin
		phi_in_phi_6 = valid ? concat_204_out : concat_204_out;
		phi_last_block_phi_6 = valid ? bb_3_predecessor_in_state_1_out_data : bb_3_predecessor_in_state_1_out_data;
		phi_s_phi_6 = valid ? concat_205_out : concat_205_out;
	end
	// controller for ram_0.raddr_ram_0_reg
	always @(*) begin
		if (andOp_198_out) begin 
			raddr_ram_0_reg = 32'd0;
		end else if (andOp_200_out) begin 
			raddr_ram_0_reg = 32'd0;
		end else begin
			raddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.waddr_ram_0_reg
	always @(*) begin
		if (andOp_197_out) begin 
			waddr_ram_0_reg = 32'd0;
		end else if (andOp_199_out) begin 
			waddr_ram_0_reg = 32'd0;
		end else begin
			waddr_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wdata_ram_0_reg
	always @(*) begin
		if (andOp_197_out) begin 
			wdata_ram_0_reg = 32'd0;
		end else if (andOp_199_out) begin 
			wdata_ram_0_reg = add_out_add_12;
		end else begin
			wdata_ram_0_reg = 0;
		end
	end
	// controller for ram_0.wen_ram_0_reg
	always @(*) begin
		if (andOp_197_out) begin 
			wen_ram_0_reg = 1'd1;
		end else if (andOp_199_out) begin 
			wen_ram_0_reg = 1'd1;
		end else begin
			wen_ram_0_reg = 0;
		end
	end
	// controller for ret_19.valid_reg
	always @(*) begin
		if (andOp_215_out) begin 
			valid_reg = 1'd1;
		end else begin
			valid_reg = 0;
		end
	end
	// controller for tmp_output_210.tmp_output_210_in_data
	always @(*) begin
		if (eq_211_out) begin 
			tmp_output_210_in_data = in_out_data;
		end else begin
			tmp_output_210_in_data = 0;
		end
	end
	// Register controllers
	always @(posedge clk) begin
		if (rst) begin
			add_tmp_4 <= 0;
		end else begin
			if (andOp_240_out) begin
				add_tmp_4 <= add_out_add_14;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			call_tmp_6 <= 0;
		end else begin
			if (andOp_242_out) begin
				call_tmp_6 <= in_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_0 <= 0;
		end else begin
			if (andOp_255_out) begin
				data_store_0_0 <= phi_out_phi_6;
			end
			if (andOp_257_out) begin
				data_store_0_0 <= data_in_0_1_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_10 <= 0;
		end else begin
			if (andOp_280_out) begin
				data_store_0_10 <= in_read_ready;
			end
			if (andOp_282_out) begin
				data_store_0_10 <= data_in_0_11_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_12 <= 0;
		end else begin
			if (andOp_285_out) begin
				data_store_0_12 <= in_out_data;
			end
			if (andOp_287_out) begin
				data_store_0_12 <= data_in_0_13_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_14 <= 0;
		end else begin
			if (andOp_290_out) begin
				data_store_0_14 <= out_write_ready;
			end
			if (andOp_292_out) begin
				data_store_0_14 <= data_in_0_15_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_16 <= 0;
		end else begin
			if (andOp_295_out) begin
				data_store_0_16 <= rdata_ram_0;
			end
			if (andOp_297_out) begin
				data_store_0_16 <= data_in_0_17_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_2 <= 0;
		end else begin
			if (andOp_260_out) begin
				data_store_0_2 <= rdata_ram_0;
			end
			if (andOp_262_out) begin
				data_store_0_2 <= data_in_0_3_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_4 <= 0;
		end else begin
			if (andOp_265_out) begin
				data_store_0_4 <= add_out_add_12;
			end
			if (andOp_267_out) begin
				data_store_0_4 <= data_in_0_5_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_6 <= 0;
		end else begin
			if (andOp_270_out) begin
				data_store_0_6 <= add_out_add_14;
			end
			if (andOp_272_out) begin
				data_store_0_6 <= data_in_0_7_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_0_8 <= 0;
		end else begin
			if (andOp_275_out) begin
				data_store_0_8 <= cmp_out_icmp_15;
			end
			if (andOp_277_out) begin
				data_store_0_8 <= data_in_0_9_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_18 <= 0;
		end else begin
			if (andOp_310_out) begin
				data_store_1_18 <= phi_out_phi_6;
			end
			if (andOp_312_out) begin
				data_store_1_18 <= data_in_1_19_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_20 <= 0;
		end else begin
			if (andOp_315_out) begin
				data_store_1_20 <= rdata_ram_0;
			end
			if (andOp_317_out) begin
				data_store_1_20 <= data_in_1_21_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_22 <= 0;
		end else begin
			if (andOp_320_out) begin
				data_store_1_22 <= add_out_add_12;
			end
			if (andOp_322_out) begin
				data_store_1_22 <= data_in_1_23_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_24 <= 0;
		end else begin
			if (andOp_325_out) begin
				data_store_1_24 <= add_out_add_14;
			end
			if (andOp_327_out) begin
				data_store_1_24 <= data_in_1_25_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_26 <= 0;
		end else begin
			if (andOp_330_out) begin
				data_store_1_26 <= cmp_out_icmp_15;
			end
			if (andOp_332_out) begin
				data_store_1_26 <= data_in_1_27_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_28 <= 0;
		end else begin
			if (andOp_335_out) begin
				data_store_1_28 <= in_read_ready;
			end
			if (andOp_337_out) begin
				data_store_1_28 <= data_in_1_29_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_30 <= 0;
		end else begin
			if (andOp_340_out) begin
				data_store_1_30 <= in_out_data;
			end
			if (andOp_342_out) begin
				data_store_1_30 <= data_in_1_31_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_32 <= 0;
		end else begin
			if (andOp_345_out) begin
				data_store_1_32 <= out_write_ready;
			end
			if (andOp_347_out) begin
				data_store_1_32 <= data_in_1_33_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_1_34 <= 0;
		end else begin
			if (andOp_350_out) begin
				data_store_1_34 <= rdata_ram_0;
			end
			if (andOp_352_out) begin
				data_store_1_34 <= data_in_1_35_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_36 <= 0;
		end else begin
			if (andOp_365_out) begin
				data_store_2_36 <= phi_out_phi_6;
			end
			if (andOp_367_out) begin
				data_store_2_36 <= data_in_2_37_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_38 <= 0;
		end else begin
			if (andOp_370_out) begin
				data_store_2_38 <= rdata_ram_0;
			end
			if (andOp_372_out) begin
				data_store_2_38 <= data_in_2_39_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_40 <= 0;
		end else begin
			if (andOp_375_out) begin
				data_store_2_40 <= add_out_add_12;
			end
			if (andOp_377_out) begin
				data_store_2_40 <= data_in_2_41_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_42 <= 0;
		end else begin
			if (andOp_380_out) begin
				data_store_2_42 <= add_out_add_14;
			end
			if (andOp_382_out) begin
				data_store_2_42 <= data_in_2_43_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_44 <= 0;
		end else begin
			if (andOp_385_out) begin
				data_store_2_44 <= cmp_out_icmp_15;
			end
			if (andOp_387_out) begin
				data_store_2_44 <= data_in_2_45_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_46 <= 0;
		end else begin
			if (andOp_390_out) begin
				data_store_2_46 <= in_read_ready;
			end
			if (andOp_392_out) begin
				data_store_2_46 <= data_in_2_47_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_48 <= 0;
		end else begin
			if (andOp_395_out) begin
				data_store_2_48 <= in_out_data;
			end
			if (andOp_397_out) begin
				data_store_2_48 <= data_in_2_49_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_50 <= 0;
		end else begin
			if (andOp_400_out) begin
				data_store_2_50 <= out_write_ready;
			end
			if (andOp_402_out) begin
				data_store_2_50 <= data_in_2_51_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_2_52 <= 0;
		end else begin
			if (andOp_405_out) begin
				data_store_2_52 <= rdata_ram_0;
			end
			if (andOp_407_out) begin
				data_store_2_52 <= data_in_2_53_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_54 <= 0;
		end else begin
			if (andOp_420_out) begin
				data_store_3_54 <= phi_out_phi_6;
			end
			if (andOp_422_out) begin
				data_store_3_54 <= data_in_3_55_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_56 <= 0;
		end else begin
			if (andOp_425_out) begin
				data_store_3_56 <= rdata_ram_0;
			end
			if (andOp_427_out) begin
				data_store_3_56 <= data_in_3_57_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_58 <= 0;
		end else begin
			if (andOp_430_out) begin
				data_store_3_58 <= add_out_add_12;
			end
			if (andOp_432_out) begin
				data_store_3_58 <= data_in_3_59_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_60 <= 0;
		end else begin
			if (andOp_435_out) begin
				data_store_3_60 <= add_out_add_14;
			end
			if (andOp_437_out) begin
				data_store_3_60 <= data_in_3_61_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_62 <= 0;
		end else begin
			if (andOp_440_out) begin
				data_store_3_62 <= cmp_out_icmp_15;
			end
			if (andOp_442_out) begin
				data_store_3_62 <= data_in_3_63_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_64 <= 0;
		end else begin
			if (andOp_445_out) begin
				data_store_3_64 <= in_read_ready;
			end
			if (andOp_447_out) begin
				data_store_3_64 <= data_in_3_65_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_66 <= 0;
		end else begin
			if (andOp_450_out) begin
				data_store_3_66 <= in_out_data;
			end
			if (andOp_452_out) begin
				data_store_3_66 <= data_in_3_67_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_68 <= 0;
		end else begin
			if (andOp_455_out) begin
				data_store_3_68 <= out_write_ready;
			end
			if (andOp_457_out) begin
				data_store_3_68 <= data_in_3_69_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_3_70 <= 0;
		end else begin
			if (andOp_460_out) begin
				data_store_3_70 <= rdata_ram_0;
			end
			if (andOp_462_out) begin
				data_store_3_70 <= data_in_3_71_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_72 <= 0;
		end else begin
			if (andOp_475_out) begin
				data_store_4_72 <= phi_out_phi_6;
			end
			if (andOp_477_out) begin
				data_store_4_72 <= data_in_4_73_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_74 <= 0;
		end else begin
			if (andOp_480_out) begin
				data_store_4_74 <= rdata_ram_0;
			end
			if (andOp_482_out) begin
				data_store_4_74 <= data_in_4_75_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_76 <= 0;
		end else begin
			if (andOp_485_out) begin
				data_store_4_76 <= add_out_add_12;
			end
			if (andOp_487_out) begin
				data_store_4_76 <= data_in_4_77_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_78 <= 0;
		end else begin
			if (andOp_490_out) begin
				data_store_4_78 <= add_out_add_14;
			end
			if (andOp_492_out) begin
				data_store_4_78 <= data_in_4_79_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_80 <= 0;
		end else begin
			if (andOp_495_out) begin
				data_store_4_80 <= cmp_out_icmp_15;
			end
			if (andOp_497_out) begin
				data_store_4_80 <= data_in_4_81_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_82 <= 0;
		end else begin
			if (andOp_500_out) begin
				data_store_4_82 <= in_read_ready;
			end
			if (andOp_502_out) begin
				data_store_4_82 <= data_in_4_83_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_84 <= 0;
		end else begin
			if (andOp_505_out) begin
				data_store_4_84 <= in_out_data;
			end
			if (andOp_507_out) begin
				data_store_4_84 <= data_in_4_85_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_86 <= 0;
		end else begin
			if (andOp_510_out) begin
				data_store_4_86 <= out_write_ready;
			end
			if (andOp_512_out) begin
				data_store_4_86 <= data_in_4_87_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			data_store_4_88 <= 0;
		end else begin
			if (andOp_515_out) begin
				data_store_4_88 <= rdata_ram_0;
			end
			if (andOp_517_out) begin
				data_store_4_88 <= data_in_4_89_out_data;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			global_state <= 0;
		end else begin
			if (andOp_102_out) begin
				global_state <= 32'd2;
			end
			if (andOp_104_out) begin
				global_state <= 32'd1;
			end
			if (andOp_119_out) begin
				global_state <= 32'd1;
			end
			if (andOp_131_out) begin
				global_state <= 32'd4;
			end
			if (andOp_219_out) begin
				global_state <= 32'd1;
			end
			if (andOp_220_out) begin
				global_state <= 32'd3;
			end
			if (andOp_221_out) begin
				global_state <= 32'd4;
			end
			if (andOp_222_out) begin
				global_state <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			icmp_tmp_5 <= 0;
		end else begin
			if (andOp_241_out) begin
				icmp_tmp_5 <= cmp_out_icmp_15;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			phi_tmp_0 <= 0;
		end else begin
			if (andOp_239_out) begin
				phi_tmp_0 <= phi_out_phi_6;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_entry_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_is_active <= 1;
		end else begin
			if (1'd1) begin
				state_0_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_BB_reg <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_0_last_state <= 0;
		end else begin
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_entry_BB_reg <= 0;
		end else begin
			if (andOp_104_out) begin
				state_1_entry_BB_reg <= 32'd9;
			end
			if (andOp_119_out) begin
				state_1_entry_BB_reg <= 32'd3;
			end
			if (andOp_219_out) begin
				state_1_entry_BB_reg <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_is_active <= 0;
		end else begin
			if (andOp_104_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_119_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_219_out) begin
				state_1_is_active <= 1'd1;
			end
			if (andOp_228_out) begin
				state_1_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_BB_reg <= 0;
		end else begin
			if (andOp_104_out) begin
				state_1_last_BB_reg <= 32'd9;
			end
			if (andOp_119_out) begin
				state_1_last_BB_reg <= 32'd4;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_1_last_state <= 0;
		end else begin
			if (andOp_104_out) begin
				state_1_last_state <= 32'd1;
			end
			if (andOp_119_out) begin
				state_1_last_state <= 32'd4;
			end
			if (andOp_219_out) begin
				state_1_last_state <= 32'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_entry_BB_reg <= 0;
		end else begin
			if (andOp_102_out) begin
				state_2_entry_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_is_active <= 0;
		end else begin
			if (andOp_102_out) begin
				state_2_is_active <= 1'd1;
			end
			if (andOp_230_out) begin
				state_2_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_BB_reg <= 0;
		end else begin
			if (andOp_102_out) begin
				state_2_last_BB_reg <= 32'd9;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_2_last_state <= 0;
		end else begin
			if (andOp_102_out) begin
				state_2_last_state <= 32'd1;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_entry_BB_reg <= 0;
		end else begin
			if (andOp_220_out) begin
				state_3_entry_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_is_active <= 0;
		end else begin
			if (andOp_220_out) begin
				state_3_is_active <= 1'd1;
			end
			if (andOp_232_out) begin
				state_3_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_BB_reg <= 0;
		end else begin
			if (andOp_109_out) begin
				state_3_last_BB_reg <= 32'd10;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_3_last_state <= 0;
		end else begin
			if (andOp_220_out) begin
				state_3_last_state <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_entry_BB_reg <= 0;
		end else begin
			if (andOp_131_out) begin
				state_4_entry_BB_reg <= 32'd6;
			end
			if (andOp_221_out) begin
				state_4_entry_BB_reg <= 32'd4;
			end
			if (andOp_222_out) begin
				state_4_entry_BB_reg <= 32'd2;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_is_active <= 0;
		end else begin
			if (andOp_131_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_221_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_222_out) begin
				state_4_is_active <= 1'd1;
			end
			if (andOp_238_out) begin
				state_4_is_active <= 1'd0;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_BB_reg <= 0;
		end else begin
			if (andOp_131_out) begin
				state_4_last_BB_reg <= 32'd6;
			end
			if (andOp_133_out) begin
				state_4_last_BB_reg <= 32'd7;
			end
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state_4_last_state <= 0;
		end else begin
			if (andOp_131_out) begin
				state_4_last_state <= 32'd4;
			end
			if (andOp_221_out) begin
				state_4_last_state <= 32'd3;
			end
			if (andOp_222_out) begin
				state_4_last_state <= 32'd4;
			end
		end
	end

endmodule

